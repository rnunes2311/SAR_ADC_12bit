magic
tech sky130A
magscale 1 2
timestamp 1715456343
<< pwell >>
rect -400 23970 -220 24000
rect -115 23970 70 24000
rect -400 23940 70 23970
rect 12740 23940 13140 24000
rect -400 -330 13140 23940
<< psubdiff >>
rect -304 23840 -280 23880
rect 13000 23840 13024 23880
rect -370 23740 -330 23770
rect -370 -100 -330 -70
rect -304 -210 -280 -170
rect 13000 -210 13024 -170
<< psubdiffcont >>
rect -280 23840 13000 23880
rect -370 -70 -330 23740
rect -280 -210 13000 -170
<< locali >>
rect -215 24130 -155 24170
rect -205 23880 -165 24130
rect 12980 24075 13040 24115
rect 12995 23880 13035 24075
rect -370 23740 -330 23880
rect -296 23840 -280 23880
rect 13000 23840 13035 23880
rect -370 -140 -330 -70
rect -296 -210 -280 -170
rect 13000 -210 13016 -170
<< viali >>
rect -255 24130 -215 24170
rect -155 24130 -115 24170
rect 12940 24075 12980 24115
rect 13040 24075 13080 24115
rect -270 23840 12910 23880
rect -370 -50 -330 23740
rect -220 -210 12960 -170
<< metal1 >>
rect -275 24120 -265 24180
rect -205 24025 -165 24180
rect -105 24120 -95 24180
rect 12920 24065 12930 24125
rect 12990 24025 13030 24125
rect 13090 24065 13100 24125
rect -370 24015 0 24025
rect -370 23955 -366 24015
rect -314 23955 -56 24015
rect -4 23955 0 24015
rect -370 23886 0 23955
rect 30 24015 400 24025
rect 30 23955 34 24015
rect 86 23955 344 24015
rect 396 23955 400 24015
rect 30 23886 400 23955
rect 430 24015 800 24025
rect 430 23955 434 24015
rect 486 23955 744 24015
rect 796 23955 800 24015
rect 430 23886 800 23955
rect 830 24015 1200 24025
rect 830 23955 834 24015
rect 886 23955 1144 24015
rect 1196 23955 1200 24015
rect 830 23886 1200 23955
rect 1230 24015 1600 24025
rect 1230 23955 1234 24015
rect 1286 23955 1544 24015
rect 1596 23955 1600 24015
rect 1230 23886 1600 23955
rect 1630 24015 2000 24025
rect 1630 23955 1634 24015
rect 1686 23955 1944 24015
rect 1996 23955 2000 24015
rect 1630 23886 2000 23955
rect 2030 24015 2400 24025
rect 2030 23955 2034 24015
rect 2086 23955 2344 24015
rect 2396 23955 2400 24015
rect 2030 23886 2400 23955
rect 2430 24015 2800 24025
rect 2430 23955 2434 24015
rect 2486 23955 2744 24015
rect 2796 23955 2800 24015
rect 2430 23886 2800 23955
rect 2830 24015 3200 24025
rect 2830 23955 2834 24015
rect 2886 23955 3144 24015
rect 3196 23955 3200 24015
rect 2830 23886 3200 23955
rect 3230 24015 3600 24025
rect 3230 23955 3234 24015
rect 3286 23955 3544 24015
rect 3596 23955 3600 24015
rect 3230 23886 3600 23955
rect 3630 24015 4000 24025
rect 3630 23955 3634 24015
rect 3686 23955 3944 24015
rect 3996 23955 4000 24015
rect 3630 23886 4000 23955
rect 4030 24015 4400 24025
rect 4030 23955 4034 24015
rect 4086 23955 4344 24015
rect 4396 23955 4400 24015
rect 4030 23886 4400 23955
rect 4430 24015 4800 24025
rect 4430 23955 4434 24015
rect 4486 23955 4744 24015
rect 4796 23955 4800 24015
rect 4430 23886 4800 23955
rect 4830 24015 5200 24025
rect 4830 23955 4834 24015
rect 4886 23955 5144 24015
rect 5196 23955 5200 24015
rect 4830 23886 5200 23955
rect 5230 24015 5600 24025
rect 5230 23955 5234 24015
rect 5286 23955 5544 24015
rect 5596 23955 5600 24015
rect 5230 23886 5600 23955
rect 5630 24015 6000 24025
rect 5630 23955 5634 24015
rect 5686 23955 5944 24015
rect 5996 23955 6000 24015
rect 5630 23886 6000 23955
rect 6030 24015 6400 24025
rect 6030 23955 6034 24015
rect 6086 23955 6344 24015
rect 6396 23955 6400 24015
rect 6030 23886 6400 23955
rect 6430 24015 6800 24025
rect 6430 23955 6434 24015
rect 6486 23955 6744 24015
rect 6796 23955 6800 24015
rect 6430 23886 6800 23955
rect 6830 24015 7200 24025
rect 6830 23955 6834 24015
rect 6886 23955 7144 24015
rect 7196 23955 7200 24015
rect 6830 23886 7200 23955
rect 7230 24015 7600 24025
rect 7230 23955 7234 24015
rect 7286 23955 7544 24015
rect 7596 23955 7600 24015
rect 7230 23886 7600 23955
rect 7630 24015 8000 24025
rect 7630 23955 7634 24015
rect 7686 23955 7944 24015
rect 7996 23955 8000 24015
rect 7630 23886 8000 23955
rect 8030 24015 8400 24025
rect 8030 23955 8034 24015
rect 8086 23955 8344 24015
rect 8396 23955 8400 24015
rect 8030 23886 8400 23955
rect 8430 24015 8800 24025
rect 8430 23955 8434 24015
rect 8486 23955 8744 24015
rect 8796 23955 8800 24015
rect 8430 23886 8800 23955
rect 8830 24015 9200 24025
rect 8830 23955 8834 24015
rect 8886 23955 9144 24015
rect 9196 23955 9200 24015
rect 8830 23886 9200 23955
rect 9230 24015 9600 24025
rect 9230 23955 9234 24015
rect 9286 23955 9544 24015
rect 9596 23955 9600 24015
rect 9230 23886 9600 23955
rect 9630 24015 10000 24025
rect 9630 23955 9634 24015
rect 9686 23955 9944 24015
rect 9996 23955 10000 24015
rect 9630 23886 10000 23955
rect 10030 24015 10400 24025
rect 10030 23955 10034 24015
rect 10086 23955 10344 24015
rect 10396 23955 10400 24015
rect 10030 23886 10400 23955
rect 10430 24015 10800 24025
rect 10430 23955 10434 24015
rect 10486 23955 10744 24015
rect 10796 23955 10800 24015
rect 10430 23886 10800 23955
rect 10830 24015 11200 24025
rect 10830 23955 10834 24015
rect 10886 23955 11144 24015
rect 11196 23955 11200 24015
rect 10830 23886 11200 23955
rect 11230 24015 11600 24025
rect 11230 23955 11234 24015
rect 11286 23955 11544 24015
rect 11596 23955 11600 24015
rect 11230 23886 11600 23955
rect 11630 24015 12000 24025
rect 11630 23955 11634 24015
rect 11686 23955 11944 24015
rect 11996 23955 12000 24015
rect 11630 23886 12000 23955
rect 12030 24015 12400 24025
rect 12030 23955 12034 24015
rect 12086 23955 12344 24015
rect 12396 23955 12400 24015
rect 12030 23886 12400 23955
rect 12430 24015 12800 24025
rect 12430 23955 12434 24015
rect 12486 23955 12744 24015
rect 12796 23955 12800 24015
rect 12430 23886 12800 23955
rect 12830 24015 13200 24025
rect 12830 23955 12834 24015
rect 12886 23955 13144 24015
rect 13196 23955 13200 24015
rect 12830 23886 13200 23955
rect -370 23880 13200 23886
rect -370 23840 -270 23880
rect 12910 23840 13200 23880
rect -370 23834 13200 23840
rect -370 23793 0 23834
rect -376 23755 0 23793
rect -376 23740 -366 23755
rect -376 -50 -370 23740
rect -314 23695 -56 23755
rect -4 23695 0 23755
rect -330 23685 0 23695
rect 30 23755 400 23834
rect 30 23695 34 23755
rect 86 23695 344 23755
rect 396 23695 400 23755
rect 30 23685 400 23695
rect 430 23755 800 23834
rect 430 23695 434 23755
rect 486 23695 744 23755
rect 796 23695 800 23755
rect 430 23685 800 23695
rect 830 23755 1200 23834
rect 830 23695 834 23755
rect 886 23695 1144 23755
rect 1196 23695 1200 23755
rect 830 23685 1200 23695
rect 1230 23755 1600 23834
rect 1230 23695 1234 23755
rect 1286 23695 1544 23755
rect 1596 23695 1600 23755
rect 1230 23685 1600 23695
rect 1630 23755 2000 23834
rect 1630 23695 1634 23755
rect 1686 23695 1944 23755
rect 1996 23695 2000 23755
rect 1630 23685 2000 23695
rect 2030 23755 2400 23834
rect 2030 23695 2034 23755
rect 2086 23695 2344 23755
rect 2396 23695 2400 23755
rect 2030 23685 2400 23695
rect 2430 23755 2800 23834
rect 2430 23695 2434 23755
rect 2486 23695 2744 23755
rect 2796 23695 2800 23755
rect 2430 23685 2800 23695
rect 2830 23755 3200 23834
rect 2830 23695 2834 23755
rect 2886 23695 3144 23755
rect 3196 23695 3200 23755
rect 2830 23685 3200 23695
rect 3230 23755 3600 23834
rect 3230 23695 3234 23755
rect 3286 23695 3544 23755
rect 3596 23695 3600 23755
rect 3230 23685 3600 23695
rect 3630 23755 4000 23834
rect 3630 23695 3634 23755
rect 3686 23695 3944 23755
rect 3996 23695 4000 23755
rect 3630 23685 4000 23695
rect 4030 23755 4400 23834
rect 4030 23695 4034 23755
rect 4086 23695 4344 23755
rect 4396 23695 4400 23755
rect 4030 23685 4400 23695
rect 4430 23755 4800 23834
rect 4430 23695 4434 23755
rect 4486 23695 4744 23755
rect 4796 23695 4800 23755
rect 4430 23685 4800 23695
rect 4830 23755 5200 23834
rect 4830 23695 4834 23755
rect 4886 23695 5144 23755
rect 5196 23695 5200 23755
rect 4830 23685 5200 23695
rect 5230 23755 5600 23834
rect 5230 23695 5234 23755
rect 5286 23695 5544 23755
rect 5596 23695 5600 23755
rect 5230 23685 5600 23695
rect 5630 23755 6000 23834
rect 5630 23695 5634 23755
rect 5686 23695 5944 23755
rect 5996 23695 6000 23755
rect 5630 23685 6000 23695
rect 6030 23755 6400 23834
rect 6030 23695 6034 23755
rect 6086 23695 6344 23755
rect 6396 23695 6400 23755
rect 6030 23685 6400 23695
rect 6430 23755 6800 23834
rect 6430 23695 6434 23755
rect 6486 23695 6744 23755
rect 6796 23695 6800 23755
rect 6430 23685 6800 23695
rect 6830 23755 7200 23834
rect 6830 23695 6834 23755
rect 6886 23695 7144 23755
rect 7196 23695 7200 23755
rect 6830 23685 7200 23695
rect 7230 23755 7600 23834
rect 7230 23695 7234 23755
rect 7286 23695 7544 23755
rect 7596 23695 7600 23755
rect 7230 23685 7600 23695
rect 7630 23755 8000 23834
rect 7630 23695 7634 23755
rect 7686 23695 7944 23755
rect 7996 23695 8000 23755
rect 7630 23685 8000 23695
rect 8030 23755 8400 23834
rect 8030 23695 8034 23755
rect 8086 23695 8344 23755
rect 8396 23695 8400 23755
rect 8030 23685 8400 23695
rect 8430 23755 8800 23834
rect 8430 23695 8434 23755
rect 8486 23695 8744 23755
rect 8796 23695 8800 23755
rect 8430 23685 8800 23695
rect 8830 23755 9200 23834
rect 8830 23695 8834 23755
rect 8886 23695 9144 23755
rect 9196 23695 9200 23755
rect 8830 23685 9200 23695
rect 9230 23755 9600 23834
rect 9230 23695 9234 23755
rect 9286 23695 9544 23755
rect 9596 23695 9600 23755
rect 9230 23685 9600 23695
rect 9630 23755 10000 23834
rect 9630 23695 9634 23755
rect 9686 23695 9944 23755
rect 9996 23695 10000 23755
rect 9630 23685 10000 23695
rect 10030 23755 10400 23834
rect 10030 23695 10034 23755
rect 10086 23695 10344 23755
rect 10396 23695 10400 23755
rect 10030 23685 10400 23695
rect 10430 23755 10800 23834
rect 10430 23695 10434 23755
rect 10486 23695 10744 23755
rect 10796 23695 10800 23755
rect 10430 23685 10800 23695
rect 10830 23755 11200 23834
rect 10830 23695 10834 23755
rect 10886 23695 11144 23755
rect 11196 23695 11200 23755
rect 10830 23685 11200 23695
rect 11230 23755 11600 23834
rect 11230 23695 11234 23755
rect 11286 23695 11544 23755
rect 11596 23695 11600 23755
rect 11230 23685 11600 23695
rect 11630 23755 12000 23834
rect 11630 23695 11634 23755
rect 11686 23695 11944 23755
rect 11996 23695 12000 23755
rect 11630 23685 12000 23695
rect 12030 23755 12400 23834
rect 12030 23695 12034 23755
rect 12086 23695 12344 23755
rect 12396 23695 12400 23755
rect 12030 23685 12400 23695
rect 12430 23755 12800 23834
rect 12430 23695 12434 23755
rect 12486 23695 12744 23755
rect 12796 23695 12800 23755
rect 12430 23685 12800 23695
rect 12830 23755 13200 23834
rect 12830 23695 12834 23755
rect 12886 23695 13144 23755
rect 13196 23695 13200 23755
rect 12830 23685 13200 23695
rect -330 23655 -324 23685
rect -330 23645 0 23655
rect -314 23585 -56 23645
rect -4 23585 0 23645
rect -330 23385 0 23585
rect -314 23325 -56 23385
rect -4 23325 0 23385
rect -330 23315 0 23325
rect 30 23645 400 23655
rect 30 23585 34 23645
rect 86 23585 344 23645
rect 396 23585 400 23645
rect 30 23510 400 23585
rect 430 23645 800 23655
rect 430 23585 434 23645
rect 486 23585 744 23645
rect 796 23585 800 23645
rect 430 23510 800 23585
rect 830 23645 1200 23655
rect 830 23585 834 23645
rect 886 23585 1144 23645
rect 1196 23585 1200 23645
rect 830 23510 1200 23585
rect 1230 23645 1600 23655
rect 1230 23585 1234 23645
rect 1286 23585 1544 23645
rect 1596 23585 1600 23645
rect 1230 23510 1600 23585
rect 1630 23645 2000 23655
rect 1630 23585 1634 23645
rect 1686 23585 1944 23645
rect 1996 23585 2000 23645
rect 1630 23510 2000 23585
rect 2030 23645 2400 23655
rect 2030 23585 2034 23645
rect 2086 23585 2344 23645
rect 2396 23585 2400 23645
rect 2030 23510 2400 23585
rect 2430 23645 2800 23655
rect 2430 23585 2434 23645
rect 2486 23585 2744 23645
rect 2796 23585 2800 23645
rect 2430 23510 2800 23585
rect 2830 23645 3200 23655
rect 2830 23585 2834 23645
rect 2886 23585 3144 23645
rect 3196 23585 3200 23645
rect 2830 23510 3200 23585
rect 3230 23645 3600 23655
rect 3230 23585 3234 23645
rect 3286 23585 3544 23645
rect 3596 23585 3600 23645
rect 3230 23510 3600 23585
rect 3630 23645 4000 23655
rect 3630 23585 3634 23645
rect 3686 23585 3944 23645
rect 3996 23585 4000 23645
rect 3630 23510 4000 23585
rect 4030 23645 4400 23655
rect 4030 23585 4034 23645
rect 4086 23585 4344 23645
rect 4396 23585 4400 23645
rect 4030 23510 4400 23585
rect 4430 23645 4800 23655
rect 4430 23585 4434 23645
rect 4486 23585 4744 23645
rect 4796 23585 4800 23645
rect 4430 23510 4800 23585
rect 4830 23645 5200 23655
rect 4830 23585 4834 23645
rect 4886 23585 5144 23645
rect 5196 23585 5200 23645
rect 4830 23510 5200 23585
rect 5230 23645 5600 23655
rect 5230 23585 5234 23645
rect 5286 23585 5544 23645
rect 5596 23585 5600 23645
rect 5230 23510 5600 23585
rect 5630 23645 6000 23655
rect 5630 23585 5634 23645
rect 5686 23585 5944 23645
rect 5996 23585 6000 23645
rect 5630 23510 6000 23585
rect 6030 23645 6400 23655
rect 6030 23585 6034 23645
rect 6086 23585 6344 23645
rect 6396 23585 6400 23645
rect 6030 23510 6400 23585
rect 6430 23645 6800 23655
rect 6430 23585 6434 23645
rect 6486 23585 6744 23645
rect 6796 23585 6800 23645
rect 6430 23510 6800 23585
rect 6830 23645 7200 23655
rect 6830 23585 6834 23645
rect 6886 23585 7144 23645
rect 7196 23585 7200 23645
rect 6830 23510 7200 23585
rect 7230 23645 7600 23655
rect 7230 23585 7234 23645
rect 7286 23585 7544 23645
rect 7596 23585 7600 23645
rect 7230 23510 7600 23585
rect 7630 23645 8000 23655
rect 7630 23585 7634 23645
rect 7686 23585 7944 23645
rect 7996 23585 8000 23645
rect 7630 23510 8000 23585
rect 8030 23645 8400 23655
rect 8030 23585 8034 23645
rect 8086 23585 8344 23645
rect 8396 23585 8400 23645
rect 8030 23510 8400 23585
rect 8430 23645 8800 23655
rect 8430 23585 8434 23645
rect 8486 23585 8744 23645
rect 8796 23585 8800 23645
rect 8430 23510 8800 23585
rect 8830 23645 9200 23655
rect 8830 23585 8834 23645
rect 8886 23585 9144 23645
rect 9196 23585 9200 23645
rect 8830 23510 9200 23585
rect 9230 23645 9600 23655
rect 9230 23585 9234 23645
rect 9286 23585 9544 23645
rect 9596 23585 9600 23645
rect 9230 23510 9600 23585
rect 9630 23645 10000 23655
rect 9630 23585 9634 23645
rect 9686 23585 9944 23645
rect 9996 23585 10000 23645
rect 9630 23510 10000 23585
rect 10030 23645 10400 23655
rect 10030 23585 10034 23645
rect 10086 23585 10344 23645
rect 10396 23585 10400 23645
rect 10030 23510 10400 23585
rect 10430 23645 10800 23655
rect 10430 23585 10434 23645
rect 10486 23585 10744 23645
rect 10796 23585 10800 23645
rect 10430 23510 10800 23585
rect 10830 23645 11200 23655
rect 10830 23585 10834 23645
rect 10886 23585 11144 23645
rect 11196 23585 11200 23645
rect 10830 23510 11200 23585
rect 11230 23645 11600 23655
rect 11230 23585 11234 23645
rect 11286 23585 11544 23645
rect 11596 23585 11600 23645
rect 11230 23510 11600 23585
rect 11630 23645 12000 23655
rect 11630 23585 11634 23645
rect 11686 23585 11944 23645
rect 11996 23585 12000 23645
rect 11630 23510 12000 23585
rect 12030 23645 12400 23655
rect 12030 23585 12034 23645
rect 12086 23585 12344 23645
rect 12396 23585 12400 23645
rect 12030 23510 12400 23585
rect 12430 23645 12800 23655
rect 12430 23585 12434 23645
rect 12486 23585 12744 23645
rect 12796 23585 12800 23645
rect 12430 23510 12800 23585
rect 12830 23645 13200 23655
rect 12830 23585 12834 23645
rect 12886 23585 13144 23645
rect 13196 23585 13200 23645
rect 12830 23510 13200 23585
rect 30 23470 13200 23510
rect 30 23385 400 23470
rect 30 23325 34 23385
rect 86 23325 344 23385
rect 396 23325 400 23385
rect 30 23315 400 23325
rect 430 23385 800 23470
rect 430 23325 434 23385
rect 486 23325 744 23385
rect 796 23325 800 23385
rect 430 23315 800 23325
rect 830 23385 1200 23470
rect 830 23325 834 23385
rect 886 23325 1144 23385
rect 1196 23325 1200 23385
rect 830 23315 1200 23325
rect 1230 23385 1600 23470
rect 1230 23325 1234 23385
rect 1286 23325 1544 23385
rect 1596 23325 1600 23385
rect 1230 23315 1600 23325
rect 1630 23385 2000 23470
rect 1630 23325 1634 23385
rect 1686 23325 1944 23385
rect 1996 23325 2000 23385
rect 1630 23315 2000 23325
rect 2030 23385 2400 23470
rect 2030 23325 2034 23385
rect 2086 23325 2344 23385
rect 2396 23325 2400 23385
rect 2030 23315 2400 23325
rect 2430 23385 2800 23470
rect 2430 23325 2434 23385
rect 2486 23325 2744 23385
rect 2796 23325 2800 23385
rect 2430 23315 2800 23325
rect 2830 23385 3200 23470
rect 2830 23325 2834 23385
rect 2886 23325 3144 23385
rect 3196 23325 3200 23385
rect 2830 23315 3200 23325
rect 3230 23385 3600 23470
rect 3230 23325 3234 23385
rect 3286 23325 3544 23385
rect 3596 23325 3600 23385
rect 3230 23315 3600 23325
rect 3630 23385 4000 23470
rect 3630 23325 3634 23385
rect 3686 23325 3944 23385
rect 3996 23325 4000 23385
rect 3630 23315 4000 23325
rect 4030 23385 4400 23470
rect 4030 23325 4034 23385
rect 4086 23325 4344 23385
rect 4396 23325 4400 23385
rect 4030 23315 4400 23325
rect 4430 23385 4800 23470
rect 4430 23325 4434 23385
rect 4486 23325 4744 23385
rect 4796 23325 4800 23385
rect 4430 23315 4800 23325
rect 4830 23385 5200 23470
rect 4830 23325 4834 23385
rect 4886 23325 5144 23385
rect 5196 23325 5200 23385
rect 4830 23315 5200 23325
rect 5230 23385 5600 23470
rect 5230 23325 5234 23385
rect 5286 23325 5544 23385
rect 5596 23325 5600 23385
rect 5230 23315 5600 23325
rect 5630 23385 6000 23470
rect 5630 23325 5634 23385
rect 5686 23325 5944 23385
rect 5996 23325 6000 23385
rect 5630 23315 6000 23325
rect 6030 23385 6400 23470
rect 6030 23325 6034 23385
rect 6086 23325 6344 23385
rect 6396 23325 6400 23385
rect 6030 23315 6400 23325
rect 6430 23385 6800 23470
rect 6430 23325 6434 23385
rect 6486 23325 6744 23385
rect 6796 23325 6800 23385
rect 6430 23315 6800 23325
rect 6830 23385 7200 23470
rect 6830 23325 6834 23385
rect 6886 23325 7144 23385
rect 7196 23325 7200 23385
rect 6830 23315 7200 23325
rect 7230 23385 7600 23470
rect 7230 23325 7234 23385
rect 7286 23325 7544 23385
rect 7596 23325 7600 23385
rect 7230 23315 7600 23325
rect 7630 23385 8000 23470
rect 7630 23325 7634 23385
rect 7686 23325 7944 23385
rect 7996 23325 8000 23385
rect 7630 23315 8000 23325
rect 8030 23385 8400 23470
rect 8030 23325 8034 23385
rect 8086 23325 8344 23385
rect 8396 23325 8400 23385
rect 8030 23315 8400 23325
rect 8430 23385 8800 23470
rect 8430 23325 8434 23385
rect 8486 23325 8744 23385
rect 8796 23325 8800 23385
rect 8430 23315 8800 23325
rect 8830 23385 9200 23470
rect 8830 23325 8834 23385
rect 8886 23325 9144 23385
rect 9196 23325 9200 23385
rect 8830 23315 9200 23325
rect 9230 23385 9600 23470
rect 9230 23325 9234 23385
rect 9286 23325 9544 23385
rect 9596 23325 9600 23385
rect 9230 23315 9600 23325
rect 9630 23385 10000 23470
rect 9630 23325 9634 23385
rect 9686 23325 9944 23385
rect 9996 23325 10000 23385
rect 9630 23315 10000 23325
rect 10030 23385 10400 23470
rect 10030 23325 10034 23385
rect 10086 23325 10344 23385
rect 10396 23325 10400 23385
rect 10030 23315 10400 23325
rect 10430 23385 10800 23470
rect 10430 23325 10434 23385
rect 10486 23325 10744 23385
rect 10796 23325 10800 23385
rect 10430 23315 10800 23325
rect 10830 23385 11200 23470
rect 10830 23325 10834 23385
rect 10886 23325 11144 23385
rect 11196 23325 11200 23385
rect 10830 23315 11200 23325
rect 11230 23385 11600 23470
rect 11230 23325 11234 23385
rect 11286 23325 11544 23385
rect 11596 23325 11600 23385
rect 11230 23315 11600 23325
rect 11630 23385 12000 23470
rect 11630 23325 11634 23385
rect 11686 23325 11944 23385
rect 11996 23325 12000 23385
rect 11630 23315 12000 23325
rect 12030 23385 12400 23470
rect 12030 23325 12034 23385
rect 12086 23325 12344 23385
rect 12396 23325 12400 23385
rect 12030 23315 12400 23325
rect 12430 23385 12800 23470
rect 12430 23325 12434 23385
rect 12486 23325 12744 23385
rect 12796 23325 12800 23385
rect 12430 23315 12800 23325
rect 12830 23385 13200 23470
rect 12830 23325 12834 23385
rect 12886 23325 13144 23385
rect 13196 23325 13200 23385
rect 12830 23315 13200 23325
rect -330 23285 -324 23315
rect 30 23285 70 23315
rect 430 23285 470 23315
rect 830 23285 870 23315
rect 1230 23285 1270 23315
rect 1630 23285 1670 23315
rect 2030 23285 2070 23315
rect 2430 23285 2470 23315
rect 2830 23285 2870 23315
rect 3230 23285 3270 23315
rect 3630 23285 3670 23315
rect 4030 23285 4070 23315
rect 4430 23285 4470 23315
rect 4830 23285 4870 23315
rect 5230 23285 5270 23315
rect 5630 23285 5670 23315
rect 6030 23285 6070 23315
rect 6430 23285 6470 23315
rect 6830 23285 6870 23315
rect 7230 23285 7270 23315
rect 7630 23285 7670 23315
rect 8030 23285 8070 23315
rect 8430 23285 8470 23315
rect 8830 23285 8870 23315
rect 9230 23285 9270 23315
rect 9630 23285 9670 23315
rect 10030 23285 10070 23315
rect 10430 23285 10470 23315
rect 10830 23285 10870 23315
rect 11230 23285 11270 23315
rect 11630 23285 11670 23315
rect 12030 23285 12070 23315
rect 12430 23285 12470 23315
rect -330 23275 0 23285
rect -314 23215 -56 23275
rect -4 23215 0 23275
rect -330 23015 0 23215
rect -314 22955 -56 23015
rect -4 22955 0 23015
rect -330 22945 0 22955
rect 30 23275 400 23285
rect 30 23215 34 23275
rect 86 23215 344 23275
rect 396 23215 400 23275
rect 30 23140 400 23215
rect 430 23275 800 23285
rect 430 23215 434 23275
rect 486 23215 744 23275
rect 796 23215 800 23275
rect 430 23140 800 23215
rect 830 23275 1200 23285
rect 830 23215 834 23275
rect 886 23215 1144 23275
rect 1196 23215 1200 23275
rect 830 23140 1200 23215
rect 1230 23275 1600 23285
rect 1230 23215 1234 23275
rect 1286 23215 1544 23275
rect 1596 23215 1600 23275
rect 1230 23140 1600 23215
rect 1630 23275 2000 23285
rect 1630 23215 1634 23275
rect 1686 23215 1944 23275
rect 1996 23215 2000 23275
rect 1630 23140 2000 23215
rect 2030 23275 2400 23285
rect 2030 23215 2034 23275
rect 2086 23215 2344 23275
rect 2396 23215 2400 23275
rect 2030 23140 2400 23215
rect 2430 23275 2800 23285
rect 2430 23215 2434 23275
rect 2486 23215 2744 23275
rect 2796 23215 2800 23275
rect 2430 23140 2800 23215
rect 2830 23275 3200 23285
rect 2830 23215 2834 23275
rect 2886 23215 3144 23275
rect 3196 23215 3200 23275
rect 2830 23140 3200 23215
rect 3230 23275 3600 23285
rect 3230 23215 3234 23275
rect 3286 23215 3544 23275
rect 3596 23215 3600 23275
rect 3230 23140 3600 23215
rect 3630 23275 4000 23285
rect 3630 23215 3634 23275
rect 3686 23215 3944 23275
rect 3996 23215 4000 23275
rect 3630 23140 4000 23215
rect 4030 23275 4400 23285
rect 4030 23215 4034 23275
rect 4086 23215 4344 23275
rect 4396 23215 4400 23275
rect 4030 23140 4400 23215
rect 4430 23275 4800 23285
rect 4430 23215 4434 23275
rect 4486 23215 4744 23275
rect 4796 23215 4800 23275
rect 4430 23140 4800 23215
rect 4830 23275 5200 23285
rect 4830 23215 4834 23275
rect 4886 23215 5144 23275
rect 5196 23215 5200 23275
rect 4830 23140 5200 23215
rect 5230 23275 5600 23285
rect 5230 23215 5234 23275
rect 5286 23215 5544 23275
rect 5596 23215 5600 23275
rect 5230 23140 5600 23215
rect 5630 23275 6000 23285
rect 5630 23215 5634 23275
rect 5686 23215 5944 23275
rect 5996 23215 6000 23275
rect 5630 23140 6000 23215
rect 6030 23275 6400 23285
rect 6030 23215 6034 23275
rect 6086 23215 6344 23275
rect 6396 23215 6400 23275
rect 6030 23140 6400 23215
rect 6430 23275 6800 23285
rect 6430 23215 6434 23275
rect 6486 23215 6744 23275
rect 6796 23215 6800 23275
rect 6430 23140 6800 23215
rect 6830 23275 7200 23285
rect 6830 23215 6834 23275
rect 6886 23215 7144 23275
rect 7196 23215 7200 23275
rect 6830 23140 7200 23215
rect 7230 23275 7600 23285
rect 7230 23215 7234 23275
rect 7286 23215 7544 23275
rect 7596 23215 7600 23275
rect 7230 23140 7600 23215
rect 7630 23275 8000 23285
rect 7630 23215 7634 23275
rect 7686 23215 7944 23275
rect 7996 23215 8000 23275
rect 7630 23140 8000 23215
rect 8030 23275 8400 23285
rect 8030 23215 8034 23275
rect 8086 23215 8344 23275
rect 8396 23215 8400 23275
rect 8030 23140 8400 23215
rect 8430 23275 8800 23285
rect 8430 23215 8434 23275
rect 8486 23215 8744 23275
rect 8796 23215 8800 23275
rect 8430 23140 8800 23215
rect 8830 23275 9200 23285
rect 8830 23215 8834 23275
rect 8886 23215 9144 23275
rect 9196 23215 9200 23275
rect 8830 23140 9200 23215
rect 9230 23275 9600 23285
rect 9230 23215 9234 23275
rect 9286 23215 9544 23275
rect 9596 23215 9600 23275
rect 9230 23140 9600 23215
rect 9630 23275 10000 23285
rect 9630 23215 9634 23275
rect 9686 23215 9944 23275
rect 9996 23215 10000 23275
rect 9630 23140 10000 23215
rect 10030 23275 10400 23285
rect 10030 23215 10034 23275
rect 10086 23215 10344 23275
rect 10396 23215 10400 23275
rect 10030 23140 10400 23215
rect 10430 23275 10800 23285
rect 10430 23215 10434 23275
rect 10486 23215 10744 23275
rect 10796 23215 10800 23275
rect 10430 23140 10800 23215
rect 10830 23275 11200 23285
rect 10830 23215 10834 23275
rect 10886 23215 11144 23275
rect 11196 23215 11200 23275
rect 10830 23140 11200 23215
rect 11230 23275 11600 23285
rect 11230 23215 11234 23275
rect 11286 23215 11544 23275
rect 11596 23215 11600 23275
rect 11230 23140 11600 23215
rect 11630 23275 12000 23285
rect 11630 23215 11634 23275
rect 11686 23215 11944 23275
rect 11996 23215 12000 23275
rect 11630 23140 12000 23215
rect 12030 23275 12400 23285
rect 12030 23215 12034 23275
rect 12086 23215 12344 23275
rect 12396 23215 12400 23275
rect 12030 23140 12400 23215
rect 12430 23275 12800 23285
rect 12430 23215 12434 23275
rect 12486 23215 12744 23275
rect 12796 23215 12800 23275
rect 12430 23140 12800 23215
rect 12830 23275 13200 23285
rect 12830 23215 12834 23275
rect 12886 23215 13144 23275
rect 13196 23215 13200 23275
rect 12830 23140 13200 23215
rect 30 23100 13200 23140
rect 30 23015 400 23100
rect 30 22955 34 23015
rect 86 22955 344 23015
rect 396 22955 400 23015
rect 30 22945 400 22955
rect 430 23015 800 23100
rect 430 22955 434 23015
rect 486 22955 744 23015
rect 796 22955 800 23015
rect 430 22945 800 22955
rect 830 23015 1200 23100
rect 830 22955 834 23015
rect 886 22955 1144 23015
rect 1196 22955 1200 23015
rect 830 22945 1200 22955
rect 1230 23015 1600 23100
rect 1230 22955 1234 23015
rect 1286 22955 1544 23015
rect 1596 22955 1600 23015
rect 1230 22945 1600 22955
rect 1630 23015 2000 23100
rect 1630 22955 1634 23015
rect 1686 22955 1944 23015
rect 1996 22955 2000 23015
rect 1630 22945 2000 22955
rect 2030 23015 2400 23100
rect 2030 22955 2034 23015
rect 2086 22955 2344 23015
rect 2396 22955 2400 23015
rect 2030 22945 2400 22955
rect 2430 23015 2800 23100
rect 2430 22955 2434 23015
rect 2486 22955 2744 23015
rect 2796 22955 2800 23015
rect 2430 22945 2800 22955
rect 2830 23015 3200 23100
rect 2830 22955 2834 23015
rect 2886 22955 3144 23015
rect 3196 22955 3200 23015
rect 2830 22945 3200 22955
rect 3230 23015 3600 23100
rect 3230 22955 3234 23015
rect 3286 22955 3544 23015
rect 3596 22955 3600 23015
rect 3230 22945 3600 22955
rect 3630 23015 4000 23100
rect 3630 22955 3634 23015
rect 3686 22955 3944 23015
rect 3996 22955 4000 23015
rect 3630 22945 4000 22955
rect 4030 23015 4400 23100
rect 4030 22955 4034 23015
rect 4086 22955 4344 23015
rect 4396 22955 4400 23015
rect 4030 22945 4400 22955
rect 4430 23015 4800 23100
rect 4430 22955 4434 23015
rect 4486 22955 4744 23015
rect 4796 22955 4800 23015
rect 4430 22945 4800 22955
rect 4830 23015 5200 23100
rect 4830 22955 4834 23015
rect 4886 22955 5144 23015
rect 5196 22955 5200 23015
rect 4830 22945 5200 22955
rect 5230 23015 5600 23100
rect 5230 22955 5234 23015
rect 5286 22955 5544 23015
rect 5596 22955 5600 23015
rect 5230 22945 5600 22955
rect 5630 23015 6000 23100
rect 5630 22955 5634 23015
rect 5686 22955 5944 23015
rect 5996 22955 6000 23015
rect 5630 22945 6000 22955
rect 6030 23015 6400 23100
rect 6030 22955 6034 23015
rect 6086 22955 6344 23015
rect 6396 22955 6400 23015
rect 6030 22945 6400 22955
rect 6430 23015 6800 23100
rect 6430 22955 6434 23015
rect 6486 22955 6744 23015
rect 6796 22955 6800 23015
rect 6430 22945 6800 22955
rect 6830 23015 7200 23100
rect 6830 22955 6834 23015
rect 6886 22955 7144 23015
rect 7196 22955 7200 23015
rect 6830 22945 7200 22955
rect 7230 23015 7600 23100
rect 7230 22955 7234 23015
rect 7286 22955 7544 23015
rect 7596 22955 7600 23015
rect 7230 22945 7600 22955
rect 7630 23015 8000 23100
rect 7630 22955 7634 23015
rect 7686 22955 7944 23015
rect 7996 22955 8000 23015
rect 7630 22945 8000 22955
rect 8030 23015 8400 23100
rect 8030 22955 8034 23015
rect 8086 22955 8344 23015
rect 8396 22955 8400 23015
rect 8030 22945 8400 22955
rect 8430 23015 8800 23100
rect 8430 22955 8434 23015
rect 8486 22955 8744 23015
rect 8796 22955 8800 23015
rect 8430 22945 8800 22955
rect 8830 23015 9200 23100
rect 8830 22955 8834 23015
rect 8886 22955 9144 23015
rect 9196 22955 9200 23015
rect 8830 22945 9200 22955
rect 9230 23015 9600 23100
rect 9230 22955 9234 23015
rect 9286 22955 9544 23015
rect 9596 22955 9600 23015
rect 9230 22945 9600 22955
rect 9630 23015 10000 23100
rect 9630 22955 9634 23015
rect 9686 22955 9944 23015
rect 9996 22955 10000 23015
rect 9630 22945 10000 22955
rect 10030 23015 10400 23100
rect 10030 22955 10034 23015
rect 10086 22955 10344 23015
rect 10396 22955 10400 23015
rect 10030 22945 10400 22955
rect 10430 23015 10800 23100
rect 10430 22955 10434 23015
rect 10486 22955 10744 23015
rect 10796 22955 10800 23015
rect 10430 22945 10800 22955
rect 10830 23015 11200 23100
rect 10830 22955 10834 23015
rect 10886 22955 11144 23015
rect 11196 22955 11200 23015
rect 10830 22945 11200 22955
rect 11230 23015 11600 23100
rect 11230 22955 11234 23015
rect 11286 22955 11544 23015
rect 11596 22955 11600 23015
rect 11230 22945 11600 22955
rect 11630 23015 12000 23100
rect 11630 22955 11634 23015
rect 11686 22955 11944 23015
rect 11996 22955 12000 23015
rect 11630 22945 12000 22955
rect 12030 23015 12400 23100
rect 12030 22955 12034 23015
rect 12086 22955 12344 23015
rect 12396 22955 12400 23015
rect 12030 22945 12400 22955
rect 12430 23015 12800 23100
rect 12430 22955 12434 23015
rect 12486 22955 12744 23015
rect 12796 22955 12800 23015
rect 12430 22945 12800 22955
rect 12830 23015 13200 23100
rect 12830 22955 12834 23015
rect 12886 22955 13144 23015
rect 13196 22955 13200 23015
rect 12830 22945 13200 22955
rect -330 22915 -324 22945
rect 30 22915 70 22945
rect 430 22915 470 22945
rect 830 22915 870 22945
rect 1230 22915 1270 22945
rect 1630 22915 1670 22945
rect 2030 22915 2070 22945
rect 2430 22915 2470 22945
rect 2830 22915 2870 22945
rect 3230 22915 3270 22945
rect 3630 22915 3670 22945
rect 4030 22915 4070 22945
rect 4430 22915 4470 22945
rect 4830 22915 4870 22945
rect 5230 22915 5270 22945
rect 5630 22915 5670 22945
rect 6030 22915 6070 22945
rect 6430 22915 6470 22945
rect 6830 22915 6870 22945
rect 7230 22915 7270 22945
rect 7630 22915 7670 22945
rect 8030 22915 8070 22945
rect 8430 22915 8470 22945
rect 8830 22915 8870 22945
rect 9230 22915 9270 22945
rect 9630 22915 9670 22945
rect 10030 22915 10070 22945
rect 10430 22915 10470 22945
rect 10830 22915 10870 22945
rect 11230 22915 11270 22945
rect 11630 22915 11670 22945
rect 12030 22915 12070 22945
rect 12430 22915 12470 22945
rect -330 22905 0 22915
rect -314 22845 -56 22905
rect -4 22845 0 22905
rect -330 22645 0 22845
rect -314 22585 -56 22645
rect -4 22585 0 22645
rect -330 22575 0 22585
rect 30 22905 400 22915
rect 30 22845 34 22905
rect 86 22845 344 22905
rect 396 22845 400 22905
rect 30 22770 400 22845
rect 430 22905 800 22915
rect 430 22845 434 22905
rect 486 22845 744 22905
rect 796 22845 800 22905
rect 430 22770 800 22845
rect 830 22905 1200 22915
rect 830 22845 834 22905
rect 886 22845 1144 22905
rect 1196 22845 1200 22905
rect 830 22770 1200 22845
rect 1230 22905 1600 22915
rect 1230 22845 1234 22905
rect 1286 22845 1544 22905
rect 1596 22845 1600 22905
rect 1230 22770 1600 22845
rect 1630 22905 2000 22915
rect 1630 22845 1634 22905
rect 1686 22845 1944 22905
rect 1996 22845 2000 22905
rect 1630 22770 2000 22845
rect 2030 22905 2400 22915
rect 2030 22845 2034 22905
rect 2086 22845 2344 22905
rect 2396 22845 2400 22905
rect 2030 22770 2400 22845
rect 2430 22905 2800 22915
rect 2430 22845 2434 22905
rect 2486 22845 2744 22905
rect 2796 22845 2800 22905
rect 2430 22770 2800 22845
rect 2830 22905 3200 22915
rect 2830 22845 2834 22905
rect 2886 22845 3144 22905
rect 3196 22845 3200 22905
rect 2830 22770 3200 22845
rect 3230 22905 3600 22915
rect 3230 22845 3234 22905
rect 3286 22845 3544 22905
rect 3596 22845 3600 22905
rect 3230 22770 3600 22845
rect 3630 22905 4000 22915
rect 3630 22845 3634 22905
rect 3686 22845 3944 22905
rect 3996 22845 4000 22905
rect 3630 22770 4000 22845
rect 4030 22905 4400 22915
rect 4030 22845 4034 22905
rect 4086 22845 4344 22905
rect 4396 22845 4400 22905
rect 4030 22770 4400 22845
rect 4430 22905 4800 22915
rect 4430 22845 4434 22905
rect 4486 22845 4744 22905
rect 4796 22845 4800 22905
rect 4430 22770 4800 22845
rect 4830 22905 5200 22915
rect 4830 22845 4834 22905
rect 4886 22845 5144 22905
rect 5196 22845 5200 22905
rect 4830 22770 5200 22845
rect 5230 22905 5600 22915
rect 5230 22845 5234 22905
rect 5286 22845 5544 22905
rect 5596 22845 5600 22905
rect 5230 22770 5600 22845
rect 5630 22905 6000 22915
rect 5630 22845 5634 22905
rect 5686 22845 5944 22905
rect 5996 22845 6000 22905
rect 5630 22770 6000 22845
rect 6030 22905 6400 22915
rect 6030 22845 6034 22905
rect 6086 22845 6344 22905
rect 6396 22845 6400 22905
rect 6030 22770 6400 22845
rect 6430 22905 6800 22915
rect 6430 22845 6434 22905
rect 6486 22845 6744 22905
rect 6796 22845 6800 22905
rect 6430 22770 6800 22845
rect 6830 22905 7200 22915
rect 6830 22845 6834 22905
rect 6886 22845 7144 22905
rect 7196 22845 7200 22905
rect 6830 22770 7200 22845
rect 7230 22905 7600 22915
rect 7230 22845 7234 22905
rect 7286 22845 7544 22905
rect 7596 22845 7600 22905
rect 7230 22770 7600 22845
rect 7630 22905 8000 22915
rect 7630 22845 7634 22905
rect 7686 22845 7944 22905
rect 7996 22845 8000 22905
rect 7630 22770 8000 22845
rect 8030 22905 8400 22915
rect 8030 22845 8034 22905
rect 8086 22845 8344 22905
rect 8396 22845 8400 22905
rect 8030 22770 8400 22845
rect 8430 22905 8800 22915
rect 8430 22845 8434 22905
rect 8486 22845 8744 22905
rect 8796 22845 8800 22905
rect 8430 22770 8800 22845
rect 8830 22905 9200 22915
rect 8830 22845 8834 22905
rect 8886 22845 9144 22905
rect 9196 22845 9200 22905
rect 8830 22770 9200 22845
rect 9230 22905 9600 22915
rect 9230 22845 9234 22905
rect 9286 22845 9544 22905
rect 9596 22845 9600 22905
rect 9230 22770 9600 22845
rect 9630 22905 10000 22915
rect 9630 22845 9634 22905
rect 9686 22845 9944 22905
rect 9996 22845 10000 22905
rect 9630 22770 10000 22845
rect 10030 22905 10400 22915
rect 10030 22845 10034 22905
rect 10086 22845 10344 22905
rect 10396 22845 10400 22905
rect 10030 22770 10400 22845
rect 10430 22905 10800 22915
rect 10430 22845 10434 22905
rect 10486 22845 10744 22905
rect 10796 22845 10800 22905
rect 10430 22770 10800 22845
rect 10830 22905 11200 22915
rect 10830 22845 10834 22905
rect 10886 22845 11144 22905
rect 11196 22845 11200 22905
rect 10830 22770 11200 22845
rect 11230 22905 11600 22915
rect 11230 22845 11234 22905
rect 11286 22845 11544 22905
rect 11596 22845 11600 22905
rect 11230 22770 11600 22845
rect 11630 22905 12000 22915
rect 11630 22845 11634 22905
rect 11686 22845 11944 22905
rect 11996 22845 12000 22905
rect 11630 22770 12000 22845
rect 12030 22905 12400 22915
rect 12030 22845 12034 22905
rect 12086 22845 12344 22905
rect 12396 22845 12400 22905
rect 12030 22770 12400 22845
rect 12430 22905 12800 22915
rect 12430 22845 12434 22905
rect 12486 22845 12744 22905
rect 12796 22845 12800 22905
rect 12430 22770 12800 22845
rect 12830 22905 13200 22915
rect 12830 22845 12834 22905
rect 12886 22845 13144 22905
rect 13196 22845 13200 22905
rect 12830 22770 13200 22845
rect 30 22730 13200 22770
rect 30 22645 400 22730
rect 30 22585 34 22645
rect 86 22585 344 22645
rect 396 22585 400 22645
rect 30 22575 400 22585
rect 430 22645 800 22730
rect 430 22585 434 22645
rect 486 22585 744 22645
rect 796 22585 800 22645
rect 430 22575 800 22585
rect 830 22645 1200 22730
rect 830 22585 834 22645
rect 886 22585 1144 22645
rect 1196 22585 1200 22645
rect 830 22575 1200 22585
rect 1230 22645 1600 22730
rect 1230 22585 1234 22645
rect 1286 22585 1544 22645
rect 1596 22585 1600 22645
rect 1230 22575 1600 22585
rect 1630 22645 2000 22730
rect 1630 22585 1634 22645
rect 1686 22585 1944 22645
rect 1996 22585 2000 22645
rect 1630 22575 2000 22585
rect 2030 22645 2400 22730
rect 2030 22585 2034 22645
rect 2086 22585 2344 22645
rect 2396 22585 2400 22645
rect 2030 22575 2400 22585
rect 2430 22645 2800 22730
rect 2430 22585 2434 22645
rect 2486 22585 2744 22645
rect 2796 22585 2800 22645
rect 2430 22575 2800 22585
rect 2830 22645 3200 22730
rect 2830 22585 2834 22645
rect 2886 22585 3144 22645
rect 3196 22585 3200 22645
rect 2830 22575 3200 22585
rect 3230 22645 3600 22730
rect 3230 22585 3234 22645
rect 3286 22585 3544 22645
rect 3596 22585 3600 22645
rect 3230 22575 3600 22585
rect 3630 22645 4000 22730
rect 3630 22585 3634 22645
rect 3686 22585 3944 22645
rect 3996 22585 4000 22645
rect 3630 22575 4000 22585
rect 4030 22645 4400 22730
rect 4030 22585 4034 22645
rect 4086 22585 4344 22645
rect 4396 22585 4400 22645
rect 4030 22575 4400 22585
rect 4430 22645 4800 22730
rect 4430 22585 4434 22645
rect 4486 22585 4744 22645
rect 4796 22585 4800 22645
rect 4430 22575 4800 22585
rect 4830 22645 5200 22730
rect 4830 22585 4834 22645
rect 4886 22585 5144 22645
rect 5196 22585 5200 22645
rect 4830 22575 5200 22585
rect 5230 22645 5600 22730
rect 5230 22585 5234 22645
rect 5286 22585 5544 22645
rect 5596 22585 5600 22645
rect 5230 22575 5600 22585
rect 5630 22645 6000 22730
rect 5630 22585 5634 22645
rect 5686 22585 5944 22645
rect 5996 22585 6000 22645
rect 5630 22575 6000 22585
rect 6030 22645 6400 22730
rect 6030 22585 6034 22645
rect 6086 22585 6344 22645
rect 6396 22585 6400 22645
rect 6030 22575 6400 22585
rect 6430 22645 6800 22730
rect 6430 22585 6434 22645
rect 6486 22585 6744 22645
rect 6796 22585 6800 22645
rect 6430 22575 6800 22585
rect 6830 22645 7200 22730
rect 6830 22585 6834 22645
rect 6886 22585 7144 22645
rect 7196 22585 7200 22645
rect 6830 22575 7200 22585
rect 7230 22645 7600 22730
rect 7230 22585 7234 22645
rect 7286 22585 7544 22645
rect 7596 22585 7600 22645
rect 7230 22575 7600 22585
rect 7630 22645 8000 22730
rect 7630 22585 7634 22645
rect 7686 22585 7944 22645
rect 7996 22585 8000 22645
rect 7630 22575 8000 22585
rect 8030 22645 8400 22730
rect 8030 22585 8034 22645
rect 8086 22585 8344 22645
rect 8396 22585 8400 22645
rect 8030 22575 8400 22585
rect 8430 22645 8800 22730
rect 8430 22585 8434 22645
rect 8486 22585 8744 22645
rect 8796 22585 8800 22645
rect 8430 22575 8800 22585
rect 8830 22645 9200 22730
rect 8830 22585 8834 22645
rect 8886 22585 9144 22645
rect 9196 22585 9200 22645
rect 8830 22575 9200 22585
rect 9230 22645 9600 22730
rect 9230 22585 9234 22645
rect 9286 22585 9544 22645
rect 9596 22585 9600 22645
rect 9230 22575 9600 22585
rect 9630 22645 10000 22730
rect 9630 22585 9634 22645
rect 9686 22585 9944 22645
rect 9996 22585 10000 22645
rect 9630 22575 10000 22585
rect 10030 22645 10400 22730
rect 10030 22585 10034 22645
rect 10086 22585 10344 22645
rect 10396 22585 10400 22645
rect 10030 22575 10400 22585
rect 10430 22645 10800 22730
rect 10430 22585 10434 22645
rect 10486 22585 10744 22645
rect 10796 22585 10800 22645
rect 10430 22575 10800 22585
rect 10830 22645 11200 22730
rect 10830 22585 10834 22645
rect 10886 22585 11144 22645
rect 11196 22585 11200 22645
rect 10830 22575 11200 22585
rect 11230 22645 11600 22730
rect 11230 22585 11234 22645
rect 11286 22585 11544 22645
rect 11596 22585 11600 22645
rect 11230 22575 11600 22585
rect 11630 22645 12000 22730
rect 11630 22585 11634 22645
rect 11686 22585 11944 22645
rect 11996 22585 12000 22645
rect 11630 22575 12000 22585
rect 12030 22645 12400 22730
rect 12030 22585 12034 22645
rect 12086 22585 12344 22645
rect 12396 22585 12400 22645
rect 12030 22575 12400 22585
rect 12430 22645 12800 22730
rect 12430 22585 12434 22645
rect 12486 22585 12744 22645
rect 12796 22585 12800 22645
rect 12430 22575 12800 22585
rect 12830 22645 13200 22730
rect 12830 22585 12834 22645
rect 12886 22585 13144 22645
rect 13196 22585 13200 22645
rect 12830 22575 13200 22585
rect -330 22545 -324 22575
rect 30 22545 70 22575
rect 430 22545 470 22575
rect 830 22545 870 22575
rect 1230 22545 1270 22575
rect 1630 22545 1670 22575
rect 2030 22545 2070 22575
rect 2430 22545 2470 22575
rect 2830 22545 2870 22575
rect 3230 22545 3270 22575
rect 3630 22545 3670 22575
rect 4030 22545 4070 22575
rect 4430 22545 4470 22575
rect 4830 22545 4870 22575
rect 5230 22545 5270 22575
rect 5630 22545 5670 22575
rect 6030 22545 6070 22575
rect 6430 22545 6470 22575
rect 6830 22545 6870 22575
rect 7230 22545 7270 22575
rect 7630 22545 7670 22575
rect 8030 22545 8070 22575
rect 8430 22545 8470 22575
rect 8830 22545 8870 22575
rect 9230 22545 9270 22575
rect 9630 22545 9670 22575
rect 10030 22545 10070 22575
rect 10430 22545 10470 22575
rect 10830 22545 10870 22575
rect 11230 22545 11270 22575
rect 11630 22545 11670 22575
rect 12030 22545 12070 22575
rect 12430 22545 12470 22575
rect -330 22535 0 22545
rect -314 22475 -56 22535
rect -4 22475 0 22535
rect -330 22275 0 22475
rect -314 22215 -56 22275
rect -4 22215 0 22275
rect -330 22205 0 22215
rect 30 22535 400 22545
rect 30 22475 34 22535
rect 86 22475 344 22535
rect 396 22475 400 22535
rect 30 22400 400 22475
rect 430 22535 800 22545
rect 430 22475 434 22535
rect 486 22475 744 22535
rect 796 22475 800 22535
rect 430 22400 800 22475
rect 830 22535 1200 22545
rect 830 22475 834 22535
rect 886 22475 1144 22535
rect 1196 22475 1200 22535
rect 830 22400 1200 22475
rect 1230 22535 1600 22545
rect 1230 22475 1234 22535
rect 1286 22475 1544 22535
rect 1596 22475 1600 22535
rect 1230 22400 1600 22475
rect 1630 22535 2000 22545
rect 1630 22475 1634 22535
rect 1686 22475 1944 22535
rect 1996 22475 2000 22535
rect 1630 22400 2000 22475
rect 2030 22535 2400 22545
rect 2030 22475 2034 22535
rect 2086 22475 2344 22535
rect 2396 22475 2400 22535
rect 2030 22400 2400 22475
rect 2430 22535 2800 22545
rect 2430 22475 2434 22535
rect 2486 22475 2744 22535
rect 2796 22475 2800 22535
rect 2430 22400 2800 22475
rect 2830 22535 3200 22545
rect 2830 22475 2834 22535
rect 2886 22475 3144 22535
rect 3196 22475 3200 22535
rect 2830 22400 3200 22475
rect 3230 22535 3600 22545
rect 3230 22475 3234 22535
rect 3286 22475 3544 22535
rect 3596 22475 3600 22535
rect 3230 22400 3600 22475
rect 3630 22535 4000 22545
rect 3630 22475 3634 22535
rect 3686 22475 3944 22535
rect 3996 22475 4000 22535
rect 3630 22400 4000 22475
rect 4030 22535 4400 22545
rect 4030 22475 4034 22535
rect 4086 22475 4344 22535
rect 4396 22475 4400 22535
rect 4030 22400 4400 22475
rect 4430 22535 4800 22545
rect 4430 22475 4434 22535
rect 4486 22475 4744 22535
rect 4796 22475 4800 22535
rect 4430 22400 4800 22475
rect 4830 22535 5200 22545
rect 4830 22475 4834 22535
rect 4886 22475 5144 22535
rect 5196 22475 5200 22535
rect 4830 22400 5200 22475
rect 5230 22535 5600 22545
rect 5230 22475 5234 22535
rect 5286 22475 5544 22535
rect 5596 22475 5600 22535
rect 5230 22400 5600 22475
rect 5630 22535 6000 22545
rect 5630 22475 5634 22535
rect 5686 22475 5944 22535
rect 5996 22475 6000 22535
rect 5630 22400 6000 22475
rect 6030 22535 6400 22545
rect 6030 22475 6034 22535
rect 6086 22475 6344 22535
rect 6396 22475 6400 22535
rect 6030 22400 6400 22475
rect 6430 22535 6800 22545
rect 6430 22475 6434 22535
rect 6486 22475 6744 22535
rect 6796 22475 6800 22535
rect 6430 22400 6800 22475
rect 6830 22535 7200 22545
rect 6830 22475 6834 22535
rect 6886 22475 7144 22535
rect 7196 22475 7200 22535
rect 6830 22400 7200 22475
rect 7230 22535 7600 22545
rect 7230 22475 7234 22535
rect 7286 22475 7544 22535
rect 7596 22475 7600 22535
rect 7230 22400 7600 22475
rect 7630 22535 8000 22545
rect 7630 22475 7634 22535
rect 7686 22475 7944 22535
rect 7996 22475 8000 22535
rect 7630 22400 8000 22475
rect 8030 22535 8400 22545
rect 8030 22475 8034 22535
rect 8086 22475 8344 22535
rect 8396 22475 8400 22535
rect 8030 22400 8400 22475
rect 8430 22535 8800 22545
rect 8430 22475 8434 22535
rect 8486 22475 8744 22535
rect 8796 22475 8800 22535
rect 8430 22400 8800 22475
rect 8830 22535 9200 22545
rect 8830 22475 8834 22535
rect 8886 22475 9144 22535
rect 9196 22475 9200 22535
rect 8830 22400 9200 22475
rect 9230 22535 9600 22545
rect 9230 22475 9234 22535
rect 9286 22475 9544 22535
rect 9596 22475 9600 22535
rect 9230 22400 9600 22475
rect 9630 22535 10000 22545
rect 9630 22475 9634 22535
rect 9686 22475 9944 22535
rect 9996 22475 10000 22535
rect 9630 22400 10000 22475
rect 10030 22535 10400 22545
rect 10030 22475 10034 22535
rect 10086 22475 10344 22535
rect 10396 22475 10400 22535
rect 10030 22400 10400 22475
rect 10430 22535 10800 22545
rect 10430 22475 10434 22535
rect 10486 22475 10744 22535
rect 10796 22475 10800 22535
rect 10430 22400 10800 22475
rect 10830 22535 11200 22545
rect 10830 22475 10834 22535
rect 10886 22475 11144 22535
rect 11196 22475 11200 22535
rect 10830 22400 11200 22475
rect 11230 22535 11600 22545
rect 11230 22475 11234 22535
rect 11286 22475 11544 22535
rect 11596 22475 11600 22535
rect 11230 22400 11600 22475
rect 11630 22535 12000 22545
rect 11630 22475 11634 22535
rect 11686 22475 11944 22535
rect 11996 22475 12000 22535
rect 11630 22400 12000 22475
rect 12030 22535 12400 22545
rect 12030 22475 12034 22535
rect 12086 22475 12344 22535
rect 12396 22475 12400 22535
rect 12030 22400 12400 22475
rect 12430 22535 12800 22545
rect 12430 22475 12434 22535
rect 12486 22475 12744 22535
rect 12796 22475 12800 22535
rect 12430 22400 12800 22475
rect 12830 22535 13200 22545
rect 12830 22475 12834 22535
rect 12886 22475 13144 22535
rect 13196 22475 13200 22535
rect 12830 22400 13200 22475
rect 30 22360 13200 22400
rect 30 22275 400 22360
rect 30 22215 34 22275
rect 86 22215 344 22275
rect 396 22215 400 22275
rect 30 22205 400 22215
rect 430 22275 800 22360
rect 430 22215 434 22275
rect 486 22215 744 22275
rect 796 22215 800 22275
rect 430 22205 800 22215
rect 830 22275 1200 22360
rect 830 22215 834 22275
rect 886 22215 1144 22275
rect 1196 22215 1200 22275
rect 830 22205 1200 22215
rect 1230 22275 1600 22360
rect 1230 22215 1234 22275
rect 1286 22215 1544 22275
rect 1596 22215 1600 22275
rect 1230 22205 1600 22215
rect 1630 22275 2000 22360
rect 1630 22215 1634 22275
rect 1686 22215 1944 22275
rect 1996 22215 2000 22275
rect 1630 22205 2000 22215
rect 2030 22275 2400 22360
rect 2030 22215 2034 22275
rect 2086 22215 2344 22275
rect 2396 22215 2400 22275
rect 2030 22205 2400 22215
rect 2430 22275 2800 22360
rect 2430 22215 2434 22275
rect 2486 22215 2744 22275
rect 2796 22215 2800 22275
rect 2430 22205 2800 22215
rect 2830 22275 3200 22360
rect 2830 22215 2834 22275
rect 2886 22215 3144 22275
rect 3196 22215 3200 22275
rect 2830 22205 3200 22215
rect 3230 22275 3600 22360
rect 3230 22215 3234 22275
rect 3286 22215 3544 22275
rect 3596 22215 3600 22275
rect 3230 22205 3600 22215
rect 3630 22275 4000 22360
rect 3630 22215 3634 22275
rect 3686 22215 3944 22275
rect 3996 22215 4000 22275
rect 3630 22205 4000 22215
rect 4030 22275 4400 22360
rect 4030 22215 4034 22275
rect 4086 22215 4344 22275
rect 4396 22215 4400 22275
rect 4030 22205 4400 22215
rect 4430 22275 4800 22360
rect 4430 22215 4434 22275
rect 4486 22215 4744 22275
rect 4796 22215 4800 22275
rect 4430 22205 4800 22215
rect 4830 22275 5200 22360
rect 4830 22215 4834 22275
rect 4886 22215 5144 22275
rect 5196 22215 5200 22275
rect 4830 22205 5200 22215
rect 5230 22275 5600 22360
rect 5230 22215 5234 22275
rect 5286 22215 5544 22275
rect 5596 22215 5600 22275
rect 5230 22205 5600 22215
rect 5630 22275 6000 22360
rect 5630 22215 5634 22275
rect 5686 22215 5944 22275
rect 5996 22215 6000 22275
rect 5630 22205 6000 22215
rect 6030 22275 6400 22360
rect 6030 22215 6034 22275
rect 6086 22215 6344 22275
rect 6396 22215 6400 22275
rect 6030 22205 6400 22215
rect 6430 22275 6800 22360
rect 6430 22215 6434 22275
rect 6486 22215 6744 22275
rect 6796 22215 6800 22275
rect 6430 22205 6800 22215
rect 6830 22275 7200 22360
rect 6830 22215 6834 22275
rect 6886 22215 7144 22275
rect 7196 22215 7200 22275
rect 6830 22205 7200 22215
rect 7230 22275 7600 22360
rect 7230 22215 7234 22275
rect 7286 22215 7544 22275
rect 7596 22215 7600 22275
rect 7230 22205 7600 22215
rect 7630 22275 8000 22360
rect 7630 22215 7634 22275
rect 7686 22215 7944 22275
rect 7996 22215 8000 22275
rect 7630 22205 8000 22215
rect 8030 22275 8400 22360
rect 8030 22215 8034 22275
rect 8086 22215 8344 22275
rect 8396 22215 8400 22275
rect 8030 22205 8400 22215
rect 8430 22275 8800 22360
rect 8430 22215 8434 22275
rect 8486 22215 8744 22275
rect 8796 22215 8800 22275
rect 8430 22205 8800 22215
rect 8830 22275 9200 22360
rect 8830 22215 8834 22275
rect 8886 22215 9144 22275
rect 9196 22215 9200 22275
rect 8830 22205 9200 22215
rect 9230 22275 9600 22360
rect 9230 22215 9234 22275
rect 9286 22215 9544 22275
rect 9596 22215 9600 22275
rect 9230 22205 9600 22215
rect 9630 22275 10000 22360
rect 9630 22215 9634 22275
rect 9686 22215 9944 22275
rect 9996 22215 10000 22275
rect 9630 22205 10000 22215
rect 10030 22275 10400 22360
rect 10030 22215 10034 22275
rect 10086 22215 10344 22275
rect 10396 22215 10400 22275
rect 10030 22205 10400 22215
rect 10430 22275 10800 22360
rect 10430 22215 10434 22275
rect 10486 22215 10744 22275
rect 10796 22215 10800 22275
rect 10430 22205 10800 22215
rect 10830 22275 11200 22360
rect 10830 22215 10834 22275
rect 10886 22215 11144 22275
rect 11196 22215 11200 22275
rect 10830 22205 11200 22215
rect 11230 22275 11600 22360
rect 11230 22215 11234 22275
rect 11286 22215 11544 22275
rect 11596 22215 11600 22275
rect 11230 22205 11600 22215
rect 11630 22275 12000 22360
rect 11630 22215 11634 22275
rect 11686 22215 11944 22275
rect 11996 22215 12000 22275
rect 11630 22205 12000 22215
rect 12030 22275 12400 22360
rect 12030 22215 12034 22275
rect 12086 22215 12344 22275
rect 12396 22215 12400 22275
rect 12030 22205 12400 22215
rect 12430 22275 12800 22360
rect 12430 22215 12434 22275
rect 12486 22215 12744 22275
rect 12796 22215 12800 22275
rect 12430 22205 12800 22215
rect 12830 22275 13200 22360
rect 12830 22215 12834 22275
rect 12886 22215 13144 22275
rect 13196 22215 13200 22275
rect 12830 22205 13200 22215
rect -330 22175 -324 22205
rect 30 22175 70 22205
rect 430 22175 470 22205
rect 830 22175 870 22205
rect 1230 22175 1270 22205
rect 1630 22175 1670 22205
rect 2030 22175 2070 22205
rect 2430 22175 2470 22205
rect 2830 22175 2870 22205
rect 3230 22175 3270 22205
rect 3630 22175 3670 22205
rect 4030 22175 4070 22205
rect 4430 22175 4470 22205
rect 4830 22175 4870 22205
rect 5230 22175 5270 22205
rect 5630 22175 5670 22205
rect 6030 22175 6070 22205
rect 6430 22175 6470 22205
rect 6830 22175 6870 22205
rect 7230 22175 7270 22205
rect 7630 22175 7670 22205
rect 8030 22175 8070 22205
rect 8430 22175 8470 22205
rect 8830 22175 8870 22205
rect 9230 22175 9270 22205
rect 9630 22175 9670 22205
rect 10030 22175 10070 22205
rect 10430 22175 10470 22205
rect 10830 22175 10870 22205
rect 11230 22175 11270 22205
rect 11630 22175 11670 22205
rect 12030 22175 12070 22205
rect 12430 22175 12470 22205
rect -330 22165 0 22175
rect -314 22105 -56 22165
rect -4 22105 0 22165
rect -330 21905 0 22105
rect -314 21845 -56 21905
rect -4 21845 0 21905
rect -330 21835 0 21845
rect 30 22165 400 22175
rect 30 22105 34 22165
rect 86 22105 344 22165
rect 396 22105 400 22165
rect 30 22030 400 22105
rect 430 22165 800 22175
rect 430 22105 434 22165
rect 486 22105 744 22165
rect 796 22105 800 22165
rect 430 22030 800 22105
rect 830 22165 1200 22175
rect 830 22105 834 22165
rect 886 22105 1144 22165
rect 1196 22105 1200 22165
rect 830 22030 1200 22105
rect 1230 22165 1600 22175
rect 1230 22105 1234 22165
rect 1286 22105 1544 22165
rect 1596 22105 1600 22165
rect 1230 22030 1600 22105
rect 1630 22165 2000 22175
rect 1630 22105 1634 22165
rect 1686 22105 1944 22165
rect 1996 22105 2000 22165
rect 1630 22030 2000 22105
rect 2030 22165 2400 22175
rect 2030 22105 2034 22165
rect 2086 22105 2344 22165
rect 2396 22105 2400 22165
rect 2030 22030 2400 22105
rect 2430 22165 2800 22175
rect 2430 22105 2434 22165
rect 2486 22105 2744 22165
rect 2796 22105 2800 22165
rect 2430 22030 2800 22105
rect 2830 22165 3200 22175
rect 2830 22105 2834 22165
rect 2886 22105 3144 22165
rect 3196 22105 3200 22165
rect 2830 22030 3200 22105
rect 3230 22165 3600 22175
rect 3230 22105 3234 22165
rect 3286 22105 3544 22165
rect 3596 22105 3600 22165
rect 3230 22030 3600 22105
rect 3630 22165 4000 22175
rect 3630 22105 3634 22165
rect 3686 22105 3944 22165
rect 3996 22105 4000 22165
rect 3630 22030 4000 22105
rect 4030 22165 4400 22175
rect 4030 22105 4034 22165
rect 4086 22105 4344 22165
rect 4396 22105 4400 22165
rect 4030 22030 4400 22105
rect 4430 22165 4800 22175
rect 4430 22105 4434 22165
rect 4486 22105 4744 22165
rect 4796 22105 4800 22165
rect 4430 22030 4800 22105
rect 4830 22165 5200 22175
rect 4830 22105 4834 22165
rect 4886 22105 5144 22165
rect 5196 22105 5200 22165
rect 4830 22030 5200 22105
rect 5230 22165 5600 22175
rect 5230 22105 5234 22165
rect 5286 22105 5544 22165
rect 5596 22105 5600 22165
rect 5230 22030 5600 22105
rect 5630 22165 6000 22175
rect 5630 22105 5634 22165
rect 5686 22105 5944 22165
rect 5996 22105 6000 22165
rect 5630 22030 6000 22105
rect 6030 22165 6400 22175
rect 6030 22105 6034 22165
rect 6086 22105 6344 22165
rect 6396 22105 6400 22165
rect 6030 22030 6400 22105
rect 6430 22165 6800 22175
rect 6430 22105 6434 22165
rect 6486 22105 6744 22165
rect 6796 22105 6800 22165
rect 6430 22030 6800 22105
rect 6830 22165 7200 22175
rect 6830 22105 6834 22165
rect 6886 22105 7144 22165
rect 7196 22105 7200 22165
rect 6830 22030 7200 22105
rect 7230 22165 7600 22175
rect 7230 22105 7234 22165
rect 7286 22105 7544 22165
rect 7596 22105 7600 22165
rect 7230 22030 7600 22105
rect 7630 22165 8000 22175
rect 7630 22105 7634 22165
rect 7686 22105 7944 22165
rect 7996 22105 8000 22165
rect 7630 22030 8000 22105
rect 8030 22165 8400 22175
rect 8030 22105 8034 22165
rect 8086 22105 8344 22165
rect 8396 22105 8400 22165
rect 8030 22030 8400 22105
rect 8430 22165 8800 22175
rect 8430 22105 8434 22165
rect 8486 22105 8744 22165
rect 8796 22105 8800 22165
rect 8430 22030 8800 22105
rect 8830 22165 9200 22175
rect 8830 22105 8834 22165
rect 8886 22105 9144 22165
rect 9196 22105 9200 22165
rect 8830 22030 9200 22105
rect 9230 22165 9600 22175
rect 9230 22105 9234 22165
rect 9286 22105 9544 22165
rect 9596 22105 9600 22165
rect 9230 22030 9600 22105
rect 9630 22165 10000 22175
rect 9630 22105 9634 22165
rect 9686 22105 9944 22165
rect 9996 22105 10000 22165
rect 9630 22030 10000 22105
rect 10030 22165 10400 22175
rect 10030 22105 10034 22165
rect 10086 22105 10344 22165
rect 10396 22105 10400 22165
rect 10030 22030 10400 22105
rect 10430 22165 10800 22175
rect 10430 22105 10434 22165
rect 10486 22105 10744 22165
rect 10796 22105 10800 22165
rect 10430 22030 10800 22105
rect 10830 22165 11200 22175
rect 10830 22105 10834 22165
rect 10886 22105 11144 22165
rect 11196 22105 11200 22165
rect 10830 22030 11200 22105
rect 11230 22165 11600 22175
rect 11230 22105 11234 22165
rect 11286 22105 11544 22165
rect 11596 22105 11600 22165
rect 11230 22030 11600 22105
rect 11630 22165 12000 22175
rect 11630 22105 11634 22165
rect 11686 22105 11944 22165
rect 11996 22105 12000 22165
rect 11630 22030 12000 22105
rect 12030 22165 12400 22175
rect 12030 22105 12034 22165
rect 12086 22105 12344 22165
rect 12396 22105 12400 22165
rect 12030 22030 12400 22105
rect 12430 22165 12800 22175
rect 12430 22105 12434 22165
rect 12486 22105 12744 22165
rect 12796 22105 12800 22165
rect 12430 22030 12800 22105
rect 12830 22165 13200 22175
rect 12830 22105 12834 22165
rect 12886 22105 13144 22165
rect 13196 22105 13200 22165
rect 12830 22030 13200 22105
rect 30 21990 13200 22030
rect 30 21905 400 21990
rect 30 21845 34 21905
rect 86 21845 344 21905
rect 396 21845 400 21905
rect 30 21835 400 21845
rect 430 21905 800 21990
rect 430 21845 434 21905
rect 486 21845 744 21905
rect 796 21845 800 21905
rect 430 21835 800 21845
rect 830 21905 1200 21990
rect 830 21845 834 21905
rect 886 21845 1144 21905
rect 1196 21845 1200 21905
rect 830 21835 1200 21845
rect 1230 21905 1600 21990
rect 1230 21845 1234 21905
rect 1286 21845 1544 21905
rect 1596 21845 1600 21905
rect 1230 21835 1600 21845
rect 1630 21905 2000 21990
rect 1630 21845 1634 21905
rect 1686 21845 1944 21905
rect 1996 21845 2000 21905
rect 1630 21835 2000 21845
rect 2030 21905 2400 21990
rect 2030 21845 2034 21905
rect 2086 21845 2344 21905
rect 2396 21845 2400 21905
rect 2030 21835 2400 21845
rect 2430 21905 2800 21990
rect 2430 21845 2434 21905
rect 2486 21845 2744 21905
rect 2796 21845 2800 21905
rect 2430 21835 2800 21845
rect 2830 21905 3200 21990
rect 2830 21845 2834 21905
rect 2886 21845 3144 21905
rect 3196 21845 3200 21905
rect 2830 21835 3200 21845
rect 3230 21905 3600 21990
rect 3230 21845 3234 21905
rect 3286 21845 3544 21905
rect 3596 21845 3600 21905
rect 3230 21835 3600 21845
rect 3630 21905 4000 21990
rect 3630 21845 3634 21905
rect 3686 21845 3944 21905
rect 3996 21845 4000 21905
rect 3630 21835 4000 21845
rect 4030 21905 4400 21990
rect 4030 21845 4034 21905
rect 4086 21845 4344 21905
rect 4396 21845 4400 21905
rect 4030 21835 4400 21845
rect 4430 21905 4800 21990
rect 4430 21845 4434 21905
rect 4486 21845 4744 21905
rect 4796 21845 4800 21905
rect 4430 21835 4800 21845
rect 4830 21905 5200 21990
rect 4830 21845 4834 21905
rect 4886 21845 5144 21905
rect 5196 21845 5200 21905
rect 4830 21835 5200 21845
rect 5230 21905 5600 21990
rect 5230 21845 5234 21905
rect 5286 21845 5544 21905
rect 5596 21845 5600 21905
rect 5230 21835 5600 21845
rect 5630 21905 6000 21990
rect 5630 21845 5634 21905
rect 5686 21845 5944 21905
rect 5996 21845 6000 21905
rect 5630 21835 6000 21845
rect 6030 21905 6400 21990
rect 6030 21845 6034 21905
rect 6086 21845 6344 21905
rect 6396 21845 6400 21905
rect 6030 21835 6400 21845
rect 6430 21905 6800 21990
rect 6430 21845 6434 21905
rect 6486 21845 6744 21905
rect 6796 21845 6800 21905
rect 6430 21835 6800 21845
rect 6830 21905 7200 21990
rect 6830 21845 6834 21905
rect 6886 21845 7144 21905
rect 7196 21845 7200 21905
rect 6830 21835 7200 21845
rect 7230 21905 7600 21990
rect 7230 21845 7234 21905
rect 7286 21845 7544 21905
rect 7596 21845 7600 21905
rect 7230 21835 7600 21845
rect 7630 21905 8000 21990
rect 7630 21845 7634 21905
rect 7686 21845 7944 21905
rect 7996 21845 8000 21905
rect 7630 21835 8000 21845
rect 8030 21905 8400 21990
rect 8030 21845 8034 21905
rect 8086 21845 8344 21905
rect 8396 21845 8400 21905
rect 8030 21835 8400 21845
rect 8430 21905 8800 21990
rect 8430 21845 8434 21905
rect 8486 21845 8744 21905
rect 8796 21845 8800 21905
rect 8430 21835 8800 21845
rect 8830 21905 9200 21990
rect 8830 21845 8834 21905
rect 8886 21845 9144 21905
rect 9196 21845 9200 21905
rect 8830 21835 9200 21845
rect 9230 21905 9600 21990
rect 9230 21845 9234 21905
rect 9286 21845 9544 21905
rect 9596 21845 9600 21905
rect 9230 21835 9600 21845
rect 9630 21905 10000 21990
rect 9630 21845 9634 21905
rect 9686 21845 9944 21905
rect 9996 21845 10000 21905
rect 9630 21835 10000 21845
rect 10030 21905 10400 21990
rect 10030 21845 10034 21905
rect 10086 21845 10344 21905
rect 10396 21845 10400 21905
rect 10030 21835 10400 21845
rect 10430 21905 10800 21990
rect 10430 21845 10434 21905
rect 10486 21845 10744 21905
rect 10796 21845 10800 21905
rect 10430 21835 10800 21845
rect 10830 21905 11200 21990
rect 10830 21845 10834 21905
rect 10886 21845 11144 21905
rect 11196 21845 11200 21905
rect 10830 21835 11200 21845
rect 11230 21905 11600 21990
rect 11230 21845 11234 21905
rect 11286 21845 11544 21905
rect 11596 21845 11600 21905
rect 11230 21835 11600 21845
rect 11630 21905 12000 21990
rect 11630 21845 11634 21905
rect 11686 21845 11944 21905
rect 11996 21845 12000 21905
rect 11630 21835 12000 21845
rect 12030 21905 12400 21990
rect 12030 21845 12034 21905
rect 12086 21845 12344 21905
rect 12396 21845 12400 21905
rect 12030 21835 12400 21845
rect 12430 21905 12800 21990
rect 12430 21845 12434 21905
rect 12486 21845 12744 21905
rect 12796 21845 12800 21905
rect 12430 21835 12800 21845
rect 12830 21905 13200 21990
rect 12830 21845 12834 21905
rect 12886 21845 13144 21905
rect 13196 21845 13200 21905
rect 12830 21835 13200 21845
rect -330 21805 -324 21835
rect 30 21805 70 21835
rect 430 21805 470 21835
rect 830 21805 870 21835
rect 1230 21805 1270 21835
rect 1630 21805 1670 21835
rect 2030 21805 2070 21835
rect 2430 21805 2470 21835
rect 2830 21805 2870 21835
rect 3230 21805 3270 21835
rect 3630 21805 3670 21835
rect 4030 21805 4070 21835
rect 4430 21805 4470 21835
rect 4830 21805 4870 21835
rect 5230 21805 5270 21835
rect 5630 21805 5670 21835
rect 6030 21805 6070 21835
rect 6430 21805 6470 21835
rect 6830 21805 6870 21835
rect 7230 21805 7270 21835
rect 7630 21805 7670 21835
rect 8030 21805 8070 21835
rect 8430 21805 8470 21835
rect 8830 21805 8870 21835
rect 9230 21805 9270 21835
rect 9630 21805 9670 21835
rect 10030 21805 10070 21835
rect 10430 21805 10470 21835
rect 10830 21805 10870 21835
rect 11230 21805 11270 21835
rect 11630 21805 11670 21835
rect 12030 21805 12070 21835
rect 12430 21805 12470 21835
rect -330 21795 0 21805
rect -314 21735 -56 21795
rect -4 21735 0 21795
rect -330 21535 0 21735
rect -314 21475 -56 21535
rect -4 21475 0 21535
rect -330 21465 0 21475
rect 30 21795 400 21805
rect 30 21735 34 21795
rect 86 21735 344 21795
rect 396 21735 400 21795
rect 30 21660 400 21735
rect 430 21795 800 21805
rect 430 21735 434 21795
rect 486 21735 744 21795
rect 796 21735 800 21795
rect 430 21660 800 21735
rect 830 21795 1200 21805
rect 830 21735 834 21795
rect 886 21735 1144 21795
rect 1196 21735 1200 21795
rect 830 21660 1200 21735
rect 1230 21795 1600 21805
rect 1230 21735 1234 21795
rect 1286 21735 1544 21795
rect 1596 21735 1600 21795
rect 1230 21660 1600 21735
rect 1630 21795 2000 21805
rect 1630 21735 1634 21795
rect 1686 21735 1944 21795
rect 1996 21735 2000 21795
rect 1630 21660 2000 21735
rect 2030 21795 2400 21805
rect 2030 21735 2034 21795
rect 2086 21735 2344 21795
rect 2396 21735 2400 21795
rect 2030 21660 2400 21735
rect 2430 21795 2800 21805
rect 2430 21735 2434 21795
rect 2486 21735 2744 21795
rect 2796 21735 2800 21795
rect 2430 21660 2800 21735
rect 2830 21795 3200 21805
rect 2830 21735 2834 21795
rect 2886 21735 3144 21795
rect 3196 21735 3200 21795
rect 2830 21660 3200 21735
rect 3230 21795 3600 21805
rect 3230 21735 3234 21795
rect 3286 21735 3544 21795
rect 3596 21735 3600 21795
rect 3230 21660 3600 21735
rect 3630 21795 4000 21805
rect 3630 21735 3634 21795
rect 3686 21735 3944 21795
rect 3996 21735 4000 21795
rect 3630 21660 4000 21735
rect 4030 21795 4400 21805
rect 4030 21735 4034 21795
rect 4086 21735 4344 21795
rect 4396 21735 4400 21795
rect 4030 21660 4400 21735
rect 4430 21795 4800 21805
rect 4430 21735 4434 21795
rect 4486 21735 4744 21795
rect 4796 21735 4800 21795
rect 4430 21660 4800 21735
rect 4830 21795 5200 21805
rect 4830 21735 4834 21795
rect 4886 21735 5144 21795
rect 5196 21735 5200 21795
rect 4830 21660 5200 21735
rect 5230 21795 5600 21805
rect 5230 21735 5234 21795
rect 5286 21735 5544 21795
rect 5596 21735 5600 21795
rect 5230 21660 5600 21735
rect 5630 21795 6000 21805
rect 5630 21735 5634 21795
rect 5686 21735 5944 21795
rect 5996 21735 6000 21795
rect 5630 21660 6000 21735
rect 6030 21795 6400 21805
rect 6030 21735 6034 21795
rect 6086 21735 6344 21795
rect 6396 21735 6400 21795
rect 6030 21660 6400 21735
rect 6430 21795 6800 21805
rect 6430 21735 6434 21795
rect 6486 21735 6744 21795
rect 6796 21735 6800 21795
rect 6430 21660 6800 21735
rect 6830 21795 7200 21805
rect 6830 21735 6834 21795
rect 6886 21735 7144 21795
rect 7196 21735 7200 21795
rect 6830 21660 7200 21735
rect 7230 21795 7600 21805
rect 7230 21735 7234 21795
rect 7286 21735 7544 21795
rect 7596 21735 7600 21795
rect 7230 21660 7600 21735
rect 7630 21795 8000 21805
rect 7630 21735 7634 21795
rect 7686 21735 7944 21795
rect 7996 21735 8000 21795
rect 7630 21660 8000 21735
rect 8030 21795 8400 21805
rect 8030 21735 8034 21795
rect 8086 21735 8344 21795
rect 8396 21735 8400 21795
rect 8030 21660 8400 21735
rect 8430 21795 8800 21805
rect 8430 21735 8434 21795
rect 8486 21735 8744 21795
rect 8796 21735 8800 21795
rect 8430 21660 8800 21735
rect 8830 21795 9200 21805
rect 8830 21735 8834 21795
rect 8886 21735 9144 21795
rect 9196 21735 9200 21795
rect 8830 21660 9200 21735
rect 9230 21795 9600 21805
rect 9230 21735 9234 21795
rect 9286 21735 9544 21795
rect 9596 21735 9600 21795
rect 9230 21660 9600 21735
rect 9630 21795 10000 21805
rect 9630 21735 9634 21795
rect 9686 21735 9944 21795
rect 9996 21735 10000 21795
rect 9630 21660 10000 21735
rect 10030 21795 10400 21805
rect 10030 21735 10034 21795
rect 10086 21735 10344 21795
rect 10396 21735 10400 21795
rect 10030 21660 10400 21735
rect 10430 21795 10800 21805
rect 10430 21735 10434 21795
rect 10486 21735 10744 21795
rect 10796 21735 10800 21795
rect 10430 21660 10800 21735
rect 10830 21795 11200 21805
rect 10830 21735 10834 21795
rect 10886 21735 11144 21795
rect 11196 21735 11200 21795
rect 10830 21660 11200 21735
rect 11230 21795 11600 21805
rect 11230 21735 11234 21795
rect 11286 21735 11544 21795
rect 11596 21735 11600 21795
rect 11230 21660 11600 21735
rect 11630 21795 12000 21805
rect 11630 21735 11634 21795
rect 11686 21735 11944 21795
rect 11996 21735 12000 21795
rect 11630 21660 12000 21735
rect 12030 21795 12400 21805
rect 12030 21735 12034 21795
rect 12086 21735 12344 21795
rect 12396 21735 12400 21795
rect 12030 21660 12400 21735
rect 12430 21795 12800 21805
rect 12430 21735 12434 21795
rect 12486 21735 12744 21795
rect 12796 21735 12800 21795
rect 12430 21660 12800 21735
rect 12830 21795 13200 21805
rect 12830 21735 12834 21795
rect 12886 21735 13144 21795
rect 13196 21735 13200 21795
rect 12830 21660 13200 21735
rect 30 21620 13200 21660
rect 30 21535 400 21620
rect 30 21475 34 21535
rect 86 21475 344 21535
rect 396 21475 400 21535
rect 30 21465 400 21475
rect 430 21535 800 21620
rect 430 21475 434 21535
rect 486 21475 744 21535
rect 796 21475 800 21535
rect 430 21465 800 21475
rect 830 21535 1200 21620
rect 830 21475 834 21535
rect 886 21475 1144 21535
rect 1196 21475 1200 21535
rect 830 21465 1200 21475
rect 1230 21535 1600 21620
rect 1230 21475 1234 21535
rect 1286 21475 1544 21535
rect 1596 21475 1600 21535
rect 1230 21465 1600 21475
rect 1630 21535 2000 21620
rect 1630 21475 1634 21535
rect 1686 21475 1944 21535
rect 1996 21475 2000 21535
rect 1630 21465 2000 21475
rect 2030 21535 2400 21620
rect 2030 21475 2034 21535
rect 2086 21475 2344 21535
rect 2396 21475 2400 21535
rect 2030 21465 2400 21475
rect 2430 21535 2800 21620
rect 2430 21475 2434 21535
rect 2486 21475 2744 21535
rect 2796 21475 2800 21535
rect 2430 21465 2800 21475
rect 2830 21535 3200 21620
rect 2830 21475 2834 21535
rect 2886 21475 3144 21535
rect 3196 21475 3200 21535
rect 2830 21465 3200 21475
rect 3230 21535 3600 21620
rect 3230 21475 3234 21535
rect 3286 21475 3544 21535
rect 3596 21475 3600 21535
rect 3230 21465 3600 21475
rect 3630 21535 4000 21620
rect 3630 21475 3634 21535
rect 3686 21475 3944 21535
rect 3996 21475 4000 21535
rect 3630 21465 4000 21475
rect 4030 21535 4400 21620
rect 4030 21475 4034 21535
rect 4086 21475 4344 21535
rect 4396 21475 4400 21535
rect 4030 21465 4400 21475
rect 4430 21535 4800 21620
rect 4430 21475 4434 21535
rect 4486 21475 4744 21535
rect 4796 21475 4800 21535
rect 4430 21465 4800 21475
rect 4830 21535 5200 21620
rect 4830 21475 4834 21535
rect 4886 21475 5144 21535
rect 5196 21475 5200 21535
rect 4830 21465 5200 21475
rect 5230 21535 5600 21620
rect 5230 21475 5234 21535
rect 5286 21475 5544 21535
rect 5596 21475 5600 21535
rect 5230 21465 5600 21475
rect 5630 21535 6000 21620
rect 5630 21475 5634 21535
rect 5686 21475 5944 21535
rect 5996 21475 6000 21535
rect 5630 21465 6000 21475
rect 6030 21535 6400 21620
rect 6030 21475 6034 21535
rect 6086 21475 6344 21535
rect 6396 21475 6400 21535
rect 6030 21465 6400 21475
rect 6430 21535 6800 21620
rect 6430 21475 6434 21535
rect 6486 21475 6744 21535
rect 6796 21475 6800 21535
rect 6430 21465 6800 21475
rect 6830 21535 7200 21620
rect 6830 21475 6834 21535
rect 6886 21475 7144 21535
rect 7196 21475 7200 21535
rect 6830 21465 7200 21475
rect 7230 21535 7600 21620
rect 7230 21475 7234 21535
rect 7286 21475 7544 21535
rect 7596 21475 7600 21535
rect 7230 21465 7600 21475
rect 7630 21535 8000 21620
rect 7630 21475 7634 21535
rect 7686 21475 7944 21535
rect 7996 21475 8000 21535
rect 7630 21465 8000 21475
rect 8030 21535 8400 21620
rect 8030 21475 8034 21535
rect 8086 21475 8344 21535
rect 8396 21475 8400 21535
rect 8030 21465 8400 21475
rect 8430 21535 8800 21620
rect 8430 21475 8434 21535
rect 8486 21475 8744 21535
rect 8796 21475 8800 21535
rect 8430 21465 8800 21475
rect 8830 21535 9200 21620
rect 8830 21475 8834 21535
rect 8886 21475 9144 21535
rect 9196 21475 9200 21535
rect 8830 21465 9200 21475
rect 9230 21535 9600 21620
rect 9230 21475 9234 21535
rect 9286 21475 9544 21535
rect 9596 21475 9600 21535
rect 9230 21465 9600 21475
rect 9630 21535 10000 21620
rect 9630 21475 9634 21535
rect 9686 21475 9944 21535
rect 9996 21475 10000 21535
rect 9630 21465 10000 21475
rect 10030 21535 10400 21620
rect 10030 21475 10034 21535
rect 10086 21475 10344 21535
rect 10396 21475 10400 21535
rect 10030 21465 10400 21475
rect 10430 21535 10800 21620
rect 10430 21475 10434 21535
rect 10486 21475 10744 21535
rect 10796 21475 10800 21535
rect 10430 21465 10800 21475
rect 10830 21535 11200 21620
rect 10830 21475 10834 21535
rect 10886 21475 11144 21535
rect 11196 21475 11200 21535
rect 10830 21465 11200 21475
rect 11230 21535 11600 21620
rect 11230 21475 11234 21535
rect 11286 21475 11544 21535
rect 11596 21475 11600 21535
rect 11230 21465 11600 21475
rect 11630 21535 12000 21620
rect 11630 21475 11634 21535
rect 11686 21475 11944 21535
rect 11996 21475 12000 21535
rect 11630 21465 12000 21475
rect 12030 21535 12400 21620
rect 12030 21475 12034 21535
rect 12086 21475 12344 21535
rect 12396 21475 12400 21535
rect 12030 21465 12400 21475
rect 12430 21535 12800 21620
rect 12430 21475 12434 21535
rect 12486 21475 12744 21535
rect 12796 21475 12800 21535
rect 12430 21465 12800 21475
rect 12830 21535 13200 21620
rect 12830 21475 12834 21535
rect 12886 21475 13144 21535
rect 13196 21475 13200 21535
rect 12830 21465 13200 21475
rect -330 21435 -324 21465
rect 30 21435 70 21465
rect 430 21435 470 21465
rect 830 21435 870 21465
rect 1230 21435 1270 21465
rect 1630 21435 1670 21465
rect 2030 21435 2070 21465
rect 2430 21435 2470 21465
rect 2830 21435 2870 21465
rect 3230 21435 3270 21465
rect 3630 21435 3670 21465
rect 4030 21435 4070 21465
rect 4430 21435 4470 21465
rect 4830 21435 4870 21465
rect 5230 21435 5270 21465
rect 5630 21435 5670 21465
rect 6030 21435 6070 21465
rect 6430 21435 6470 21465
rect 6830 21435 6870 21465
rect 7230 21435 7270 21465
rect 7630 21435 7670 21465
rect 8030 21435 8070 21465
rect 8430 21435 8470 21465
rect 8830 21435 8870 21465
rect 9230 21435 9270 21465
rect 9630 21435 9670 21465
rect 10030 21435 10070 21465
rect 10430 21435 10470 21465
rect 10830 21435 10870 21465
rect 11230 21435 11270 21465
rect 11630 21435 11670 21465
rect 12030 21435 12070 21465
rect 12430 21435 12470 21465
rect -330 21425 0 21435
rect -314 21365 -56 21425
rect -4 21365 0 21425
rect -330 21165 0 21365
rect -314 21105 -56 21165
rect -4 21105 0 21165
rect -330 21095 0 21105
rect 30 21425 400 21435
rect 30 21365 34 21425
rect 86 21365 344 21425
rect 396 21365 400 21425
rect 30 21290 400 21365
rect 430 21425 800 21435
rect 430 21365 434 21425
rect 486 21365 744 21425
rect 796 21365 800 21425
rect 430 21290 800 21365
rect 830 21425 1200 21435
rect 830 21365 834 21425
rect 886 21365 1144 21425
rect 1196 21365 1200 21425
rect 830 21290 1200 21365
rect 1230 21425 1600 21435
rect 1230 21365 1234 21425
rect 1286 21365 1544 21425
rect 1596 21365 1600 21425
rect 1230 21290 1600 21365
rect 1630 21425 2000 21435
rect 1630 21365 1634 21425
rect 1686 21365 1944 21425
rect 1996 21365 2000 21425
rect 1630 21290 2000 21365
rect 2030 21425 2400 21435
rect 2030 21365 2034 21425
rect 2086 21365 2344 21425
rect 2396 21365 2400 21425
rect 2030 21290 2400 21365
rect 2430 21425 2800 21435
rect 2430 21365 2434 21425
rect 2486 21365 2744 21425
rect 2796 21365 2800 21425
rect 2430 21290 2800 21365
rect 2830 21425 3200 21435
rect 2830 21365 2834 21425
rect 2886 21365 3144 21425
rect 3196 21365 3200 21425
rect 2830 21290 3200 21365
rect 3230 21425 3600 21435
rect 3230 21365 3234 21425
rect 3286 21365 3544 21425
rect 3596 21365 3600 21425
rect 3230 21290 3600 21365
rect 3630 21425 4000 21435
rect 3630 21365 3634 21425
rect 3686 21365 3944 21425
rect 3996 21365 4000 21425
rect 3630 21290 4000 21365
rect 4030 21425 4400 21435
rect 4030 21365 4034 21425
rect 4086 21365 4344 21425
rect 4396 21365 4400 21425
rect 4030 21290 4400 21365
rect 4430 21425 4800 21435
rect 4430 21365 4434 21425
rect 4486 21365 4744 21425
rect 4796 21365 4800 21425
rect 4430 21290 4800 21365
rect 4830 21425 5200 21435
rect 4830 21365 4834 21425
rect 4886 21365 5144 21425
rect 5196 21365 5200 21425
rect 4830 21290 5200 21365
rect 5230 21425 5600 21435
rect 5230 21365 5234 21425
rect 5286 21365 5544 21425
rect 5596 21365 5600 21425
rect 5230 21290 5600 21365
rect 5630 21425 6000 21435
rect 5630 21365 5634 21425
rect 5686 21365 5944 21425
rect 5996 21365 6000 21425
rect 5630 21290 6000 21365
rect 6030 21425 6400 21435
rect 6030 21365 6034 21425
rect 6086 21365 6344 21425
rect 6396 21365 6400 21425
rect 6030 21290 6400 21365
rect 6430 21425 6800 21435
rect 6430 21365 6434 21425
rect 6486 21365 6744 21425
rect 6796 21365 6800 21425
rect 6430 21290 6800 21365
rect 6830 21425 7200 21435
rect 6830 21365 6834 21425
rect 6886 21365 7144 21425
rect 7196 21365 7200 21425
rect 6830 21290 7200 21365
rect 7230 21425 7600 21435
rect 7230 21365 7234 21425
rect 7286 21365 7544 21425
rect 7596 21365 7600 21425
rect 7230 21290 7600 21365
rect 7630 21425 8000 21435
rect 7630 21365 7634 21425
rect 7686 21365 7944 21425
rect 7996 21365 8000 21425
rect 7630 21290 8000 21365
rect 8030 21425 8400 21435
rect 8030 21365 8034 21425
rect 8086 21365 8344 21425
rect 8396 21365 8400 21425
rect 8030 21290 8400 21365
rect 8430 21425 8800 21435
rect 8430 21365 8434 21425
rect 8486 21365 8744 21425
rect 8796 21365 8800 21425
rect 8430 21290 8800 21365
rect 8830 21425 9200 21435
rect 8830 21365 8834 21425
rect 8886 21365 9144 21425
rect 9196 21365 9200 21425
rect 8830 21290 9200 21365
rect 9230 21425 9600 21435
rect 9230 21365 9234 21425
rect 9286 21365 9544 21425
rect 9596 21365 9600 21425
rect 9230 21290 9600 21365
rect 9630 21425 10000 21435
rect 9630 21365 9634 21425
rect 9686 21365 9944 21425
rect 9996 21365 10000 21425
rect 9630 21290 10000 21365
rect 10030 21425 10400 21435
rect 10030 21365 10034 21425
rect 10086 21365 10344 21425
rect 10396 21365 10400 21425
rect 10030 21290 10400 21365
rect 10430 21425 10800 21435
rect 10430 21365 10434 21425
rect 10486 21365 10744 21425
rect 10796 21365 10800 21425
rect 10430 21290 10800 21365
rect 10830 21425 11200 21435
rect 10830 21365 10834 21425
rect 10886 21365 11144 21425
rect 11196 21365 11200 21425
rect 10830 21290 11200 21365
rect 11230 21425 11600 21435
rect 11230 21365 11234 21425
rect 11286 21365 11544 21425
rect 11596 21365 11600 21425
rect 11230 21290 11600 21365
rect 11630 21425 12000 21435
rect 11630 21365 11634 21425
rect 11686 21365 11944 21425
rect 11996 21365 12000 21425
rect 11630 21290 12000 21365
rect 12030 21425 12400 21435
rect 12030 21365 12034 21425
rect 12086 21365 12344 21425
rect 12396 21365 12400 21425
rect 12030 21290 12400 21365
rect 12430 21425 12800 21435
rect 12430 21365 12434 21425
rect 12486 21365 12744 21425
rect 12796 21365 12800 21425
rect 12430 21290 12800 21365
rect 12830 21425 13200 21435
rect 12830 21365 12834 21425
rect 12886 21365 13144 21425
rect 13196 21365 13200 21425
rect 12830 21290 13200 21365
rect 30 21250 13200 21290
rect 30 21165 400 21250
rect 30 21105 34 21165
rect 86 21105 344 21165
rect 396 21105 400 21165
rect 30 21095 400 21105
rect 430 21165 800 21250
rect 430 21105 434 21165
rect 486 21105 744 21165
rect 796 21105 800 21165
rect 430 21095 800 21105
rect 830 21165 1200 21250
rect 830 21105 834 21165
rect 886 21105 1144 21165
rect 1196 21105 1200 21165
rect 830 21095 1200 21105
rect 1230 21165 1600 21250
rect 1230 21105 1234 21165
rect 1286 21105 1544 21165
rect 1596 21105 1600 21165
rect 1230 21095 1600 21105
rect 1630 21165 2000 21250
rect 1630 21105 1634 21165
rect 1686 21105 1944 21165
rect 1996 21105 2000 21165
rect 1630 21095 2000 21105
rect 2030 21165 2400 21250
rect 2030 21105 2034 21165
rect 2086 21105 2344 21165
rect 2396 21105 2400 21165
rect 2030 21095 2400 21105
rect 2430 21165 2800 21250
rect 2430 21105 2434 21165
rect 2486 21105 2744 21165
rect 2796 21105 2800 21165
rect 2430 21095 2800 21105
rect 2830 21165 3200 21250
rect 2830 21105 2834 21165
rect 2886 21105 3144 21165
rect 3196 21105 3200 21165
rect 2830 21095 3200 21105
rect 3230 21165 3600 21250
rect 3230 21105 3234 21165
rect 3286 21105 3544 21165
rect 3596 21105 3600 21165
rect 3230 21095 3600 21105
rect 3630 21165 4000 21250
rect 3630 21105 3634 21165
rect 3686 21105 3944 21165
rect 3996 21105 4000 21165
rect 3630 21095 4000 21105
rect 4030 21165 4400 21250
rect 4030 21105 4034 21165
rect 4086 21105 4344 21165
rect 4396 21105 4400 21165
rect 4030 21095 4400 21105
rect 4430 21165 4800 21250
rect 4430 21105 4434 21165
rect 4486 21105 4744 21165
rect 4796 21105 4800 21165
rect 4430 21095 4800 21105
rect 4830 21165 5200 21250
rect 4830 21105 4834 21165
rect 4886 21105 5144 21165
rect 5196 21105 5200 21165
rect 4830 21095 5200 21105
rect 5230 21165 5600 21250
rect 5230 21105 5234 21165
rect 5286 21105 5544 21165
rect 5596 21105 5600 21165
rect 5230 21095 5600 21105
rect 5630 21165 6000 21250
rect 5630 21105 5634 21165
rect 5686 21105 5944 21165
rect 5996 21105 6000 21165
rect 5630 21095 6000 21105
rect 6030 21165 6400 21250
rect 6030 21105 6034 21165
rect 6086 21105 6344 21165
rect 6396 21105 6400 21165
rect 6030 21095 6400 21105
rect 6430 21165 6800 21250
rect 6430 21105 6434 21165
rect 6486 21105 6744 21165
rect 6796 21105 6800 21165
rect 6430 21095 6800 21105
rect 6830 21165 7200 21250
rect 6830 21105 6834 21165
rect 6886 21105 7144 21165
rect 7196 21105 7200 21165
rect 6830 21095 7200 21105
rect 7230 21165 7600 21250
rect 7230 21105 7234 21165
rect 7286 21105 7544 21165
rect 7596 21105 7600 21165
rect 7230 21095 7600 21105
rect 7630 21165 8000 21250
rect 7630 21105 7634 21165
rect 7686 21105 7944 21165
rect 7996 21105 8000 21165
rect 7630 21095 8000 21105
rect 8030 21165 8400 21250
rect 8030 21105 8034 21165
rect 8086 21105 8344 21165
rect 8396 21105 8400 21165
rect 8030 21095 8400 21105
rect 8430 21165 8800 21250
rect 8430 21105 8434 21165
rect 8486 21105 8744 21165
rect 8796 21105 8800 21165
rect 8430 21095 8800 21105
rect 8830 21165 9200 21250
rect 8830 21105 8834 21165
rect 8886 21105 9144 21165
rect 9196 21105 9200 21165
rect 8830 21095 9200 21105
rect 9230 21165 9600 21250
rect 9230 21105 9234 21165
rect 9286 21105 9544 21165
rect 9596 21105 9600 21165
rect 9230 21095 9600 21105
rect 9630 21165 10000 21250
rect 9630 21105 9634 21165
rect 9686 21105 9944 21165
rect 9996 21105 10000 21165
rect 9630 21095 10000 21105
rect 10030 21165 10400 21250
rect 10030 21105 10034 21165
rect 10086 21105 10344 21165
rect 10396 21105 10400 21165
rect 10030 21095 10400 21105
rect 10430 21165 10800 21250
rect 10430 21105 10434 21165
rect 10486 21105 10744 21165
rect 10796 21105 10800 21165
rect 10430 21095 10800 21105
rect 10830 21165 11200 21250
rect 10830 21105 10834 21165
rect 10886 21105 11144 21165
rect 11196 21105 11200 21165
rect 10830 21095 11200 21105
rect 11230 21165 11600 21250
rect 11230 21105 11234 21165
rect 11286 21105 11544 21165
rect 11596 21105 11600 21165
rect 11230 21095 11600 21105
rect 11630 21165 12000 21250
rect 11630 21105 11634 21165
rect 11686 21105 11944 21165
rect 11996 21105 12000 21165
rect 11630 21095 12000 21105
rect 12030 21165 12400 21250
rect 12030 21105 12034 21165
rect 12086 21105 12344 21165
rect 12396 21105 12400 21165
rect 12030 21095 12400 21105
rect 12430 21165 12800 21250
rect 12430 21105 12434 21165
rect 12486 21105 12744 21165
rect 12796 21105 12800 21165
rect 12430 21095 12800 21105
rect 12830 21165 13200 21250
rect 12830 21105 12834 21165
rect 12886 21105 13144 21165
rect 13196 21105 13200 21165
rect 12830 21095 13200 21105
rect -330 21065 -324 21095
rect 30 21065 70 21095
rect 430 21065 470 21095
rect 830 21065 870 21095
rect 1230 21065 1270 21095
rect 1630 21065 1670 21095
rect 2030 21065 2070 21095
rect 2430 21065 2470 21095
rect 2830 21065 2870 21095
rect 3230 21065 3270 21095
rect 3630 21065 3670 21095
rect 4030 21065 4070 21095
rect 4430 21065 4470 21095
rect 4830 21065 4870 21095
rect 5230 21065 5270 21095
rect 5630 21065 5670 21095
rect 6030 21065 6070 21095
rect 6430 21065 6470 21095
rect 6830 21065 6870 21095
rect 7230 21065 7270 21095
rect 7630 21065 7670 21095
rect 8030 21065 8070 21095
rect 8430 21065 8470 21095
rect 8830 21065 8870 21095
rect 9230 21065 9270 21095
rect 9630 21065 9670 21095
rect 10030 21065 10070 21095
rect 10430 21065 10470 21095
rect 10830 21065 10870 21095
rect 11230 21065 11270 21095
rect 11630 21065 11670 21095
rect 12030 21065 12070 21095
rect 12430 21065 12470 21095
rect -330 21055 0 21065
rect -314 20995 -56 21055
rect -4 20995 0 21055
rect -330 20795 0 20995
rect -314 20735 -56 20795
rect -4 20735 0 20795
rect -330 20725 0 20735
rect 30 21055 400 21065
rect 30 20995 34 21055
rect 86 20995 344 21055
rect 396 20995 400 21055
rect 30 20920 400 20995
rect 430 21055 800 21065
rect 430 20995 434 21055
rect 486 20995 744 21055
rect 796 20995 800 21055
rect 430 20920 800 20995
rect 830 21055 1200 21065
rect 830 20995 834 21055
rect 886 20995 1144 21055
rect 1196 20995 1200 21055
rect 830 20920 1200 20995
rect 1230 21055 1600 21065
rect 1230 20995 1234 21055
rect 1286 20995 1544 21055
rect 1596 20995 1600 21055
rect 1230 20920 1600 20995
rect 1630 21055 2000 21065
rect 1630 20995 1634 21055
rect 1686 20995 1944 21055
rect 1996 20995 2000 21055
rect 1630 20920 2000 20995
rect 2030 21055 2400 21065
rect 2030 20995 2034 21055
rect 2086 20995 2344 21055
rect 2396 20995 2400 21055
rect 2030 20920 2400 20995
rect 2430 21055 2800 21065
rect 2430 20995 2434 21055
rect 2486 20995 2744 21055
rect 2796 20995 2800 21055
rect 2430 20920 2800 20995
rect 2830 21055 3200 21065
rect 2830 20995 2834 21055
rect 2886 20995 3144 21055
rect 3196 20995 3200 21055
rect 2830 20920 3200 20995
rect 3230 21055 3600 21065
rect 3230 20995 3234 21055
rect 3286 20995 3544 21055
rect 3596 20995 3600 21055
rect 3230 20920 3600 20995
rect 3630 21055 4000 21065
rect 3630 20995 3634 21055
rect 3686 20995 3944 21055
rect 3996 20995 4000 21055
rect 3630 20920 4000 20995
rect 4030 21055 4400 21065
rect 4030 20995 4034 21055
rect 4086 20995 4344 21055
rect 4396 20995 4400 21055
rect 4030 20920 4400 20995
rect 4430 21055 4800 21065
rect 4430 20995 4434 21055
rect 4486 20995 4744 21055
rect 4796 20995 4800 21055
rect 4430 20920 4800 20995
rect 4830 21055 5200 21065
rect 4830 20995 4834 21055
rect 4886 20995 5144 21055
rect 5196 20995 5200 21055
rect 4830 20920 5200 20995
rect 5230 21055 5600 21065
rect 5230 20995 5234 21055
rect 5286 20995 5544 21055
rect 5596 20995 5600 21055
rect 5230 20920 5600 20995
rect 5630 21055 6000 21065
rect 5630 20995 5634 21055
rect 5686 20995 5944 21055
rect 5996 20995 6000 21055
rect 5630 20920 6000 20995
rect 6030 21055 6400 21065
rect 6030 20995 6034 21055
rect 6086 20995 6344 21055
rect 6396 20995 6400 21055
rect 6030 20920 6400 20995
rect 6430 21055 6800 21065
rect 6430 20995 6434 21055
rect 6486 20995 6744 21055
rect 6796 20995 6800 21055
rect 6430 20920 6800 20995
rect 6830 21055 7200 21065
rect 6830 20995 6834 21055
rect 6886 20995 7144 21055
rect 7196 20995 7200 21055
rect 6830 20920 7200 20995
rect 7230 21055 7600 21065
rect 7230 20995 7234 21055
rect 7286 20995 7544 21055
rect 7596 20995 7600 21055
rect 7230 20920 7600 20995
rect 7630 21055 8000 21065
rect 7630 20995 7634 21055
rect 7686 20995 7944 21055
rect 7996 20995 8000 21055
rect 7630 20920 8000 20995
rect 8030 21055 8400 21065
rect 8030 20995 8034 21055
rect 8086 20995 8344 21055
rect 8396 20995 8400 21055
rect 8030 20920 8400 20995
rect 8430 21055 8800 21065
rect 8430 20995 8434 21055
rect 8486 20995 8744 21055
rect 8796 20995 8800 21055
rect 8430 20920 8800 20995
rect 8830 21055 9200 21065
rect 8830 20995 8834 21055
rect 8886 20995 9144 21055
rect 9196 20995 9200 21055
rect 8830 20920 9200 20995
rect 9230 21055 9600 21065
rect 9230 20995 9234 21055
rect 9286 20995 9544 21055
rect 9596 20995 9600 21055
rect 9230 20920 9600 20995
rect 9630 21055 10000 21065
rect 9630 20995 9634 21055
rect 9686 20995 9944 21055
rect 9996 20995 10000 21055
rect 9630 20920 10000 20995
rect 10030 21055 10400 21065
rect 10030 20995 10034 21055
rect 10086 20995 10344 21055
rect 10396 20995 10400 21055
rect 10030 20920 10400 20995
rect 10430 21055 10800 21065
rect 10430 20995 10434 21055
rect 10486 20995 10744 21055
rect 10796 20995 10800 21055
rect 10430 20920 10800 20995
rect 10830 21055 11200 21065
rect 10830 20995 10834 21055
rect 10886 20995 11144 21055
rect 11196 20995 11200 21055
rect 10830 20920 11200 20995
rect 11230 21055 11600 21065
rect 11230 20995 11234 21055
rect 11286 20995 11544 21055
rect 11596 20995 11600 21055
rect 11230 20920 11600 20995
rect 11630 21055 12000 21065
rect 11630 20995 11634 21055
rect 11686 20995 11944 21055
rect 11996 20995 12000 21055
rect 11630 20920 12000 20995
rect 12030 21055 12400 21065
rect 12030 20995 12034 21055
rect 12086 20995 12344 21055
rect 12396 20995 12400 21055
rect 12030 20920 12400 20995
rect 12430 21055 12800 21065
rect 12430 20995 12434 21055
rect 12486 20995 12744 21055
rect 12796 20995 12800 21055
rect 12430 20920 12800 20995
rect 12830 21055 13200 21065
rect 12830 20995 12834 21055
rect 12886 20995 13144 21055
rect 13196 20995 13200 21055
rect 12830 20920 13200 20995
rect 30 20880 13200 20920
rect 30 20795 400 20880
rect 30 20735 34 20795
rect 86 20735 344 20795
rect 396 20735 400 20795
rect 30 20725 400 20735
rect 430 20795 800 20880
rect 430 20735 434 20795
rect 486 20735 744 20795
rect 796 20735 800 20795
rect 430 20725 800 20735
rect 830 20795 1200 20880
rect 830 20735 834 20795
rect 886 20735 1144 20795
rect 1196 20735 1200 20795
rect 830 20725 1200 20735
rect 1230 20795 1600 20880
rect 1230 20735 1234 20795
rect 1286 20735 1544 20795
rect 1596 20735 1600 20795
rect 1230 20725 1600 20735
rect 1630 20795 2000 20880
rect 1630 20735 1634 20795
rect 1686 20735 1944 20795
rect 1996 20735 2000 20795
rect 1630 20725 2000 20735
rect 2030 20795 2400 20880
rect 2030 20735 2034 20795
rect 2086 20735 2344 20795
rect 2396 20735 2400 20795
rect 2030 20725 2400 20735
rect 2430 20795 2800 20880
rect 2430 20735 2434 20795
rect 2486 20735 2744 20795
rect 2796 20735 2800 20795
rect 2430 20725 2800 20735
rect 2830 20795 3200 20880
rect 2830 20735 2834 20795
rect 2886 20735 3144 20795
rect 3196 20735 3200 20795
rect 2830 20725 3200 20735
rect 3230 20795 3600 20880
rect 3230 20735 3234 20795
rect 3286 20735 3544 20795
rect 3596 20735 3600 20795
rect 3230 20725 3600 20735
rect 3630 20795 4000 20880
rect 3630 20735 3634 20795
rect 3686 20735 3944 20795
rect 3996 20735 4000 20795
rect 3630 20725 4000 20735
rect 4030 20795 4400 20880
rect 4030 20735 4034 20795
rect 4086 20735 4344 20795
rect 4396 20735 4400 20795
rect 4030 20725 4400 20735
rect 4430 20795 4800 20880
rect 4430 20735 4434 20795
rect 4486 20735 4744 20795
rect 4796 20735 4800 20795
rect 4430 20725 4800 20735
rect 4830 20795 5200 20880
rect 4830 20735 4834 20795
rect 4886 20735 5144 20795
rect 5196 20735 5200 20795
rect 4830 20725 5200 20735
rect 5230 20795 5600 20880
rect 5230 20735 5234 20795
rect 5286 20735 5544 20795
rect 5596 20735 5600 20795
rect 5230 20725 5600 20735
rect 5630 20795 6000 20880
rect 5630 20735 5634 20795
rect 5686 20735 5944 20795
rect 5996 20735 6000 20795
rect 5630 20725 6000 20735
rect 6030 20795 6400 20880
rect 6030 20735 6034 20795
rect 6086 20735 6344 20795
rect 6396 20735 6400 20795
rect 6030 20725 6400 20735
rect 6430 20795 6800 20880
rect 6430 20735 6434 20795
rect 6486 20735 6744 20795
rect 6796 20735 6800 20795
rect 6430 20725 6800 20735
rect 6830 20795 7200 20880
rect 6830 20735 6834 20795
rect 6886 20735 7144 20795
rect 7196 20735 7200 20795
rect 6830 20725 7200 20735
rect 7230 20795 7600 20880
rect 7230 20735 7234 20795
rect 7286 20735 7544 20795
rect 7596 20735 7600 20795
rect 7230 20725 7600 20735
rect 7630 20795 8000 20880
rect 7630 20735 7634 20795
rect 7686 20735 7944 20795
rect 7996 20735 8000 20795
rect 7630 20725 8000 20735
rect 8030 20795 8400 20880
rect 8030 20735 8034 20795
rect 8086 20735 8344 20795
rect 8396 20735 8400 20795
rect 8030 20725 8400 20735
rect 8430 20795 8800 20880
rect 8430 20735 8434 20795
rect 8486 20735 8744 20795
rect 8796 20735 8800 20795
rect 8430 20725 8800 20735
rect 8830 20795 9200 20880
rect 8830 20735 8834 20795
rect 8886 20735 9144 20795
rect 9196 20735 9200 20795
rect 8830 20725 9200 20735
rect 9230 20795 9600 20880
rect 9230 20735 9234 20795
rect 9286 20735 9544 20795
rect 9596 20735 9600 20795
rect 9230 20725 9600 20735
rect 9630 20795 10000 20880
rect 9630 20735 9634 20795
rect 9686 20735 9944 20795
rect 9996 20735 10000 20795
rect 9630 20725 10000 20735
rect 10030 20795 10400 20880
rect 10030 20735 10034 20795
rect 10086 20735 10344 20795
rect 10396 20735 10400 20795
rect 10030 20725 10400 20735
rect 10430 20795 10800 20880
rect 10430 20735 10434 20795
rect 10486 20735 10744 20795
rect 10796 20735 10800 20795
rect 10430 20725 10800 20735
rect 10830 20795 11200 20880
rect 10830 20735 10834 20795
rect 10886 20735 11144 20795
rect 11196 20735 11200 20795
rect 10830 20725 11200 20735
rect 11230 20795 11600 20880
rect 11230 20735 11234 20795
rect 11286 20735 11544 20795
rect 11596 20735 11600 20795
rect 11230 20725 11600 20735
rect 11630 20795 12000 20880
rect 11630 20735 11634 20795
rect 11686 20735 11944 20795
rect 11996 20735 12000 20795
rect 11630 20725 12000 20735
rect 12030 20795 12400 20880
rect 12030 20735 12034 20795
rect 12086 20735 12344 20795
rect 12396 20735 12400 20795
rect 12030 20725 12400 20735
rect 12430 20795 12800 20880
rect 12430 20735 12434 20795
rect 12486 20735 12744 20795
rect 12796 20735 12800 20795
rect 12430 20725 12800 20735
rect 12830 20795 13200 20880
rect 12830 20735 12834 20795
rect 12886 20735 13144 20795
rect 13196 20735 13200 20795
rect 12830 20725 13200 20735
rect -330 20695 -324 20725
rect 30 20695 70 20725
rect 430 20695 470 20725
rect 830 20695 870 20725
rect 1230 20695 1270 20725
rect 1630 20695 1670 20725
rect 2030 20695 2070 20725
rect 2430 20695 2470 20725
rect 2830 20695 2870 20725
rect 3230 20695 3270 20725
rect 3630 20695 3670 20725
rect 4030 20695 4070 20725
rect 4430 20695 4470 20725
rect 4830 20695 4870 20725
rect 5230 20695 5270 20725
rect 5630 20695 5670 20725
rect 6030 20695 6070 20725
rect 6430 20695 6470 20725
rect 6830 20695 6870 20725
rect 7230 20695 7270 20725
rect 7630 20695 7670 20725
rect 8030 20695 8070 20725
rect 8430 20695 8470 20725
rect 8830 20695 8870 20725
rect 9230 20695 9270 20725
rect 9630 20695 9670 20725
rect 10030 20695 10070 20725
rect 10430 20695 10470 20725
rect 10830 20695 10870 20725
rect 11230 20695 11270 20725
rect 11630 20695 11670 20725
rect 12030 20695 12070 20725
rect 12430 20695 12470 20725
rect -330 20685 0 20695
rect -314 20625 -56 20685
rect -4 20625 0 20685
rect -330 20425 0 20625
rect -314 20365 -56 20425
rect -4 20365 0 20425
rect -330 20355 0 20365
rect 30 20685 400 20695
rect 30 20625 34 20685
rect 86 20625 344 20685
rect 396 20625 400 20685
rect 30 20550 400 20625
rect 430 20685 800 20695
rect 430 20625 434 20685
rect 486 20625 744 20685
rect 796 20625 800 20685
rect 430 20550 800 20625
rect 830 20685 1200 20695
rect 830 20625 834 20685
rect 886 20625 1144 20685
rect 1196 20625 1200 20685
rect 830 20550 1200 20625
rect 1230 20685 1600 20695
rect 1230 20625 1234 20685
rect 1286 20625 1544 20685
rect 1596 20625 1600 20685
rect 1230 20550 1600 20625
rect 1630 20685 2000 20695
rect 1630 20625 1634 20685
rect 1686 20625 1944 20685
rect 1996 20625 2000 20685
rect 1630 20550 2000 20625
rect 2030 20685 2400 20695
rect 2030 20625 2034 20685
rect 2086 20625 2344 20685
rect 2396 20625 2400 20685
rect 2030 20550 2400 20625
rect 2430 20685 2800 20695
rect 2430 20625 2434 20685
rect 2486 20625 2744 20685
rect 2796 20625 2800 20685
rect 2430 20550 2800 20625
rect 2830 20685 3200 20695
rect 2830 20625 2834 20685
rect 2886 20625 3144 20685
rect 3196 20625 3200 20685
rect 2830 20550 3200 20625
rect 3230 20685 3600 20695
rect 3230 20625 3234 20685
rect 3286 20625 3544 20685
rect 3596 20625 3600 20685
rect 3230 20550 3600 20625
rect 3630 20685 4000 20695
rect 3630 20625 3634 20685
rect 3686 20625 3944 20685
rect 3996 20625 4000 20685
rect 3630 20550 4000 20625
rect 4030 20685 4400 20695
rect 4030 20625 4034 20685
rect 4086 20625 4344 20685
rect 4396 20625 4400 20685
rect 4030 20550 4400 20625
rect 4430 20685 4800 20695
rect 4430 20625 4434 20685
rect 4486 20625 4744 20685
rect 4796 20625 4800 20685
rect 4430 20550 4800 20625
rect 4830 20685 5200 20695
rect 4830 20625 4834 20685
rect 4886 20625 5144 20685
rect 5196 20625 5200 20685
rect 4830 20550 5200 20625
rect 5230 20685 5600 20695
rect 5230 20625 5234 20685
rect 5286 20625 5544 20685
rect 5596 20625 5600 20685
rect 5230 20550 5600 20625
rect 5630 20685 6000 20695
rect 5630 20625 5634 20685
rect 5686 20625 5944 20685
rect 5996 20625 6000 20685
rect 5630 20550 6000 20625
rect 6030 20685 6400 20695
rect 6030 20625 6034 20685
rect 6086 20625 6344 20685
rect 6396 20625 6400 20685
rect 6030 20550 6400 20625
rect 6430 20685 6800 20695
rect 6430 20625 6434 20685
rect 6486 20625 6744 20685
rect 6796 20625 6800 20685
rect 6430 20550 6800 20625
rect 6830 20685 7200 20695
rect 6830 20625 6834 20685
rect 6886 20625 7144 20685
rect 7196 20625 7200 20685
rect 6830 20550 7200 20625
rect 7230 20685 7600 20695
rect 7230 20625 7234 20685
rect 7286 20625 7544 20685
rect 7596 20625 7600 20685
rect 7230 20550 7600 20625
rect 7630 20685 8000 20695
rect 7630 20625 7634 20685
rect 7686 20625 7944 20685
rect 7996 20625 8000 20685
rect 7630 20550 8000 20625
rect 8030 20685 8400 20695
rect 8030 20625 8034 20685
rect 8086 20625 8344 20685
rect 8396 20625 8400 20685
rect 8030 20550 8400 20625
rect 8430 20685 8800 20695
rect 8430 20625 8434 20685
rect 8486 20625 8744 20685
rect 8796 20625 8800 20685
rect 8430 20550 8800 20625
rect 8830 20685 9200 20695
rect 8830 20625 8834 20685
rect 8886 20625 9144 20685
rect 9196 20625 9200 20685
rect 8830 20550 9200 20625
rect 9230 20685 9600 20695
rect 9230 20625 9234 20685
rect 9286 20625 9544 20685
rect 9596 20625 9600 20685
rect 9230 20550 9600 20625
rect 9630 20685 10000 20695
rect 9630 20625 9634 20685
rect 9686 20625 9944 20685
rect 9996 20625 10000 20685
rect 9630 20550 10000 20625
rect 10030 20685 10400 20695
rect 10030 20625 10034 20685
rect 10086 20625 10344 20685
rect 10396 20625 10400 20685
rect 10030 20550 10400 20625
rect 10430 20685 10800 20695
rect 10430 20625 10434 20685
rect 10486 20625 10744 20685
rect 10796 20625 10800 20685
rect 10430 20550 10800 20625
rect 10830 20685 11200 20695
rect 10830 20625 10834 20685
rect 10886 20625 11144 20685
rect 11196 20625 11200 20685
rect 10830 20550 11200 20625
rect 11230 20685 11600 20695
rect 11230 20625 11234 20685
rect 11286 20625 11544 20685
rect 11596 20625 11600 20685
rect 11230 20550 11600 20625
rect 11630 20685 12000 20695
rect 11630 20625 11634 20685
rect 11686 20625 11944 20685
rect 11996 20625 12000 20685
rect 11630 20550 12000 20625
rect 12030 20685 12400 20695
rect 12030 20625 12034 20685
rect 12086 20625 12344 20685
rect 12396 20625 12400 20685
rect 12030 20550 12400 20625
rect 12430 20685 12800 20695
rect 12430 20625 12434 20685
rect 12486 20625 12744 20685
rect 12796 20625 12800 20685
rect 12430 20550 12800 20625
rect 12830 20685 13200 20695
rect 12830 20625 12834 20685
rect 12886 20625 13144 20685
rect 13196 20625 13200 20685
rect 12830 20550 13200 20625
rect 30 20510 13200 20550
rect 30 20425 400 20510
rect 30 20365 34 20425
rect 86 20365 344 20425
rect 396 20365 400 20425
rect 30 20355 400 20365
rect 430 20425 800 20510
rect 430 20365 434 20425
rect 486 20365 744 20425
rect 796 20365 800 20425
rect 430 20355 800 20365
rect 830 20425 1200 20510
rect 830 20365 834 20425
rect 886 20365 1144 20425
rect 1196 20365 1200 20425
rect 830 20355 1200 20365
rect 1230 20425 1600 20510
rect 1230 20365 1234 20425
rect 1286 20365 1544 20425
rect 1596 20365 1600 20425
rect 1230 20355 1600 20365
rect 1630 20425 2000 20510
rect 1630 20365 1634 20425
rect 1686 20365 1944 20425
rect 1996 20365 2000 20425
rect 1630 20355 2000 20365
rect 2030 20425 2400 20510
rect 2030 20365 2034 20425
rect 2086 20365 2344 20425
rect 2396 20365 2400 20425
rect 2030 20355 2400 20365
rect 2430 20425 2800 20510
rect 2430 20365 2434 20425
rect 2486 20365 2744 20425
rect 2796 20365 2800 20425
rect 2430 20355 2800 20365
rect 2830 20425 3200 20510
rect 2830 20365 2834 20425
rect 2886 20365 3144 20425
rect 3196 20365 3200 20425
rect 2830 20355 3200 20365
rect 3230 20425 3600 20510
rect 3230 20365 3234 20425
rect 3286 20365 3544 20425
rect 3596 20365 3600 20425
rect 3230 20355 3600 20365
rect 3630 20425 4000 20510
rect 3630 20365 3634 20425
rect 3686 20365 3944 20425
rect 3996 20365 4000 20425
rect 3630 20355 4000 20365
rect 4030 20425 4400 20510
rect 4030 20365 4034 20425
rect 4086 20365 4344 20425
rect 4396 20365 4400 20425
rect 4030 20355 4400 20365
rect 4430 20425 4800 20510
rect 4430 20365 4434 20425
rect 4486 20365 4744 20425
rect 4796 20365 4800 20425
rect 4430 20355 4800 20365
rect 4830 20425 5200 20510
rect 4830 20365 4834 20425
rect 4886 20365 5144 20425
rect 5196 20365 5200 20425
rect 4830 20355 5200 20365
rect 5230 20425 5600 20510
rect 5230 20365 5234 20425
rect 5286 20365 5544 20425
rect 5596 20365 5600 20425
rect 5230 20355 5600 20365
rect 5630 20425 6000 20510
rect 5630 20365 5634 20425
rect 5686 20365 5944 20425
rect 5996 20365 6000 20425
rect 5630 20355 6000 20365
rect 6030 20425 6400 20510
rect 6030 20365 6034 20425
rect 6086 20365 6344 20425
rect 6396 20365 6400 20425
rect 6030 20355 6400 20365
rect 6430 20425 6800 20510
rect 6430 20365 6434 20425
rect 6486 20365 6744 20425
rect 6796 20365 6800 20425
rect 6430 20355 6800 20365
rect 6830 20425 7200 20510
rect 6830 20365 6834 20425
rect 6886 20365 7144 20425
rect 7196 20365 7200 20425
rect 6830 20355 7200 20365
rect 7230 20425 7600 20510
rect 7230 20365 7234 20425
rect 7286 20365 7544 20425
rect 7596 20365 7600 20425
rect 7230 20355 7600 20365
rect 7630 20425 8000 20510
rect 7630 20365 7634 20425
rect 7686 20365 7944 20425
rect 7996 20365 8000 20425
rect 7630 20355 8000 20365
rect 8030 20425 8400 20510
rect 8030 20365 8034 20425
rect 8086 20365 8344 20425
rect 8396 20365 8400 20425
rect 8030 20355 8400 20365
rect 8430 20425 8800 20510
rect 8430 20365 8434 20425
rect 8486 20365 8744 20425
rect 8796 20365 8800 20425
rect 8430 20355 8800 20365
rect 8830 20425 9200 20510
rect 8830 20365 8834 20425
rect 8886 20365 9144 20425
rect 9196 20365 9200 20425
rect 8830 20355 9200 20365
rect 9230 20425 9600 20510
rect 9230 20365 9234 20425
rect 9286 20365 9544 20425
rect 9596 20365 9600 20425
rect 9230 20355 9600 20365
rect 9630 20425 10000 20510
rect 9630 20365 9634 20425
rect 9686 20365 9944 20425
rect 9996 20365 10000 20425
rect 9630 20355 10000 20365
rect 10030 20425 10400 20510
rect 10030 20365 10034 20425
rect 10086 20365 10344 20425
rect 10396 20365 10400 20425
rect 10030 20355 10400 20365
rect 10430 20425 10800 20510
rect 10430 20365 10434 20425
rect 10486 20365 10744 20425
rect 10796 20365 10800 20425
rect 10430 20355 10800 20365
rect 10830 20425 11200 20510
rect 10830 20365 10834 20425
rect 10886 20365 11144 20425
rect 11196 20365 11200 20425
rect 10830 20355 11200 20365
rect 11230 20425 11600 20510
rect 11230 20365 11234 20425
rect 11286 20365 11544 20425
rect 11596 20365 11600 20425
rect 11230 20355 11600 20365
rect 11630 20425 12000 20510
rect 11630 20365 11634 20425
rect 11686 20365 11944 20425
rect 11996 20365 12000 20425
rect 11630 20355 12000 20365
rect 12030 20425 12400 20510
rect 12030 20365 12034 20425
rect 12086 20365 12344 20425
rect 12396 20365 12400 20425
rect 12030 20355 12400 20365
rect 12430 20425 12800 20510
rect 12430 20365 12434 20425
rect 12486 20365 12744 20425
rect 12796 20365 12800 20425
rect 12430 20355 12800 20365
rect 12830 20425 13200 20510
rect 12830 20365 12834 20425
rect 12886 20365 13144 20425
rect 13196 20365 13200 20425
rect 12830 20355 13200 20365
rect -330 20325 -324 20355
rect 30 20325 70 20355
rect 430 20325 470 20355
rect 830 20325 870 20355
rect 1230 20325 1270 20355
rect 1630 20325 1670 20355
rect 2030 20325 2070 20355
rect 2430 20325 2470 20355
rect 2830 20325 2870 20355
rect 3230 20325 3270 20355
rect 3630 20325 3670 20355
rect 4030 20325 4070 20355
rect 4430 20325 4470 20355
rect 4830 20325 4870 20355
rect 5230 20325 5270 20355
rect 5630 20325 5670 20355
rect 6030 20325 6070 20355
rect 6430 20325 6470 20355
rect 6830 20325 6870 20355
rect 7230 20325 7270 20355
rect 7630 20325 7670 20355
rect 8030 20325 8070 20355
rect 8430 20325 8470 20355
rect 8830 20325 8870 20355
rect 9230 20325 9270 20355
rect 9630 20325 9670 20355
rect 10030 20325 10070 20355
rect 10430 20325 10470 20355
rect 10830 20325 10870 20355
rect 11230 20325 11270 20355
rect 11630 20325 11670 20355
rect 12030 20325 12070 20355
rect 12430 20325 12470 20355
rect -330 20315 0 20325
rect -314 20255 -56 20315
rect -4 20255 0 20315
rect -330 20055 0 20255
rect -314 19995 -56 20055
rect -4 19995 0 20055
rect -330 19985 0 19995
rect 30 20315 400 20325
rect 30 20255 34 20315
rect 86 20255 344 20315
rect 396 20255 400 20315
rect 30 20180 400 20255
rect 430 20315 800 20325
rect 430 20255 434 20315
rect 486 20255 744 20315
rect 796 20255 800 20315
rect 430 20180 800 20255
rect 830 20315 1200 20325
rect 830 20255 834 20315
rect 886 20255 1144 20315
rect 1196 20255 1200 20315
rect 830 20180 1200 20255
rect 1230 20315 1600 20325
rect 1230 20255 1234 20315
rect 1286 20255 1544 20315
rect 1596 20255 1600 20315
rect 1230 20180 1600 20255
rect 1630 20315 2000 20325
rect 1630 20255 1634 20315
rect 1686 20255 1944 20315
rect 1996 20255 2000 20315
rect 1630 20180 2000 20255
rect 2030 20315 2400 20325
rect 2030 20255 2034 20315
rect 2086 20255 2344 20315
rect 2396 20255 2400 20315
rect 2030 20180 2400 20255
rect 2430 20315 2800 20325
rect 2430 20255 2434 20315
rect 2486 20255 2744 20315
rect 2796 20255 2800 20315
rect 2430 20180 2800 20255
rect 2830 20315 3200 20325
rect 2830 20255 2834 20315
rect 2886 20255 3144 20315
rect 3196 20255 3200 20315
rect 2830 20180 3200 20255
rect 3230 20315 3600 20325
rect 3230 20255 3234 20315
rect 3286 20255 3544 20315
rect 3596 20255 3600 20315
rect 3230 20180 3600 20255
rect 3630 20315 4000 20325
rect 3630 20255 3634 20315
rect 3686 20255 3944 20315
rect 3996 20255 4000 20315
rect 3630 20180 4000 20255
rect 4030 20315 4400 20325
rect 4030 20255 4034 20315
rect 4086 20255 4344 20315
rect 4396 20255 4400 20315
rect 4030 20180 4400 20255
rect 4430 20315 4800 20325
rect 4430 20255 4434 20315
rect 4486 20255 4744 20315
rect 4796 20255 4800 20315
rect 4430 20180 4800 20255
rect 4830 20315 5200 20325
rect 4830 20255 4834 20315
rect 4886 20255 5144 20315
rect 5196 20255 5200 20315
rect 4830 20180 5200 20255
rect 5230 20315 5600 20325
rect 5230 20255 5234 20315
rect 5286 20255 5544 20315
rect 5596 20255 5600 20315
rect 5230 20180 5600 20255
rect 5630 20315 6000 20325
rect 5630 20255 5634 20315
rect 5686 20255 5944 20315
rect 5996 20255 6000 20315
rect 5630 20180 6000 20255
rect 6030 20315 6400 20325
rect 6030 20255 6034 20315
rect 6086 20255 6344 20315
rect 6396 20255 6400 20315
rect 6030 20180 6400 20255
rect 6430 20315 6800 20325
rect 6430 20255 6434 20315
rect 6486 20255 6744 20315
rect 6796 20255 6800 20315
rect 6430 20180 6800 20255
rect 6830 20315 7200 20325
rect 6830 20255 6834 20315
rect 6886 20255 7144 20315
rect 7196 20255 7200 20315
rect 6830 20180 7200 20255
rect 7230 20315 7600 20325
rect 7230 20255 7234 20315
rect 7286 20255 7544 20315
rect 7596 20255 7600 20315
rect 7230 20180 7600 20255
rect 7630 20315 8000 20325
rect 7630 20255 7634 20315
rect 7686 20255 7944 20315
rect 7996 20255 8000 20315
rect 7630 20180 8000 20255
rect 8030 20315 8400 20325
rect 8030 20255 8034 20315
rect 8086 20255 8344 20315
rect 8396 20255 8400 20315
rect 8030 20180 8400 20255
rect 8430 20315 8800 20325
rect 8430 20255 8434 20315
rect 8486 20255 8744 20315
rect 8796 20255 8800 20315
rect 8430 20180 8800 20255
rect 8830 20315 9200 20325
rect 8830 20255 8834 20315
rect 8886 20255 9144 20315
rect 9196 20255 9200 20315
rect 8830 20180 9200 20255
rect 9230 20315 9600 20325
rect 9230 20255 9234 20315
rect 9286 20255 9544 20315
rect 9596 20255 9600 20315
rect 9230 20180 9600 20255
rect 9630 20315 10000 20325
rect 9630 20255 9634 20315
rect 9686 20255 9944 20315
rect 9996 20255 10000 20315
rect 9630 20180 10000 20255
rect 10030 20315 10400 20325
rect 10030 20255 10034 20315
rect 10086 20255 10344 20315
rect 10396 20255 10400 20315
rect 10030 20180 10400 20255
rect 10430 20315 10800 20325
rect 10430 20255 10434 20315
rect 10486 20255 10744 20315
rect 10796 20255 10800 20315
rect 10430 20180 10800 20255
rect 10830 20315 11200 20325
rect 10830 20255 10834 20315
rect 10886 20255 11144 20315
rect 11196 20255 11200 20315
rect 10830 20180 11200 20255
rect 11230 20315 11600 20325
rect 11230 20255 11234 20315
rect 11286 20255 11544 20315
rect 11596 20255 11600 20315
rect 11230 20180 11600 20255
rect 11630 20315 12000 20325
rect 11630 20255 11634 20315
rect 11686 20255 11944 20315
rect 11996 20255 12000 20315
rect 11630 20180 12000 20255
rect 12030 20315 12400 20325
rect 12030 20255 12034 20315
rect 12086 20255 12344 20315
rect 12396 20255 12400 20315
rect 12030 20180 12400 20255
rect 12430 20315 12800 20325
rect 12430 20255 12434 20315
rect 12486 20255 12744 20315
rect 12796 20255 12800 20315
rect 12430 20180 12800 20255
rect 12830 20315 13200 20325
rect 12830 20255 12834 20315
rect 12886 20255 13144 20315
rect 13196 20255 13200 20315
rect 12830 20180 13200 20255
rect 30 20140 13200 20180
rect 30 20055 400 20140
rect 30 19995 34 20055
rect 86 19995 344 20055
rect 396 19995 400 20055
rect 30 19985 400 19995
rect 430 20055 800 20140
rect 430 19995 434 20055
rect 486 19995 744 20055
rect 796 19995 800 20055
rect 430 19985 800 19995
rect 830 20055 1200 20140
rect 830 19995 834 20055
rect 886 19995 1144 20055
rect 1196 19995 1200 20055
rect 830 19985 1200 19995
rect 1230 20055 1600 20140
rect 1230 19995 1234 20055
rect 1286 19995 1544 20055
rect 1596 19995 1600 20055
rect 1230 19985 1600 19995
rect 1630 20055 2000 20140
rect 1630 19995 1634 20055
rect 1686 19995 1944 20055
rect 1996 19995 2000 20055
rect 1630 19985 2000 19995
rect 2030 20055 2400 20140
rect 2030 19995 2034 20055
rect 2086 19995 2344 20055
rect 2396 19995 2400 20055
rect 2030 19985 2400 19995
rect 2430 20055 2800 20140
rect 2430 19995 2434 20055
rect 2486 19995 2744 20055
rect 2796 19995 2800 20055
rect 2430 19985 2800 19995
rect 2830 20055 3200 20140
rect 2830 19995 2834 20055
rect 2886 19995 3144 20055
rect 3196 19995 3200 20055
rect 2830 19985 3200 19995
rect 3230 20055 3600 20140
rect 3230 19995 3234 20055
rect 3286 19995 3544 20055
rect 3596 19995 3600 20055
rect 3230 19985 3600 19995
rect 3630 20055 4000 20140
rect 3630 19995 3634 20055
rect 3686 19995 3944 20055
rect 3996 19995 4000 20055
rect 3630 19985 4000 19995
rect 4030 20055 4400 20140
rect 4030 19995 4034 20055
rect 4086 19995 4344 20055
rect 4396 19995 4400 20055
rect 4030 19985 4400 19995
rect 4430 20055 4800 20140
rect 4430 19995 4434 20055
rect 4486 19995 4744 20055
rect 4796 19995 4800 20055
rect 4430 19985 4800 19995
rect 4830 20055 5200 20140
rect 4830 19995 4834 20055
rect 4886 19995 5144 20055
rect 5196 19995 5200 20055
rect 4830 19985 5200 19995
rect 5230 20055 5600 20140
rect 5230 19995 5234 20055
rect 5286 19995 5544 20055
rect 5596 19995 5600 20055
rect 5230 19985 5600 19995
rect 5630 20055 6000 20140
rect 5630 19995 5634 20055
rect 5686 19995 5944 20055
rect 5996 19995 6000 20055
rect 5630 19985 6000 19995
rect 6030 20055 6400 20140
rect 6030 19995 6034 20055
rect 6086 19995 6344 20055
rect 6396 19995 6400 20055
rect 6030 19985 6400 19995
rect 6430 20055 6800 20140
rect 6430 19995 6434 20055
rect 6486 19995 6744 20055
rect 6796 19995 6800 20055
rect 6430 19985 6800 19995
rect 6830 20055 7200 20140
rect 6830 19995 6834 20055
rect 6886 19995 7144 20055
rect 7196 19995 7200 20055
rect 6830 19985 7200 19995
rect 7230 20055 7600 20140
rect 7230 19995 7234 20055
rect 7286 19995 7544 20055
rect 7596 19995 7600 20055
rect 7230 19985 7600 19995
rect 7630 20055 8000 20140
rect 7630 19995 7634 20055
rect 7686 19995 7944 20055
rect 7996 19995 8000 20055
rect 7630 19985 8000 19995
rect 8030 20055 8400 20140
rect 8030 19995 8034 20055
rect 8086 19995 8344 20055
rect 8396 19995 8400 20055
rect 8030 19985 8400 19995
rect 8430 20055 8800 20140
rect 8430 19995 8434 20055
rect 8486 19995 8744 20055
rect 8796 19995 8800 20055
rect 8430 19985 8800 19995
rect 8830 20055 9200 20140
rect 8830 19995 8834 20055
rect 8886 19995 9144 20055
rect 9196 19995 9200 20055
rect 8830 19985 9200 19995
rect 9230 20055 9600 20140
rect 9230 19995 9234 20055
rect 9286 19995 9544 20055
rect 9596 19995 9600 20055
rect 9230 19985 9600 19995
rect 9630 20055 10000 20140
rect 9630 19995 9634 20055
rect 9686 19995 9944 20055
rect 9996 19995 10000 20055
rect 9630 19985 10000 19995
rect 10030 20055 10400 20140
rect 10030 19995 10034 20055
rect 10086 19995 10344 20055
rect 10396 19995 10400 20055
rect 10030 19985 10400 19995
rect 10430 20055 10800 20140
rect 10430 19995 10434 20055
rect 10486 19995 10744 20055
rect 10796 19995 10800 20055
rect 10430 19985 10800 19995
rect 10830 20055 11200 20140
rect 10830 19995 10834 20055
rect 10886 19995 11144 20055
rect 11196 19995 11200 20055
rect 10830 19985 11200 19995
rect 11230 20055 11600 20140
rect 11230 19995 11234 20055
rect 11286 19995 11544 20055
rect 11596 19995 11600 20055
rect 11230 19985 11600 19995
rect 11630 20055 12000 20140
rect 11630 19995 11634 20055
rect 11686 19995 11944 20055
rect 11996 19995 12000 20055
rect 11630 19985 12000 19995
rect 12030 20055 12400 20140
rect 12030 19995 12034 20055
rect 12086 19995 12344 20055
rect 12396 19995 12400 20055
rect 12030 19985 12400 19995
rect 12430 20055 12800 20140
rect 12430 19995 12434 20055
rect 12486 19995 12744 20055
rect 12796 19995 12800 20055
rect 12430 19985 12800 19995
rect 12830 20055 13200 20140
rect 12830 19995 12834 20055
rect 12886 19995 13144 20055
rect 13196 19995 13200 20055
rect 12830 19985 13200 19995
rect -330 19955 -324 19985
rect 30 19955 70 19985
rect 430 19955 470 19985
rect 830 19955 870 19985
rect 1230 19955 1270 19985
rect 1630 19955 1670 19985
rect 2030 19955 2070 19985
rect 2430 19955 2470 19985
rect 2830 19955 2870 19985
rect 3230 19955 3270 19985
rect 3630 19955 3670 19985
rect 4030 19955 4070 19985
rect 4430 19955 4470 19985
rect 4830 19955 4870 19985
rect 5230 19955 5270 19985
rect 5630 19955 5670 19985
rect 6030 19955 6070 19985
rect 6430 19955 6470 19985
rect 6830 19955 6870 19985
rect 7230 19955 7270 19985
rect 7630 19955 7670 19985
rect 8030 19955 8070 19985
rect 8430 19955 8470 19985
rect 8830 19955 8870 19985
rect 9230 19955 9270 19985
rect 9630 19955 9670 19985
rect 10030 19955 10070 19985
rect 10430 19955 10470 19985
rect 10830 19955 10870 19985
rect 11230 19955 11270 19985
rect 11630 19955 11670 19985
rect 12030 19955 12070 19985
rect 12430 19955 12470 19985
rect -330 19945 0 19955
rect -314 19885 -56 19945
rect -4 19885 0 19945
rect -330 19685 0 19885
rect -314 19625 -56 19685
rect -4 19625 0 19685
rect -330 19615 0 19625
rect 30 19945 400 19955
rect 30 19885 34 19945
rect 86 19885 344 19945
rect 396 19885 400 19945
rect 30 19810 400 19885
rect 430 19945 800 19955
rect 430 19885 434 19945
rect 486 19885 744 19945
rect 796 19885 800 19945
rect 430 19810 800 19885
rect 830 19945 1200 19955
rect 830 19885 834 19945
rect 886 19885 1144 19945
rect 1196 19885 1200 19945
rect 830 19810 1200 19885
rect 1230 19945 1600 19955
rect 1230 19885 1234 19945
rect 1286 19885 1544 19945
rect 1596 19885 1600 19945
rect 1230 19810 1600 19885
rect 1630 19945 2000 19955
rect 1630 19885 1634 19945
rect 1686 19885 1944 19945
rect 1996 19885 2000 19945
rect 1630 19810 2000 19885
rect 2030 19945 2400 19955
rect 2030 19885 2034 19945
rect 2086 19885 2344 19945
rect 2396 19885 2400 19945
rect 2030 19810 2400 19885
rect 2430 19945 2800 19955
rect 2430 19885 2434 19945
rect 2486 19885 2744 19945
rect 2796 19885 2800 19945
rect 2430 19810 2800 19885
rect 2830 19945 3200 19955
rect 2830 19885 2834 19945
rect 2886 19885 3144 19945
rect 3196 19885 3200 19945
rect 2830 19810 3200 19885
rect 3230 19945 3600 19955
rect 3230 19885 3234 19945
rect 3286 19885 3544 19945
rect 3596 19885 3600 19945
rect 3230 19810 3600 19885
rect 3630 19945 4000 19955
rect 3630 19885 3634 19945
rect 3686 19885 3944 19945
rect 3996 19885 4000 19945
rect 3630 19810 4000 19885
rect 4030 19945 4400 19955
rect 4030 19885 4034 19945
rect 4086 19885 4344 19945
rect 4396 19885 4400 19945
rect 4030 19810 4400 19885
rect 4430 19945 4800 19955
rect 4430 19885 4434 19945
rect 4486 19885 4744 19945
rect 4796 19885 4800 19945
rect 4430 19810 4800 19885
rect 4830 19945 5200 19955
rect 4830 19885 4834 19945
rect 4886 19885 5144 19945
rect 5196 19885 5200 19945
rect 4830 19810 5200 19885
rect 5230 19945 5600 19955
rect 5230 19885 5234 19945
rect 5286 19885 5544 19945
rect 5596 19885 5600 19945
rect 5230 19810 5600 19885
rect 5630 19945 6000 19955
rect 5630 19885 5634 19945
rect 5686 19885 5944 19945
rect 5996 19885 6000 19945
rect 5630 19810 6000 19885
rect 6030 19945 6400 19955
rect 6030 19885 6034 19945
rect 6086 19885 6344 19945
rect 6396 19885 6400 19945
rect 6030 19810 6400 19885
rect 6430 19945 6800 19955
rect 6430 19885 6434 19945
rect 6486 19885 6744 19945
rect 6796 19885 6800 19945
rect 6430 19810 6800 19885
rect 6830 19945 7200 19955
rect 6830 19885 6834 19945
rect 6886 19885 7144 19945
rect 7196 19885 7200 19945
rect 6830 19810 7200 19885
rect 7230 19945 7600 19955
rect 7230 19885 7234 19945
rect 7286 19885 7544 19945
rect 7596 19885 7600 19945
rect 7230 19810 7600 19885
rect 7630 19945 8000 19955
rect 7630 19885 7634 19945
rect 7686 19885 7944 19945
rect 7996 19885 8000 19945
rect 7630 19810 8000 19885
rect 8030 19945 8400 19955
rect 8030 19885 8034 19945
rect 8086 19885 8344 19945
rect 8396 19885 8400 19945
rect 8030 19810 8400 19885
rect 8430 19945 8800 19955
rect 8430 19885 8434 19945
rect 8486 19885 8744 19945
rect 8796 19885 8800 19945
rect 8430 19810 8800 19885
rect 8830 19945 9200 19955
rect 8830 19885 8834 19945
rect 8886 19885 9144 19945
rect 9196 19885 9200 19945
rect 8830 19810 9200 19885
rect 9230 19945 9600 19955
rect 9230 19885 9234 19945
rect 9286 19885 9544 19945
rect 9596 19885 9600 19945
rect 9230 19810 9600 19885
rect 9630 19945 10000 19955
rect 9630 19885 9634 19945
rect 9686 19885 9944 19945
rect 9996 19885 10000 19945
rect 9630 19810 10000 19885
rect 10030 19945 10400 19955
rect 10030 19885 10034 19945
rect 10086 19885 10344 19945
rect 10396 19885 10400 19945
rect 10030 19810 10400 19885
rect 10430 19945 10800 19955
rect 10430 19885 10434 19945
rect 10486 19885 10744 19945
rect 10796 19885 10800 19945
rect 10430 19810 10800 19885
rect 10830 19945 11200 19955
rect 10830 19885 10834 19945
rect 10886 19885 11144 19945
rect 11196 19885 11200 19945
rect 10830 19810 11200 19885
rect 11230 19945 11600 19955
rect 11230 19885 11234 19945
rect 11286 19885 11544 19945
rect 11596 19885 11600 19945
rect 11230 19810 11600 19885
rect 11630 19945 12000 19955
rect 11630 19885 11634 19945
rect 11686 19885 11944 19945
rect 11996 19885 12000 19945
rect 11630 19810 12000 19885
rect 12030 19945 12400 19955
rect 12030 19885 12034 19945
rect 12086 19885 12344 19945
rect 12396 19885 12400 19945
rect 12030 19810 12400 19885
rect 12430 19945 12800 19955
rect 12430 19885 12434 19945
rect 12486 19885 12744 19945
rect 12796 19885 12800 19945
rect 12430 19810 12800 19885
rect 12830 19945 13200 19955
rect 12830 19885 12834 19945
rect 12886 19885 13144 19945
rect 13196 19885 13200 19945
rect 12830 19810 13200 19885
rect 30 19770 13200 19810
rect 30 19685 400 19770
rect 30 19625 34 19685
rect 86 19625 344 19685
rect 396 19625 400 19685
rect 30 19615 400 19625
rect 430 19685 800 19770
rect 430 19625 434 19685
rect 486 19625 744 19685
rect 796 19625 800 19685
rect 430 19615 800 19625
rect 830 19685 1200 19770
rect 830 19625 834 19685
rect 886 19625 1144 19685
rect 1196 19625 1200 19685
rect 830 19615 1200 19625
rect 1230 19685 1600 19770
rect 1230 19625 1234 19685
rect 1286 19625 1544 19685
rect 1596 19625 1600 19685
rect 1230 19615 1600 19625
rect 1630 19685 2000 19770
rect 1630 19625 1634 19685
rect 1686 19625 1944 19685
rect 1996 19625 2000 19685
rect 1630 19615 2000 19625
rect 2030 19685 2400 19770
rect 2030 19625 2034 19685
rect 2086 19625 2344 19685
rect 2396 19625 2400 19685
rect 2030 19615 2400 19625
rect 2430 19685 2800 19770
rect 2430 19625 2434 19685
rect 2486 19625 2744 19685
rect 2796 19625 2800 19685
rect 2430 19615 2800 19625
rect 2830 19685 3200 19770
rect 2830 19625 2834 19685
rect 2886 19625 3144 19685
rect 3196 19625 3200 19685
rect 2830 19615 3200 19625
rect 3230 19685 3600 19770
rect 3230 19625 3234 19685
rect 3286 19625 3544 19685
rect 3596 19625 3600 19685
rect 3230 19615 3600 19625
rect 3630 19685 4000 19770
rect 3630 19625 3634 19685
rect 3686 19625 3944 19685
rect 3996 19625 4000 19685
rect 3630 19615 4000 19625
rect 4030 19685 4400 19770
rect 4030 19625 4034 19685
rect 4086 19625 4344 19685
rect 4396 19625 4400 19685
rect 4030 19615 4400 19625
rect 4430 19685 4800 19770
rect 4430 19625 4434 19685
rect 4486 19625 4744 19685
rect 4796 19625 4800 19685
rect 4430 19615 4800 19625
rect 4830 19685 5200 19770
rect 4830 19625 4834 19685
rect 4886 19625 5144 19685
rect 5196 19625 5200 19685
rect 4830 19615 5200 19625
rect 5230 19685 5600 19770
rect 5230 19625 5234 19685
rect 5286 19625 5544 19685
rect 5596 19625 5600 19685
rect 5230 19615 5600 19625
rect 5630 19685 6000 19770
rect 5630 19625 5634 19685
rect 5686 19625 5944 19685
rect 5996 19625 6000 19685
rect 5630 19615 6000 19625
rect 6030 19685 6400 19770
rect 6030 19625 6034 19685
rect 6086 19625 6344 19685
rect 6396 19625 6400 19685
rect 6030 19615 6400 19625
rect 6430 19685 6800 19770
rect 6430 19625 6434 19685
rect 6486 19625 6744 19685
rect 6796 19625 6800 19685
rect 6430 19615 6800 19625
rect 6830 19685 7200 19770
rect 6830 19625 6834 19685
rect 6886 19625 7144 19685
rect 7196 19625 7200 19685
rect 6830 19615 7200 19625
rect 7230 19685 7600 19770
rect 7230 19625 7234 19685
rect 7286 19625 7544 19685
rect 7596 19625 7600 19685
rect 7230 19615 7600 19625
rect 7630 19685 8000 19770
rect 7630 19625 7634 19685
rect 7686 19625 7944 19685
rect 7996 19625 8000 19685
rect 7630 19615 8000 19625
rect 8030 19685 8400 19770
rect 8030 19625 8034 19685
rect 8086 19625 8344 19685
rect 8396 19625 8400 19685
rect 8030 19615 8400 19625
rect 8430 19685 8800 19770
rect 8430 19625 8434 19685
rect 8486 19625 8744 19685
rect 8796 19625 8800 19685
rect 8430 19615 8800 19625
rect 8830 19685 9200 19770
rect 8830 19625 8834 19685
rect 8886 19625 9144 19685
rect 9196 19625 9200 19685
rect 8830 19615 9200 19625
rect 9230 19685 9600 19770
rect 9230 19625 9234 19685
rect 9286 19625 9544 19685
rect 9596 19625 9600 19685
rect 9230 19615 9600 19625
rect 9630 19685 10000 19770
rect 9630 19625 9634 19685
rect 9686 19625 9944 19685
rect 9996 19625 10000 19685
rect 9630 19615 10000 19625
rect 10030 19685 10400 19770
rect 10030 19625 10034 19685
rect 10086 19625 10344 19685
rect 10396 19625 10400 19685
rect 10030 19615 10400 19625
rect 10430 19685 10800 19770
rect 10430 19625 10434 19685
rect 10486 19625 10744 19685
rect 10796 19625 10800 19685
rect 10430 19615 10800 19625
rect 10830 19685 11200 19770
rect 10830 19625 10834 19685
rect 10886 19625 11144 19685
rect 11196 19625 11200 19685
rect 10830 19615 11200 19625
rect 11230 19685 11600 19770
rect 11230 19625 11234 19685
rect 11286 19625 11544 19685
rect 11596 19625 11600 19685
rect 11230 19615 11600 19625
rect 11630 19685 12000 19770
rect 11630 19625 11634 19685
rect 11686 19625 11944 19685
rect 11996 19625 12000 19685
rect 11630 19615 12000 19625
rect 12030 19685 12400 19770
rect 12030 19625 12034 19685
rect 12086 19625 12344 19685
rect 12396 19625 12400 19685
rect 12030 19615 12400 19625
rect 12430 19685 12800 19770
rect 12430 19625 12434 19685
rect 12486 19625 12744 19685
rect 12796 19625 12800 19685
rect 12430 19615 12800 19625
rect 12830 19685 13200 19770
rect 12830 19625 12834 19685
rect 12886 19625 13144 19685
rect 13196 19625 13200 19685
rect 12830 19615 13200 19625
rect -330 19585 -324 19615
rect 30 19585 70 19615
rect 430 19585 470 19615
rect 830 19585 870 19615
rect 1230 19585 1270 19615
rect 1630 19585 1670 19615
rect 2030 19585 2070 19615
rect 2430 19585 2470 19615
rect 2830 19585 2870 19615
rect -330 19575 0 19585
rect -314 19515 -56 19575
rect -4 19515 0 19575
rect -330 19315 0 19515
rect -314 19255 -56 19315
rect -4 19255 0 19315
rect -330 19245 0 19255
rect 30 19575 400 19585
rect 30 19515 34 19575
rect 86 19515 344 19575
rect 396 19515 400 19575
rect 30 19440 400 19515
rect 430 19575 800 19585
rect 430 19515 434 19575
rect 486 19515 744 19575
rect 796 19515 800 19575
rect 430 19440 800 19515
rect 830 19575 1200 19585
rect 830 19515 834 19575
rect 886 19515 1144 19575
rect 1196 19515 1200 19575
rect 830 19440 1200 19515
rect 1230 19575 1600 19585
rect 1230 19515 1234 19575
rect 1286 19515 1544 19575
rect 1596 19515 1600 19575
rect 1230 19440 1600 19515
rect 1630 19575 2000 19585
rect 1630 19515 1634 19575
rect 1686 19515 1944 19575
rect 1996 19515 2000 19575
rect 1630 19440 2000 19515
rect 2030 19575 2400 19585
rect 2030 19515 2034 19575
rect 2086 19515 2344 19575
rect 2396 19515 2400 19575
rect 2030 19440 2400 19515
rect 2430 19575 2800 19585
rect 2430 19515 2434 19575
rect 2486 19515 2744 19575
rect 2796 19515 2800 19575
rect 2430 19440 2800 19515
rect 2830 19575 3200 19585
rect 2830 19515 2834 19575
rect 2886 19515 3144 19575
rect 3196 19515 3200 19575
rect 2830 19440 3200 19515
rect 30 19400 3200 19440
rect 30 19315 400 19400
rect 30 19255 34 19315
rect 86 19255 344 19315
rect 396 19255 400 19315
rect 30 19245 400 19255
rect 430 19315 800 19400
rect 430 19255 434 19315
rect 486 19255 744 19315
rect 796 19255 800 19315
rect 430 19245 800 19255
rect 830 19315 1200 19400
rect 830 19255 834 19315
rect 886 19255 1144 19315
rect 1196 19255 1200 19315
rect 830 19245 1200 19255
rect 1230 19315 1600 19400
rect 1230 19255 1234 19315
rect 1286 19255 1544 19315
rect 1596 19255 1600 19315
rect 1230 19245 1600 19255
rect 1630 19315 2000 19400
rect 1630 19255 1634 19315
rect 1686 19255 1944 19315
rect 1996 19255 2000 19315
rect 1630 19245 2000 19255
rect 2030 19315 2400 19400
rect 2030 19255 2034 19315
rect 2086 19255 2344 19315
rect 2396 19255 2400 19315
rect 2030 19245 2400 19255
rect 2430 19315 2800 19400
rect 2430 19255 2434 19315
rect 2486 19255 2744 19315
rect 2796 19255 2800 19315
rect 2430 19245 2800 19255
rect 2830 19315 3200 19400
rect 2830 19255 2834 19315
rect 2886 19255 3144 19315
rect 3196 19255 3200 19315
rect 2830 19245 3200 19255
rect 3230 19575 3600 19585
rect 3230 19515 3234 19575
rect 3286 19515 3544 19575
rect 3596 19515 3600 19575
rect 3230 19440 3600 19515
rect 3630 19575 4000 19585
rect 3630 19515 3634 19575
rect 3686 19515 3944 19575
rect 3996 19515 4000 19575
rect 3630 19440 4000 19515
rect 4030 19575 4400 19585
rect 4030 19515 4034 19575
rect 4086 19515 4344 19575
rect 4396 19515 4400 19575
rect 4030 19440 4400 19515
rect 4430 19575 4800 19585
rect 4430 19515 4434 19575
rect 4486 19515 4744 19575
rect 4796 19515 4800 19575
rect 4430 19440 4800 19515
rect 4830 19575 5200 19585
rect 4830 19515 4834 19575
rect 4886 19515 5144 19575
rect 5196 19515 5200 19575
rect 4830 19440 5200 19515
rect 5230 19575 5600 19585
rect 5230 19515 5234 19575
rect 5286 19515 5544 19575
rect 5596 19515 5600 19575
rect 5230 19440 5600 19515
rect 5630 19575 6000 19585
rect 5630 19515 5634 19575
rect 5686 19515 5944 19575
rect 5996 19515 6000 19575
rect 5630 19440 6000 19515
rect 6030 19575 6400 19585
rect 6030 19515 6034 19575
rect 6086 19515 6344 19575
rect 6396 19515 6400 19575
rect 6030 19440 6400 19515
rect 6430 19575 6800 19585
rect 6430 19515 6434 19575
rect 6486 19515 6744 19575
rect 6796 19515 6800 19575
rect 6430 19440 6800 19515
rect 6830 19575 7200 19585
rect 6830 19515 6834 19575
rect 6886 19515 7144 19575
rect 7196 19515 7200 19575
rect 6830 19440 7200 19515
rect 7230 19575 7600 19585
rect 7230 19515 7234 19575
rect 7286 19515 7544 19575
rect 7596 19515 7600 19575
rect 7230 19440 7600 19515
rect 7630 19575 8000 19585
rect 7630 19515 7634 19575
rect 7686 19515 7944 19575
rect 7996 19515 8000 19575
rect 7630 19440 8000 19515
rect 8030 19575 8400 19585
rect 8030 19515 8034 19575
rect 8086 19515 8344 19575
rect 8396 19515 8400 19575
rect 8030 19440 8400 19515
rect 8430 19575 8800 19585
rect 8430 19515 8434 19575
rect 8486 19515 8744 19575
rect 8796 19515 8800 19575
rect 8430 19440 8800 19515
rect 8830 19575 9200 19585
rect 8830 19515 8834 19575
rect 8886 19515 9144 19575
rect 9196 19515 9200 19575
rect 8830 19440 9200 19515
rect 9230 19575 9600 19585
rect 9230 19515 9234 19575
rect 9286 19515 9544 19575
rect 9596 19515 9600 19575
rect 9230 19440 9600 19515
rect 9630 19575 10000 19585
rect 9630 19515 9634 19575
rect 9686 19515 9944 19575
rect 9996 19515 10000 19575
rect 9630 19440 10000 19515
rect 10030 19575 10400 19585
rect 10030 19515 10034 19575
rect 10086 19515 10344 19575
rect 10396 19515 10400 19575
rect 10030 19440 10400 19515
rect 10430 19575 10800 19585
rect 10430 19515 10434 19575
rect 10486 19515 10744 19575
rect 10796 19515 10800 19575
rect 10430 19440 10800 19515
rect 10830 19575 11200 19585
rect 10830 19515 10834 19575
rect 10886 19515 11144 19575
rect 11196 19515 11200 19575
rect 10830 19440 11200 19515
rect 11230 19575 11600 19585
rect 11230 19515 11234 19575
rect 11286 19515 11544 19575
rect 11596 19515 11600 19575
rect 11230 19440 11600 19515
rect 11630 19575 12000 19585
rect 11630 19515 11634 19575
rect 11686 19515 11944 19575
rect 11996 19515 12000 19575
rect 11630 19440 12000 19515
rect 12030 19575 12400 19585
rect 12030 19515 12034 19575
rect 12086 19515 12344 19575
rect 12396 19515 12400 19575
rect 12030 19440 12400 19515
rect 12430 19575 12800 19585
rect 12430 19515 12434 19575
rect 12486 19515 12744 19575
rect 12796 19515 12800 19575
rect 12430 19440 12800 19515
rect 12830 19575 13200 19585
rect 12830 19515 12834 19575
rect 12886 19515 13144 19575
rect 13196 19515 13200 19575
rect 12830 19440 13200 19515
rect 3230 19400 13200 19440
rect 3230 19315 3600 19400
rect 3230 19255 3234 19315
rect 3286 19255 3544 19315
rect 3596 19255 3600 19315
rect 3230 19245 3600 19255
rect 3630 19315 4000 19400
rect 3630 19255 3634 19315
rect 3686 19255 3944 19315
rect 3996 19255 4000 19315
rect 3630 19245 4000 19255
rect 4030 19315 4400 19400
rect 4030 19255 4034 19315
rect 4086 19255 4344 19315
rect 4396 19255 4400 19315
rect 4030 19245 4400 19255
rect 4430 19315 4800 19400
rect 4430 19255 4434 19315
rect 4486 19255 4744 19315
rect 4796 19255 4800 19315
rect 4430 19245 4800 19255
rect 4830 19315 5200 19400
rect 4830 19255 4834 19315
rect 4886 19255 5144 19315
rect 5196 19255 5200 19315
rect 4830 19245 5200 19255
rect 5230 19315 5600 19400
rect 5230 19255 5234 19315
rect 5286 19255 5544 19315
rect 5596 19255 5600 19315
rect 5230 19245 5600 19255
rect 5630 19315 6000 19400
rect 5630 19255 5634 19315
rect 5686 19255 5944 19315
rect 5996 19255 6000 19315
rect 5630 19245 6000 19255
rect 6030 19315 6400 19400
rect 6030 19255 6034 19315
rect 6086 19255 6344 19315
rect 6396 19255 6400 19315
rect 6030 19245 6400 19255
rect 6430 19315 6800 19400
rect 6430 19255 6434 19315
rect 6486 19255 6744 19315
rect 6796 19255 6800 19315
rect 6430 19245 6800 19255
rect 6830 19315 7200 19400
rect 6830 19255 6834 19315
rect 6886 19255 7144 19315
rect 7196 19255 7200 19315
rect 6830 19245 7200 19255
rect 7230 19315 7600 19400
rect 7230 19255 7234 19315
rect 7286 19255 7544 19315
rect 7596 19255 7600 19315
rect 7230 19245 7600 19255
rect 7630 19315 8000 19400
rect 7630 19255 7634 19315
rect 7686 19255 7944 19315
rect 7996 19255 8000 19315
rect 7630 19245 8000 19255
rect 8030 19315 8400 19400
rect 8030 19255 8034 19315
rect 8086 19255 8344 19315
rect 8396 19255 8400 19315
rect 8030 19245 8400 19255
rect 8430 19315 8800 19400
rect 8430 19255 8434 19315
rect 8486 19255 8744 19315
rect 8796 19255 8800 19315
rect 8430 19245 8800 19255
rect 8830 19315 9200 19400
rect 8830 19255 8834 19315
rect 8886 19255 9144 19315
rect 9196 19255 9200 19315
rect 8830 19245 9200 19255
rect 9230 19315 9600 19400
rect 9230 19255 9234 19315
rect 9286 19255 9544 19315
rect 9596 19255 9600 19315
rect 9230 19245 9600 19255
rect 9630 19315 10000 19400
rect 9630 19255 9634 19315
rect 9686 19255 9944 19315
rect 9996 19255 10000 19315
rect 9630 19245 10000 19255
rect 10030 19315 10400 19400
rect 10030 19255 10034 19315
rect 10086 19255 10344 19315
rect 10396 19255 10400 19315
rect 10030 19245 10400 19255
rect 10430 19315 10800 19400
rect 10430 19255 10434 19315
rect 10486 19255 10744 19315
rect 10796 19255 10800 19315
rect 10430 19245 10800 19255
rect 10830 19315 11200 19400
rect 10830 19255 10834 19315
rect 10886 19255 11144 19315
rect 11196 19255 11200 19315
rect 10830 19245 11200 19255
rect 11230 19315 11600 19400
rect 11230 19255 11234 19315
rect 11286 19255 11544 19315
rect 11596 19255 11600 19315
rect 11230 19245 11600 19255
rect 11630 19315 12000 19400
rect 11630 19255 11634 19315
rect 11686 19255 11944 19315
rect 11996 19255 12000 19315
rect 11630 19245 12000 19255
rect 12030 19315 12400 19400
rect 12030 19255 12034 19315
rect 12086 19255 12344 19315
rect 12396 19255 12400 19315
rect 12030 19245 12400 19255
rect 12430 19315 12800 19400
rect 12430 19255 12434 19315
rect 12486 19255 12744 19315
rect 12796 19255 12800 19315
rect 12430 19245 12800 19255
rect 12830 19315 13200 19400
rect 12830 19255 12834 19315
rect 12886 19255 13144 19315
rect 13196 19255 13200 19315
rect 12830 19245 13200 19255
rect -330 19215 -324 19245
rect 30 19215 70 19245
rect 430 19215 470 19245
rect 830 19215 870 19245
rect 1230 19215 1270 19245
rect 1630 19215 1670 19245
rect 2030 19215 2070 19245
rect 2430 19215 2470 19245
rect 2830 19215 2870 19245
rect 3230 19215 3270 19245
rect 3630 19215 3670 19245
rect 4030 19215 4070 19245
rect 4430 19215 4470 19245
rect 4830 19215 4870 19245
rect 5230 19215 5270 19245
rect 5630 19215 5670 19245
rect 6030 19215 6070 19245
rect 6430 19215 6470 19245
rect 6830 19215 6870 19245
rect 7230 19215 7270 19245
rect 7630 19215 7670 19245
rect 8030 19215 8070 19245
rect 8430 19215 8470 19245
rect 8830 19215 8870 19245
rect 9230 19215 9270 19245
rect 9630 19215 9670 19245
rect 10030 19215 10070 19245
rect 10430 19215 10470 19245
rect 10830 19215 10870 19245
rect 11230 19215 11270 19245
rect 11630 19215 11670 19245
rect 12030 19215 12070 19245
rect 12430 19215 12470 19245
rect -330 19205 0 19215
rect -314 19145 -56 19205
rect -4 19145 0 19205
rect -330 18945 0 19145
rect -314 18885 -56 18945
rect -4 18885 0 18945
rect -330 18875 0 18885
rect 30 19205 400 19215
rect 30 19145 34 19205
rect 86 19145 344 19205
rect 396 19145 400 19205
rect 30 19070 400 19145
rect 430 19205 800 19215
rect 430 19145 434 19205
rect 486 19145 744 19205
rect 796 19145 800 19205
rect 430 19070 800 19145
rect 830 19205 1200 19215
rect 830 19145 834 19205
rect 886 19145 1144 19205
rect 1196 19145 1200 19205
rect 830 19070 1200 19145
rect 1230 19205 1600 19215
rect 1230 19145 1234 19205
rect 1286 19145 1544 19205
rect 1596 19145 1600 19205
rect 1230 19070 1600 19145
rect 1630 19205 2000 19215
rect 1630 19145 1634 19205
rect 1686 19145 1944 19205
rect 1996 19145 2000 19205
rect 1630 19070 2000 19145
rect 2030 19205 2400 19215
rect 2030 19145 2034 19205
rect 2086 19145 2344 19205
rect 2396 19145 2400 19205
rect 2030 19070 2400 19145
rect 2430 19205 2800 19215
rect 2430 19145 2434 19205
rect 2486 19145 2744 19205
rect 2796 19145 2800 19205
rect 2430 19070 2800 19145
rect 2830 19205 3200 19215
rect 2830 19145 2834 19205
rect 2886 19145 3144 19205
rect 3196 19145 3200 19205
rect 2830 19070 3200 19145
rect 30 19030 3200 19070
rect 30 18945 400 19030
rect 30 18885 34 18945
rect 86 18885 344 18945
rect 396 18885 400 18945
rect 30 18875 400 18885
rect 430 18945 800 19030
rect 430 18885 434 18945
rect 486 18885 744 18945
rect 796 18885 800 18945
rect 430 18875 800 18885
rect 830 18945 1200 19030
rect 830 18885 834 18945
rect 886 18885 1144 18945
rect 1196 18885 1200 18945
rect 830 18875 1200 18885
rect 1230 18945 1600 19030
rect 1230 18885 1234 18945
rect 1286 18885 1544 18945
rect 1596 18885 1600 18945
rect 1230 18875 1600 18885
rect 1630 18945 2000 19030
rect 1630 18885 1634 18945
rect 1686 18885 1944 18945
rect 1996 18885 2000 18945
rect 1630 18875 2000 18885
rect 2030 18945 2400 19030
rect 2030 18885 2034 18945
rect 2086 18885 2344 18945
rect 2396 18885 2400 18945
rect 2030 18875 2400 18885
rect 2430 18945 2800 19030
rect 2430 18885 2434 18945
rect 2486 18885 2744 18945
rect 2796 18885 2800 18945
rect 2430 18875 2800 18885
rect 2830 18945 3200 19030
rect 2830 18885 2834 18945
rect 2886 18885 3144 18945
rect 3196 18885 3200 18945
rect 2830 18875 3200 18885
rect 3230 19205 3600 19215
rect 3230 19145 3234 19205
rect 3286 19145 3544 19205
rect 3596 19145 3600 19205
rect 3230 19070 3600 19145
rect 3630 19205 4000 19215
rect 3630 19145 3634 19205
rect 3686 19145 3944 19205
rect 3996 19145 4000 19205
rect 3630 19070 4000 19145
rect 4030 19205 4400 19215
rect 4030 19145 4034 19205
rect 4086 19145 4344 19205
rect 4396 19145 4400 19205
rect 4030 19070 4400 19145
rect 4430 19205 4800 19215
rect 4430 19145 4434 19205
rect 4486 19145 4744 19205
rect 4796 19145 4800 19205
rect 4430 19070 4800 19145
rect 4830 19205 5200 19215
rect 4830 19145 4834 19205
rect 4886 19145 5144 19205
rect 5196 19145 5200 19205
rect 4830 19070 5200 19145
rect 5230 19205 5600 19215
rect 5230 19145 5234 19205
rect 5286 19145 5544 19205
rect 5596 19145 5600 19205
rect 5230 19070 5600 19145
rect 5630 19205 6000 19215
rect 5630 19145 5634 19205
rect 5686 19145 5944 19205
rect 5996 19145 6000 19205
rect 5630 19070 6000 19145
rect 6030 19205 6400 19215
rect 6030 19145 6034 19205
rect 6086 19145 6344 19205
rect 6396 19145 6400 19205
rect 6030 19070 6400 19145
rect 6430 19205 6800 19215
rect 6430 19145 6434 19205
rect 6486 19145 6744 19205
rect 6796 19145 6800 19205
rect 6430 19070 6800 19145
rect 6830 19205 7200 19215
rect 6830 19145 6834 19205
rect 6886 19145 7144 19205
rect 7196 19145 7200 19205
rect 6830 19070 7200 19145
rect 7230 19205 7600 19215
rect 7230 19145 7234 19205
rect 7286 19145 7544 19205
rect 7596 19145 7600 19205
rect 7230 19070 7600 19145
rect 7630 19205 8000 19215
rect 7630 19145 7634 19205
rect 7686 19145 7944 19205
rect 7996 19145 8000 19205
rect 7630 19070 8000 19145
rect 8030 19205 8400 19215
rect 8030 19145 8034 19205
rect 8086 19145 8344 19205
rect 8396 19145 8400 19205
rect 8030 19070 8400 19145
rect 8430 19205 8800 19215
rect 8430 19145 8434 19205
rect 8486 19145 8744 19205
rect 8796 19145 8800 19205
rect 8430 19070 8800 19145
rect 8830 19205 9200 19215
rect 8830 19145 8834 19205
rect 8886 19145 9144 19205
rect 9196 19145 9200 19205
rect 8830 19070 9200 19145
rect 9230 19205 9600 19215
rect 9230 19145 9234 19205
rect 9286 19145 9544 19205
rect 9596 19145 9600 19205
rect 9230 19070 9600 19145
rect 9630 19205 10000 19215
rect 9630 19145 9634 19205
rect 9686 19145 9944 19205
rect 9996 19145 10000 19205
rect 9630 19070 10000 19145
rect 10030 19205 10400 19215
rect 10030 19145 10034 19205
rect 10086 19145 10344 19205
rect 10396 19145 10400 19205
rect 10030 19070 10400 19145
rect 10430 19205 10800 19215
rect 10430 19145 10434 19205
rect 10486 19145 10744 19205
rect 10796 19145 10800 19205
rect 10430 19070 10800 19145
rect 10830 19205 11200 19215
rect 10830 19145 10834 19205
rect 10886 19145 11144 19205
rect 11196 19145 11200 19205
rect 10830 19070 11200 19145
rect 11230 19205 11600 19215
rect 11230 19145 11234 19205
rect 11286 19145 11544 19205
rect 11596 19145 11600 19205
rect 11230 19070 11600 19145
rect 11630 19205 12000 19215
rect 11630 19145 11634 19205
rect 11686 19145 11944 19205
rect 11996 19145 12000 19205
rect 11630 19070 12000 19145
rect 12030 19205 12400 19215
rect 12030 19145 12034 19205
rect 12086 19145 12344 19205
rect 12396 19145 12400 19205
rect 12030 19070 12400 19145
rect 12430 19205 12800 19215
rect 12430 19145 12434 19205
rect 12486 19145 12744 19205
rect 12796 19145 12800 19205
rect 12430 19070 12800 19145
rect 12830 19205 13200 19215
rect 12830 19145 12834 19205
rect 12886 19145 13144 19205
rect 13196 19145 13200 19205
rect 12830 19070 13200 19145
rect 3230 19030 13200 19070
rect 3230 18945 3600 19030
rect 3230 18885 3234 18945
rect 3286 18885 3544 18945
rect 3596 18885 3600 18945
rect 3230 18875 3600 18885
rect 3630 18945 4000 19030
rect 3630 18885 3634 18945
rect 3686 18885 3944 18945
rect 3996 18885 4000 18945
rect 3630 18875 4000 18885
rect 4030 18945 4400 19030
rect 4030 18885 4034 18945
rect 4086 18885 4344 18945
rect 4396 18885 4400 18945
rect 4030 18875 4400 18885
rect 4430 18945 4800 19030
rect 4430 18885 4434 18945
rect 4486 18885 4744 18945
rect 4796 18885 4800 18945
rect 4430 18875 4800 18885
rect 4830 18945 5200 19030
rect 4830 18885 4834 18945
rect 4886 18885 5144 18945
rect 5196 18885 5200 18945
rect 4830 18875 5200 18885
rect 5230 18945 5600 19030
rect 5230 18885 5234 18945
rect 5286 18885 5544 18945
rect 5596 18885 5600 18945
rect 5230 18875 5600 18885
rect 5630 18945 6000 19030
rect 5630 18885 5634 18945
rect 5686 18885 5944 18945
rect 5996 18885 6000 18945
rect 5630 18875 6000 18885
rect 6030 18945 6400 19030
rect 6030 18885 6034 18945
rect 6086 18885 6344 18945
rect 6396 18885 6400 18945
rect 6030 18875 6400 18885
rect 6430 18945 6800 19030
rect 6430 18885 6434 18945
rect 6486 18885 6744 18945
rect 6796 18885 6800 18945
rect 6430 18875 6800 18885
rect 6830 18945 7200 19030
rect 6830 18885 6834 18945
rect 6886 18885 7144 18945
rect 7196 18885 7200 18945
rect 6830 18875 7200 18885
rect 7230 18945 7600 19030
rect 7230 18885 7234 18945
rect 7286 18885 7544 18945
rect 7596 18885 7600 18945
rect 7230 18875 7600 18885
rect 7630 18945 8000 19030
rect 7630 18885 7634 18945
rect 7686 18885 7944 18945
rect 7996 18885 8000 18945
rect 7630 18875 8000 18885
rect 8030 18945 8400 19030
rect 8030 18885 8034 18945
rect 8086 18885 8344 18945
rect 8396 18885 8400 18945
rect 8030 18875 8400 18885
rect 8430 18945 8800 19030
rect 8430 18885 8434 18945
rect 8486 18885 8744 18945
rect 8796 18885 8800 18945
rect 8430 18875 8800 18885
rect 8830 18945 9200 19030
rect 8830 18885 8834 18945
rect 8886 18885 9144 18945
rect 9196 18885 9200 18945
rect 8830 18875 9200 18885
rect 9230 18945 9600 19030
rect 9230 18885 9234 18945
rect 9286 18885 9544 18945
rect 9596 18885 9600 18945
rect 9230 18875 9600 18885
rect 9630 18945 10000 19030
rect 9630 18885 9634 18945
rect 9686 18885 9944 18945
rect 9996 18885 10000 18945
rect 9630 18875 10000 18885
rect 10030 18945 10400 19030
rect 10030 18885 10034 18945
rect 10086 18885 10344 18945
rect 10396 18885 10400 18945
rect 10030 18875 10400 18885
rect 10430 18945 10800 19030
rect 10430 18885 10434 18945
rect 10486 18885 10744 18945
rect 10796 18885 10800 18945
rect 10430 18875 10800 18885
rect 10830 18945 11200 19030
rect 10830 18885 10834 18945
rect 10886 18885 11144 18945
rect 11196 18885 11200 18945
rect 10830 18875 11200 18885
rect 11230 18945 11600 19030
rect 11230 18885 11234 18945
rect 11286 18885 11544 18945
rect 11596 18885 11600 18945
rect 11230 18875 11600 18885
rect 11630 18945 12000 19030
rect 11630 18885 11634 18945
rect 11686 18885 11944 18945
rect 11996 18885 12000 18945
rect 11630 18875 12000 18885
rect 12030 18945 12400 19030
rect 12030 18885 12034 18945
rect 12086 18885 12344 18945
rect 12396 18885 12400 18945
rect 12030 18875 12400 18885
rect 12430 18945 12800 19030
rect 12430 18885 12434 18945
rect 12486 18885 12744 18945
rect 12796 18885 12800 18945
rect 12430 18875 12800 18885
rect 12830 18945 13200 19030
rect 12830 18885 12834 18945
rect 12886 18885 13144 18945
rect 13196 18885 13200 18945
rect 12830 18875 13200 18885
rect -330 18845 -324 18875
rect 30 18845 70 18875
rect 430 18845 470 18875
rect 830 18845 870 18875
rect 1230 18845 1270 18875
rect 1630 18845 1670 18875
rect 2030 18845 2070 18875
rect 2430 18845 2470 18875
rect 2830 18845 2870 18875
rect 3230 18845 3270 18875
rect 3630 18845 3670 18875
rect 4030 18845 4070 18875
rect 4430 18845 4470 18875
rect 4830 18845 4870 18875
rect 5230 18845 5270 18875
rect 5630 18845 5670 18875
rect 6030 18845 6070 18875
rect 6430 18845 6470 18875
rect 6830 18845 6870 18875
rect 7230 18845 7270 18875
rect 7630 18845 7670 18875
rect 8030 18845 8070 18875
rect 8430 18845 8470 18875
rect 8830 18845 8870 18875
rect 9230 18845 9270 18875
rect 9630 18845 9670 18875
rect 10030 18845 10070 18875
rect 10430 18845 10470 18875
rect 10830 18845 10870 18875
rect 11230 18845 11270 18875
rect 11630 18845 11670 18875
rect 12030 18845 12070 18875
rect 12430 18845 12470 18875
rect -330 18835 0 18845
rect -314 18775 -56 18835
rect -4 18775 0 18835
rect -330 18575 0 18775
rect -314 18515 -56 18575
rect -4 18515 0 18575
rect -330 18505 0 18515
rect 30 18835 400 18845
rect 30 18775 34 18835
rect 86 18775 344 18835
rect 396 18775 400 18835
rect 30 18700 400 18775
rect 430 18835 800 18845
rect 430 18775 434 18835
rect 486 18775 744 18835
rect 796 18775 800 18835
rect 430 18700 800 18775
rect 830 18835 1200 18845
rect 830 18775 834 18835
rect 886 18775 1144 18835
rect 1196 18775 1200 18835
rect 830 18700 1200 18775
rect 1230 18835 1600 18845
rect 1230 18775 1234 18835
rect 1286 18775 1544 18835
rect 1596 18775 1600 18835
rect 1230 18700 1600 18775
rect 1630 18835 2000 18845
rect 1630 18775 1634 18835
rect 1686 18775 1944 18835
rect 1996 18775 2000 18835
rect 1630 18700 2000 18775
rect 2030 18835 2400 18845
rect 2030 18775 2034 18835
rect 2086 18775 2344 18835
rect 2396 18775 2400 18835
rect 2030 18700 2400 18775
rect 2430 18835 2800 18845
rect 2430 18775 2434 18835
rect 2486 18775 2744 18835
rect 2796 18775 2800 18835
rect 2430 18700 2800 18775
rect 2830 18835 3200 18845
rect 2830 18775 2834 18835
rect 2886 18775 3144 18835
rect 3196 18775 3200 18835
rect 2830 18700 3200 18775
rect 30 18660 3200 18700
rect 30 18575 400 18660
rect 30 18515 34 18575
rect 86 18515 344 18575
rect 396 18515 400 18575
rect 30 18505 400 18515
rect 430 18575 800 18660
rect 430 18515 434 18575
rect 486 18515 744 18575
rect 796 18515 800 18575
rect 430 18505 800 18515
rect 830 18575 1200 18660
rect 830 18515 834 18575
rect 886 18515 1144 18575
rect 1196 18515 1200 18575
rect 830 18505 1200 18515
rect 1230 18575 1600 18660
rect 1230 18515 1234 18575
rect 1286 18515 1544 18575
rect 1596 18515 1600 18575
rect 1230 18505 1600 18515
rect 1630 18575 2000 18660
rect 1630 18515 1634 18575
rect 1686 18515 1944 18575
rect 1996 18515 2000 18575
rect 1630 18505 2000 18515
rect 2030 18575 2400 18660
rect 2030 18515 2034 18575
rect 2086 18515 2344 18575
rect 2396 18515 2400 18575
rect 2030 18505 2400 18515
rect 2430 18575 2800 18660
rect 2430 18515 2434 18575
rect 2486 18515 2744 18575
rect 2796 18515 2800 18575
rect 2430 18505 2800 18515
rect 2830 18575 3200 18660
rect 2830 18515 2834 18575
rect 2886 18515 3144 18575
rect 3196 18515 3200 18575
rect 2830 18505 3200 18515
rect 3230 18835 3600 18845
rect 3230 18775 3234 18835
rect 3286 18775 3544 18835
rect 3596 18775 3600 18835
rect 3230 18700 3600 18775
rect 3630 18835 4000 18845
rect 3630 18775 3634 18835
rect 3686 18775 3944 18835
rect 3996 18775 4000 18835
rect 3630 18700 4000 18775
rect 4030 18835 4400 18845
rect 4030 18775 4034 18835
rect 4086 18775 4344 18835
rect 4396 18775 4400 18835
rect 4030 18700 4400 18775
rect 4430 18835 4800 18845
rect 4430 18775 4434 18835
rect 4486 18775 4744 18835
rect 4796 18775 4800 18835
rect 4430 18700 4800 18775
rect 4830 18835 5200 18845
rect 4830 18775 4834 18835
rect 4886 18775 5144 18835
rect 5196 18775 5200 18835
rect 4830 18700 5200 18775
rect 5230 18835 5600 18845
rect 5230 18775 5234 18835
rect 5286 18775 5544 18835
rect 5596 18775 5600 18835
rect 5230 18700 5600 18775
rect 5630 18835 6000 18845
rect 5630 18775 5634 18835
rect 5686 18775 5944 18835
rect 5996 18775 6000 18835
rect 5630 18700 6000 18775
rect 6030 18835 6400 18845
rect 6030 18775 6034 18835
rect 6086 18775 6344 18835
rect 6396 18775 6400 18835
rect 6030 18700 6400 18775
rect 6430 18835 6800 18845
rect 6430 18775 6434 18835
rect 6486 18775 6744 18835
rect 6796 18775 6800 18835
rect 6430 18700 6800 18775
rect 6830 18835 7200 18845
rect 6830 18775 6834 18835
rect 6886 18775 7144 18835
rect 7196 18775 7200 18835
rect 6830 18700 7200 18775
rect 7230 18835 7600 18845
rect 7230 18775 7234 18835
rect 7286 18775 7544 18835
rect 7596 18775 7600 18835
rect 7230 18700 7600 18775
rect 7630 18835 8000 18845
rect 7630 18775 7634 18835
rect 7686 18775 7944 18835
rect 7996 18775 8000 18835
rect 7630 18700 8000 18775
rect 8030 18835 8400 18845
rect 8030 18775 8034 18835
rect 8086 18775 8344 18835
rect 8396 18775 8400 18835
rect 8030 18700 8400 18775
rect 8430 18835 8800 18845
rect 8430 18775 8434 18835
rect 8486 18775 8744 18835
rect 8796 18775 8800 18835
rect 8430 18700 8800 18775
rect 8830 18835 9200 18845
rect 8830 18775 8834 18835
rect 8886 18775 9144 18835
rect 9196 18775 9200 18835
rect 8830 18700 9200 18775
rect 9230 18835 9600 18845
rect 9230 18775 9234 18835
rect 9286 18775 9544 18835
rect 9596 18775 9600 18835
rect 9230 18700 9600 18775
rect 9630 18835 10000 18845
rect 9630 18775 9634 18835
rect 9686 18775 9944 18835
rect 9996 18775 10000 18835
rect 9630 18700 10000 18775
rect 10030 18835 10400 18845
rect 10030 18775 10034 18835
rect 10086 18775 10344 18835
rect 10396 18775 10400 18835
rect 10030 18700 10400 18775
rect 10430 18835 10800 18845
rect 10430 18775 10434 18835
rect 10486 18775 10744 18835
rect 10796 18775 10800 18835
rect 10430 18700 10800 18775
rect 10830 18835 11200 18845
rect 10830 18775 10834 18835
rect 10886 18775 11144 18835
rect 11196 18775 11200 18835
rect 10830 18700 11200 18775
rect 11230 18835 11600 18845
rect 11230 18775 11234 18835
rect 11286 18775 11544 18835
rect 11596 18775 11600 18835
rect 11230 18700 11600 18775
rect 11630 18835 12000 18845
rect 11630 18775 11634 18835
rect 11686 18775 11944 18835
rect 11996 18775 12000 18835
rect 11630 18700 12000 18775
rect 12030 18835 12400 18845
rect 12030 18775 12034 18835
rect 12086 18775 12344 18835
rect 12396 18775 12400 18835
rect 12030 18700 12400 18775
rect 12430 18835 12800 18845
rect 12430 18775 12434 18835
rect 12486 18775 12744 18835
rect 12796 18775 12800 18835
rect 12430 18700 12800 18775
rect 12830 18835 13200 18845
rect 12830 18775 12834 18835
rect 12886 18775 13144 18835
rect 13196 18775 13200 18835
rect 12830 18700 13200 18775
rect 3230 18660 13200 18700
rect 3230 18575 3600 18660
rect 3230 18515 3234 18575
rect 3286 18515 3544 18575
rect 3596 18515 3600 18575
rect 3230 18505 3600 18515
rect 3630 18575 4000 18660
rect 3630 18515 3634 18575
rect 3686 18515 3944 18575
rect 3996 18515 4000 18575
rect 3630 18505 4000 18515
rect 4030 18575 4400 18660
rect 4030 18515 4034 18575
rect 4086 18515 4344 18575
rect 4396 18515 4400 18575
rect 4030 18505 4400 18515
rect 4430 18575 4800 18660
rect 4430 18515 4434 18575
rect 4486 18515 4744 18575
rect 4796 18515 4800 18575
rect 4430 18505 4800 18515
rect 4830 18575 5200 18660
rect 4830 18515 4834 18575
rect 4886 18515 5144 18575
rect 5196 18515 5200 18575
rect 4830 18505 5200 18515
rect 5230 18575 5600 18660
rect 5230 18515 5234 18575
rect 5286 18515 5544 18575
rect 5596 18515 5600 18575
rect 5230 18505 5600 18515
rect 5630 18575 6000 18660
rect 5630 18515 5634 18575
rect 5686 18515 5944 18575
rect 5996 18515 6000 18575
rect 5630 18505 6000 18515
rect 6030 18575 6400 18660
rect 6030 18515 6034 18575
rect 6086 18515 6344 18575
rect 6396 18515 6400 18575
rect 6030 18505 6400 18515
rect 6430 18575 6800 18660
rect 6430 18515 6434 18575
rect 6486 18515 6744 18575
rect 6796 18515 6800 18575
rect 6430 18505 6800 18515
rect 6830 18575 7200 18660
rect 6830 18515 6834 18575
rect 6886 18515 7144 18575
rect 7196 18515 7200 18575
rect 6830 18505 7200 18515
rect 7230 18575 7600 18660
rect 7230 18515 7234 18575
rect 7286 18515 7544 18575
rect 7596 18515 7600 18575
rect 7230 18505 7600 18515
rect 7630 18575 8000 18660
rect 7630 18515 7634 18575
rect 7686 18515 7944 18575
rect 7996 18515 8000 18575
rect 7630 18505 8000 18515
rect 8030 18575 8400 18660
rect 8030 18515 8034 18575
rect 8086 18515 8344 18575
rect 8396 18515 8400 18575
rect 8030 18505 8400 18515
rect 8430 18575 8800 18660
rect 8430 18515 8434 18575
rect 8486 18515 8744 18575
rect 8796 18515 8800 18575
rect 8430 18505 8800 18515
rect 8830 18575 9200 18660
rect 8830 18515 8834 18575
rect 8886 18515 9144 18575
rect 9196 18515 9200 18575
rect 8830 18505 9200 18515
rect 9230 18575 9600 18660
rect 9230 18515 9234 18575
rect 9286 18515 9544 18575
rect 9596 18515 9600 18575
rect 9230 18505 9600 18515
rect 9630 18575 10000 18660
rect 9630 18515 9634 18575
rect 9686 18515 9944 18575
rect 9996 18515 10000 18575
rect 9630 18505 10000 18515
rect 10030 18575 10400 18660
rect 10030 18515 10034 18575
rect 10086 18515 10344 18575
rect 10396 18515 10400 18575
rect 10030 18505 10400 18515
rect 10430 18575 10800 18660
rect 10430 18515 10434 18575
rect 10486 18515 10744 18575
rect 10796 18515 10800 18575
rect 10430 18505 10800 18515
rect 10830 18575 11200 18660
rect 10830 18515 10834 18575
rect 10886 18515 11144 18575
rect 11196 18515 11200 18575
rect 10830 18505 11200 18515
rect 11230 18575 11600 18660
rect 11230 18515 11234 18575
rect 11286 18515 11544 18575
rect 11596 18515 11600 18575
rect 11230 18505 11600 18515
rect 11630 18575 12000 18660
rect 11630 18515 11634 18575
rect 11686 18515 11944 18575
rect 11996 18515 12000 18575
rect 11630 18505 12000 18515
rect 12030 18575 12400 18660
rect 12030 18515 12034 18575
rect 12086 18515 12344 18575
rect 12396 18515 12400 18575
rect 12030 18505 12400 18515
rect 12430 18575 12800 18660
rect 12430 18515 12434 18575
rect 12486 18515 12744 18575
rect 12796 18515 12800 18575
rect 12430 18505 12800 18515
rect 12830 18575 13200 18660
rect 12830 18515 12834 18575
rect 12886 18515 13144 18575
rect 13196 18515 13200 18575
rect 12830 18505 13200 18515
rect -330 18475 -324 18505
rect 30 18475 70 18505
rect 430 18475 470 18505
rect 830 18475 870 18505
rect 1230 18475 1270 18505
rect 1630 18475 1670 18505
rect 2030 18475 2070 18505
rect 2430 18475 2470 18505
rect 2830 18475 2870 18505
rect 3230 18475 3270 18505
rect 3630 18475 3670 18505
rect 4030 18475 4070 18505
rect 4430 18475 4470 18505
rect 4830 18475 4870 18505
rect 5230 18475 5270 18505
rect 5630 18475 5670 18505
rect 6030 18475 6070 18505
rect 6430 18475 6470 18505
rect 6830 18475 6870 18505
rect 7230 18475 7270 18505
rect 7630 18475 7670 18505
rect 8030 18475 8070 18505
rect 8430 18475 8470 18505
rect 8830 18475 8870 18505
rect 9230 18475 9270 18505
rect 9630 18475 9670 18505
rect 10030 18475 10070 18505
rect 10430 18475 10470 18505
rect 10830 18475 10870 18505
rect 11230 18475 11270 18505
rect 11630 18475 11670 18505
rect 12030 18475 12070 18505
rect 12430 18475 12470 18505
rect -330 18465 0 18475
rect -314 18405 -56 18465
rect -4 18405 0 18465
rect -330 18205 0 18405
rect -314 18145 -56 18205
rect -4 18145 0 18205
rect -330 18135 0 18145
rect 30 18465 400 18475
rect 30 18405 34 18465
rect 86 18405 344 18465
rect 396 18405 400 18465
rect 30 18330 400 18405
rect 430 18465 800 18475
rect 430 18405 434 18465
rect 486 18405 744 18465
rect 796 18405 800 18465
rect 430 18330 800 18405
rect 830 18465 1200 18475
rect 830 18405 834 18465
rect 886 18405 1144 18465
rect 1196 18405 1200 18465
rect 830 18330 1200 18405
rect 1230 18465 1600 18475
rect 1230 18405 1234 18465
rect 1286 18405 1544 18465
rect 1596 18405 1600 18465
rect 1230 18330 1600 18405
rect 1630 18465 2000 18475
rect 1630 18405 1634 18465
rect 1686 18405 1944 18465
rect 1996 18405 2000 18465
rect 1630 18330 2000 18405
rect 2030 18465 2400 18475
rect 2030 18405 2034 18465
rect 2086 18405 2344 18465
rect 2396 18405 2400 18465
rect 2030 18330 2400 18405
rect 2430 18465 2800 18475
rect 2430 18405 2434 18465
rect 2486 18405 2744 18465
rect 2796 18405 2800 18465
rect 2430 18330 2800 18405
rect 2830 18465 3200 18475
rect 2830 18405 2834 18465
rect 2886 18405 3144 18465
rect 3196 18405 3200 18465
rect 2830 18330 3200 18405
rect 30 18290 3200 18330
rect 30 18205 400 18290
rect 30 18145 34 18205
rect 86 18145 344 18205
rect 396 18145 400 18205
rect 30 18135 400 18145
rect 430 18205 800 18290
rect 430 18145 434 18205
rect 486 18145 744 18205
rect 796 18145 800 18205
rect 430 18135 800 18145
rect 830 18205 1200 18290
rect 830 18145 834 18205
rect 886 18145 1144 18205
rect 1196 18145 1200 18205
rect 830 18135 1200 18145
rect 1230 18205 1600 18290
rect 1230 18145 1234 18205
rect 1286 18145 1544 18205
rect 1596 18145 1600 18205
rect 1230 18135 1600 18145
rect 1630 18205 2000 18290
rect 1630 18145 1634 18205
rect 1686 18145 1944 18205
rect 1996 18145 2000 18205
rect 1630 18135 2000 18145
rect 2030 18205 2400 18290
rect 2030 18145 2034 18205
rect 2086 18145 2344 18205
rect 2396 18145 2400 18205
rect 2030 18135 2400 18145
rect 2430 18205 2800 18290
rect 2430 18145 2434 18205
rect 2486 18145 2744 18205
rect 2796 18145 2800 18205
rect 2430 18135 2800 18145
rect 2830 18205 3200 18290
rect 2830 18145 2834 18205
rect 2886 18145 3144 18205
rect 3196 18145 3200 18205
rect 2830 18135 3200 18145
rect 3230 18465 3600 18475
rect 3230 18405 3234 18465
rect 3286 18405 3544 18465
rect 3596 18405 3600 18465
rect 3230 18330 3600 18405
rect 3630 18465 4000 18475
rect 3630 18405 3634 18465
rect 3686 18405 3944 18465
rect 3996 18405 4000 18465
rect 3630 18330 4000 18405
rect 4030 18465 4400 18475
rect 4030 18405 4034 18465
rect 4086 18405 4344 18465
rect 4396 18405 4400 18465
rect 4030 18330 4400 18405
rect 4430 18465 4800 18475
rect 4430 18405 4434 18465
rect 4486 18405 4744 18465
rect 4796 18405 4800 18465
rect 4430 18330 4800 18405
rect 4830 18465 5200 18475
rect 4830 18405 4834 18465
rect 4886 18405 5144 18465
rect 5196 18405 5200 18465
rect 4830 18330 5200 18405
rect 5230 18465 5600 18475
rect 5230 18405 5234 18465
rect 5286 18405 5544 18465
rect 5596 18405 5600 18465
rect 5230 18330 5600 18405
rect 5630 18465 6000 18475
rect 5630 18405 5634 18465
rect 5686 18405 5944 18465
rect 5996 18405 6000 18465
rect 5630 18330 6000 18405
rect 6030 18465 6400 18475
rect 6030 18405 6034 18465
rect 6086 18405 6344 18465
rect 6396 18405 6400 18465
rect 6030 18330 6400 18405
rect 6430 18465 6800 18475
rect 6430 18405 6434 18465
rect 6486 18405 6744 18465
rect 6796 18405 6800 18465
rect 6430 18330 6800 18405
rect 6830 18465 7200 18475
rect 6830 18405 6834 18465
rect 6886 18405 7144 18465
rect 7196 18405 7200 18465
rect 6830 18330 7200 18405
rect 7230 18465 7600 18475
rect 7230 18405 7234 18465
rect 7286 18405 7544 18465
rect 7596 18405 7600 18465
rect 7230 18330 7600 18405
rect 7630 18465 8000 18475
rect 7630 18405 7634 18465
rect 7686 18405 7944 18465
rect 7996 18405 8000 18465
rect 7630 18330 8000 18405
rect 8030 18465 8400 18475
rect 8030 18405 8034 18465
rect 8086 18405 8344 18465
rect 8396 18405 8400 18465
rect 8030 18330 8400 18405
rect 8430 18465 8800 18475
rect 8430 18405 8434 18465
rect 8486 18405 8744 18465
rect 8796 18405 8800 18465
rect 8430 18330 8800 18405
rect 8830 18465 9200 18475
rect 8830 18405 8834 18465
rect 8886 18405 9144 18465
rect 9196 18405 9200 18465
rect 8830 18330 9200 18405
rect 9230 18465 9600 18475
rect 9230 18405 9234 18465
rect 9286 18405 9544 18465
rect 9596 18405 9600 18465
rect 9230 18330 9600 18405
rect 9630 18465 10000 18475
rect 9630 18405 9634 18465
rect 9686 18405 9944 18465
rect 9996 18405 10000 18465
rect 9630 18330 10000 18405
rect 10030 18465 10400 18475
rect 10030 18405 10034 18465
rect 10086 18405 10344 18465
rect 10396 18405 10400 18465
rect 10030 18330 10400 18405
rect 10430 18465 10800 18475
rect 10430 18405 10434 18465
rect 10486 18405 10744 18465
rect 10796 18405 10800 18465
rect 10430 18330 10800 18405
rect 10830 18465 11200 18475
rect 10830 18405 10834 18465
rect 10886 18405 11144 18465
rect 11196 18405 11200 18465
rect 10830 18330 11200 18405
rect 11230 18465 11600 18475
rect 11230 18405 11234 18465
rect 11286 18405 11544 18465
rect 11596 18405 11600 18465
rect 11230 18330 11600 18405
rect 11630 18465 12000 18475
rect 11630 18405 11634 18465
rect 11686 18405 11944 18465
rect 11996 18405 12000 18465
rect 11630 18330 12000 18405
rect 12030 18465 12400 18475
rect 12030 18405 12034 18465
rect 12086 18405 12344 18465
rect 12396 18405 12400 18465
rect 12030 18330 12400 18405
rect 12430 18465 12800 18475
rect 12430 18405 12434 18465
rect 12486 18405 12744 18465
rect 12796 18405 12800 18465
rect 12430 18330 12800 18405
rect 12830 18465 13200 18475
rect 12830 18405 12834 18465
rect 12886 18405 13144 18465
rect 13196 18405 13200 18465
rect 12830 18330 13200 18405
rect 3230 18290 13200 18330
rect 3230 18205 3600 18290
rect 3230 18145 3234 18205
rect 3286 18145 3544 18205
rect 3596 18145 3600 18205
rect 3230 18135 3600 18145
rect 3630 18205 4000 18290
rect 3630 18145 3634 18205
rect 3686 18145 3944 18205
rect 3996 18145 4000 18205
rect 3630 18135 4000 18145
rect 4030 18205 4400 18290
rect 4030 18145 4034 18205
rect 4086 18145 4344 18205
rect 4396 18145 4400 18205
rect 4030 18135 4400 18145
rect 4430 18205 4800 18290
rect 4430 18145 4434 18205
rect 4486 18145 4744 18205
rect 4796 18145 4800 18205
rect 4430 18135 4800 18145
rect 4830 18205 5200 18290
rect 4830 18145 4834 18205
rect 4886 18145 5144 18205
rect 5196 18145 5200 18205
rect 4830 18135 5200 18145
rect 5230 18205 5600 18290
rect 5230 18145 5234 18205
rect 5286 18145 5544 18205
rect 5596 18145 5600 18205
rect 5230 18135 5600 18145
rect 5630 18205 6000 18290
rect 5630 18145 5634 18205
rect 5686 18145 5944 18205
rect 5996 18145 6000 18205
rect 5630 18135 6000 18145
rect 6030 18205 6400 18290
rect 6030 18145 6034 18205
rect 6086 18145 6344 18205
rect 6396 18145 6400 18205
rect 6030 18135 6400 18145
rect 6430 18205 6800 18290
rect 6430 18145 6434 18205
rect 6486 18145 6744 18205
rect 6796 18145 6800 18205
rect 6430 18135 6800 18145
rect 6830 18205 7200 18290
rect 6830 18145 6834 18205
rect 6886 18145 7144 18205
rect 7196 18145 7200 18205
rect 6830 18135 7200 18145
rect 7230 18205 7600 18290
rect 7230 18145 7234 18205
rect 7286 18145 7544 18205
rect 7596 18145 7600 18205
rect 7230 18135 7600 18145
rect 7630 18205 8000 18290
rect 7630 18145 7634 18205
rect 7686 18145 7944 18205
rect 7996 18145 8000 18205
rect 7630 18135 8000 18145
rect 8030 18205 8400 18290
rect 8030 18145 8034 18205
rect 8086 18145 8344 18205
rect 8396 18145 8400 18205
rect 8030 18135 8400 18145
rect 8430 18205 8800 18290
rect 8430 18145 8434 18205
rect 8486 18145 8744 18205
rect 8796 18145 8800 18205
rect 8430 18135 8800 18145
rect 8830 18205 9200 18290
rect 8830 18145 8834 18205
rect 8886 18145 9144 18205
rect 9196 18145 9200 18205
rect 8830 18135 9200 18145
rect 9230 18205 9600 18290
rect 9230 18145 9234 18205
rect 9286 18145 9544 18205
rect 9596 18145 9600 18205
rect 9230 18135 9600 18145
rect 9630 18205 10000 18290
rect 9630 18145 9634 18205
rect 9686 18145 9944 18205
rect 9996 18145 10000 18205
rect 9630 18135 10000 18145
rect 10030 18205 10400 18290
rect 10030 18145 10034 18205
rect 10086 18145 10344 18205
rect 10396 18145 10400 18205
rect 10030 18135 10400 18145
rect 10430 18205 10800 18290
rect 10430 18145 10434 18205
rect 10486 18145 10744 18205
rect 10796 18145 10800 18205
rect 10430 18135 10800 18145
rect 10830 18205 11200 18290
rect 10830 18145 10834 18205
rect 10886 18145 11144 18205
rect 11196 18145 11200 18205
rect 10830 18135 11200 18145
rect 11230 18205 11600 18290
rect 11230 18145 11234 18205
rect 11286 18145 11544 18205
rect 11596 18145 11600 18205
rect 11230 18135 11600 18145
rect 11630 18205 12000 18290
rect 11630 18145 11634 18205
rect 11686 18145 11944 18205
rect 11996 18145 12000 18205
rect 11630 18135 12000 18145
rect 12030 18205 12400 18290
rect 12030 18145 12034 18205
rect 12086 18145 12344 18205
rect 12396 18145 12400 18205
rect 12030 18135 12400 18145
rect 12430 18205 12800 18290
rect 12430 18145 12434 18205
rect 12486 18145 12744 18205
rect 12796 18145 12800 18205
rect 12430 18135 12800 18145
rect 12830 18205 13200 18290
rect 12830 18145 12834 18205
rect 12886 18145 13144 18205
rect 13196 18145 13200 18205
rect 12830 18135 13200 18145
rect -330 18105 -324 18135
rect 30 18105 70 18135
rect 430 18105 470 18135
rect 830 18105 870 18135
rect 1230 18105 1270 18135
rect 1630 18105 1670 18135
rect 2030 18105 2070 18135
rect 2430 18105 2470 18135
rect 2830 18105 2870 18135
rect 3230 18105 3270 18135
rect 3630 18105 3670 18135
rect 4030 18105 4070 18135
rect 4430 18105 4470 18135
rect 4830 18105 4870 18135
rect 5230 18105 5270 18135
rect 5630 18105 5670 18135
rect 6030 18105 6070 18135
rect 6430 18105 6470 18135
rect 6830 18105 6870 18135
rect 7230 18105 7270 18135
rect 7630 18105 7670 18135
rect 8030 18105 8070 18135
rect 8430 18105 8470 18135
rect 8830 18105 8870 18135
rect 9230 18105 9270 18135
rect 9630 18105 9670 18135
rect 10030 18105 10070 18135
rect 10430 18105 10470 18135
rect 10830 18105 10870 18135
rect 11230 18105 11270 18135
rect 11630 18105 11670 18135
rect 12030 18105 12070 18135
rect 12430 18105 12470 18135
rect -330 18095 0 18105
rect -314 18035 -56 18095
rect -4 18035 0 18095
rect -330 17835 0 18035
rect -314 17775 -56 17835
rect -4 17775 0 17835
rect -330 17765 0 17775
rect 30 18095 400 18105
rect 30 18035 34 18095
rect 86 18035 344 18095
rect 396 18035 400 18095
rect 30 17960 400 18035
rect 430 18095 800 18105
rect 430 18035 434 18095
rect 486 18035 744 18095
rect 796 18035 800 18095
rect 430 17960 800 18035
rect 830 18095 1200 18105
rect 830 18035 834 18095
rect 886 18035 1144 18095
rect 1196 18035 1200 18095
rect 830 17960 1200 18035
rect 1230 18095 1600 18105
rect 1230 18035 1234 18095
rect 1286 18035 1544 18095
rect 1596 18035 1600 18095
rect 1230 17960 1600 18035
rect 1630 18095 2000 18105
rect 1630 18035 1634 18095
rect 1686 18035 1944 18095
rect 1996 18035 2000 18095
rect 1630 17960 2000 18035
rect 2030 18095 2400 18105
rect 2030 18035 2034 18095
rect 2086 18035 2344 18095
rect 2396 18035 2400 18095
rect 2030 17960 2400 18035
rect 2430 18095 2800 18105
rect 2430 18035 2434 18095
rect 2486 18035 2744 18095
rect 2796 18035 2800 18095
rect 2430 17960 2800 18035
rect 2830 18095 3200 18105
rect 2830 18035 2834 18095
rect 2886 18035 3144 18095
rect 3196 18035 3200 18095
rect 2830 17960 3200 18035
rect 30 17920 3200 17960
rect 30 17835 400 17920
rect 30 17775 34 17835
rect 86 17775 344 17835
rect 396 17775 400 17835
rect 30 17765 400 17775
rect 430 17835 800 17920
rect 430 17775 434 17835
rect 486 17775 744 17835
rect 796 17775 800 17835
rect 430 17765 800 17775
rect 830 17835 1200 17920
rect 830 17775 834 17835
rect 886 17775 1144 17835
rect 1196 17775 1200 17835
rect 830 17765 1200 17775
rect 1230 17835 1600 17920
rect 1230 17775 1234 17835
rect 1286 17775 1544 17835
rect 1596 17775 1600 17835
rect 1230 17765 1600 17775
rect 1630 17835 2000 17920
rect 1630 17775 1634 17835
rect 1686 17775 1944 17835
rect 1996 17775 2000 17835
rect 1630 17765 2000 17775
rect 2030 17835 2400 17920
rect 2030 17775 2034 17835
rect 2086 17775 2344 17835
rect 2396 17775 2400 17835
rect 2030 17765 2400 17775
rect 2430 17835 2800 17920
rect 2430 17775 2434 17835
rect 2486 17775 2744 17835
rect 2796 17775 2800 17835
rect 2430 17765 2800 17775
rect 2830 17835 3200 17920
rect 2830 17775 2834 17835
rect 2886 17775 3144 17835
rect 3196 17775 3200 17835
rect 2830 17765 3200 17775
rect 3230 18095 3600 18105
rect 3230 18035 3234 18095
rect 3286 18035 3544 18095
rect 3596 18035 3600 18095
rect 3230 17960 3600 18035
rect 3630 18095 4000 18105
rect 3630 18035 3634 18095
rect 3686 18035 3944 18095
rect 3996 18035 4000 18095
rect 3630 17960 4000 18035
rect 4030 18095 4400 18105
rect 4030 18035 4034 18095
rect 4086 18035 4344 18095
rect 4396 18035 4400 18095
rect 4030 17960 4400 18035
rect 4430 18095 4800 18105
rect 4430 18035 4434 18095
rect 4486 18035 4744 18095
rect 4796 18035 4800 18095
rect 4430 17960 4800 18035
rect 4830 18095 5200 18105
rect 4830 18035 4834 18095
rect 4886 18035 5144 18095
rect 5196 18035 5200 18095
rect 4830 17960 5200 18035
rect 5230 18095 5600 18105
rect 5230 18035 5234 18095
rect 5286 18035 5544 18095
rect 5596 18035 5600 18095
rect 5230 17960 5600 18035
rect 5630 18095 6000 18105
rect 5630 18035 5634 18095
rect 5686 18035 5944 18095
rect 5996 18035 6000 18095
rect 5630 17960 6000 18035
rect 6030 18095 6400 18105
rect 6030 18035 6034 18095
rect 6086 18035 6344 18095
rect 6396 18035 6400 18095
rect 6030 17960 6400 18035
rect 6430 18095 6800 18105
rect 6430 18035 6434 18095
rect 6486 18035 6744 18095
rect 6796 18035 6800 18095
rect 6430 17960 6800 18035
rect 6830 18095 7200 18105
rect 6830 18035 6834 18095
rect 6886 18035 7144 18095
rect 7196 18035 7200 18095
rect 6830 17960 7200 18035
rect 7230 18095 7600 18105
rect 7230 18035 7234 18095
rect 7286 18035 7544 18095
rect 7596 18035 7600 18095
rect 7230 17960 7600 18035
rect 7630 18095 8000 18105
rect 7630 18035 7634 18095
rect 7686 18035 7944 18095
rect 7996 18035 8000 18095
rect 7630 17960 8000 18035
rect 8030 18095 8400 18105
rect 8030 18035 8034 18095
rect 8086 18035 8344 18095
rect 8396 18035 8400 18095
rect 8030 17960 8400 18035
rect 8430 18095 8800 18105
rect 8430 18035 8434 18095
rect 8486 18035 8744 18095
rect 8796 18035 8800 18095
rect 8430 17960 8800 18035
rect 8830 18095 9200 18105
rect 8830 18035 8834 18095
rect 8886 18035 9144 18095
rect 9196 18035 9200 18095
rect 8830 17960 9200 18035
rect 9230 18095 9600 18105
rect 9230 18035 9234 18095
rect 9286 18035 9544 18095
rect 9596 18035 9600 18095
rect 9230 17960 9600 18035
rect 9630 18095 10000 18105
rect 9630 18035 9634 18095
rect 9686 18035 9944 18095
rect 9996 18035 10000 18095
rect 9630 17960 10000 18035
rect 10030 18095 10400 18105
rect 10030 18035 10034 18095
rect 10086 18035 10344 18095
rect 10396 18035 10400 18095
rect 10030 17960 10400 18035
rect 10430 18095 10800 18105
rect 10430 18035 10434 18095
rect 10486 18035 10744 18095
rect 10796 18035 10800 18095
rect 10430 17960 10800 18035
rect 10830 18095 11200 18105
rect 10830 18035 10834 18095
rect 10886 18035 11144 18095
rect 11196 18035 11200 18095
rect 10830 17960 11200 18035
rect 11230 18095 11600 18105
rect 11230 18035 11234 18095
rect 11286 18035 11544 18095
rect 11596 18035 11600 18095
rect 11230 17960 11600 18035
rect 11630 18095 12000 18105
rect 11630 18035 11634 18095
rect 11686 18035 11944 18095
rect 11996 18035 12000 18095
rect 11630 17960 12000 18035
rect 12030 18095 12400 18105
rect 12030 18035 12034 18095
rect 12086 18035 12344 18095
rect 12396 18035 12400 18095
rect 12030 17960 12400 18035
rect 12430 18095 12800 18105
rect 12430 18035 12434 18095
rect 12486 18035 12744 18095
rect 12796 18035 12800 18095
rect 12430 17960 12800 18035
rect 12830 18095 13200 18105
rect 12830 18035 12834 18095
rect 12886 18035 13144 18095
rect 13196 18035 13200 18095
rect 12830 17960 13200 18035
rect 3230 17920 13200 17960
rect 3230 17835 3600 17920
rect 3230 17775 3234 17835
rect 3286 17775 3544 17835
rect 3596 17775 3600 17835
rect 3230 17765 3600 17775
rect 3630 17835 4000 17920
rect 3630 17775 3634 17835
rect 3686 17775 3944 17835
rect 3996 17775 4000 17835
rect 3630 17765 4000 17775
rect 4030 17835 4400 17920
rect 4030 17775 4034 17835
rect 4086 17775 4344 17835
rect 4396 17775 4400 17835
rect 4030 17765 4400 17775
rect 4430 17835 4800 17920
rect 4430 17775 4434 17835
rect 4486 17775 4744 17835
rect 4796 17775 4800 17835
rect 4430 17765 4800 17775
rect 4830 17835 5200 17920
rect 4830 17775 4834 17835
rect 4886 17775 5144 17835
rect 5196 17775 5200 17835
rect 4830 17765 5200 17775
rect 5230 17835 5600 17920
rect 5230 17775 5234 17835
rect 5286 17775 5544 17835
rect 5596 17775 5600 17835
rect 5230 17765 5600 17775
rect 5630 17835 6000 17920
rect 5630 17775 5634 17835
rect 5686 17775 5944 17835
rect 5996 17775 6000 17835
rect 5630 17765 6000 17775
rect 6030 17835 6400 17920
rect 6030 17775 6034 17835
rect 6086 17775 6344 17835
rect 6396 17775 6400 17835
rect 6030 17765 6400 17775
rect 6430 17835 6800 17920
rect 6430 17775 6434 17835
rect 6486 17775 6744 17835
rect 6796 17775 6800 17835
rect 6430 17765 6800 17775
rect 6830 17835 7200 17920
rect 6830 17775 6834 17835
rect 6886 17775 7144 17835
rect 7196 17775 7200 17835
rect 6830 17765 7200 17775
rect 7230 17835 7600 17920
rect 7230 17775 7234 17835
rect 7286 17775 7544 17835
rect 7596 17775 7600 17835
rect 7230 17765 7600 17775
rect 7630 17835 8000 17920
rect 7630 17775 7634 17835
rect 7686 17775 7944 17835
rect 7996 17775 8000 17835
rect 7630 17765 8000 17775
rect 8030 17835 8400 17920
rect 8030 17775 8034 17835
rect 8086 17775 8344 17835
rect 8396 17775 8400 17835
rect 8030 17765 8400 17775
rect 8430 17835 8800 17920
rect 8430 17775 8434 17835
rect 8486 17775 8744 17835
rect 8796 17775 8800 17835
rect 8430 17765 8800 17775
rect 8830 17835 9200 17920
rect 8830 17775 8834 17835
rect 8886 17775 9144 17835
rect 9196 17775 9200 17835
rect 8830 17765 9200 17775
rect 9230 17835 9600 17920
rect 9230 17775 9234 17835
rect 9286 17775 9544 17835
rect 9596 17775 9600 17835
rect 9230 17765 9600 17775
rect 9630 17835 10000 17920
rect 9630 17775 9634 17835
rect 9686 17775 9944 17835
rect 9996 17775 10000 17835
rect 9630 17765 10000 17775
rect 10030 17835 10400 17920
rect 10030 17775 10034 17835
rect 10086 17775 10344 17835
rect 10396 17775 10400 17835
rect 10030 17765 10400 17775
rect 10430 17835 10800 17920
rect 10430 17775 10434 17835
rect 10486 17775 10744 17835
rect 10796 17775 10800 17835
rect 10430 17765 10800 17775
rect 10830 17835 11200 17920
rect 10830 17775 10834 17835
rect 10886 17775 11144 17835
rect 11196 17775 11200 17835
rect 10830 17765 11200 17775
rect 11230 17835 11600 17920
rect 11230 17775 11234 17835
rect 11286 17775 11544 17835
rect 11596 17775 11600 17835
rect 11230 17765 11600 17775
rect 11630 17835 12000 17920
rect 11630 17775 11634 17835
rect 11686 17775 11944 17835
rect 11996 17775 12000 17835
rect 11630 17765 12000 17775
rect 12030 17835 12400 17920
rect 12030 17775 12034 17835
rect 12086 17775 12344 17835
rect 12396 17775 12400 17835
rect 12030 17765 12400 17775
rect 12430 17835 12800 17920
rect 12430 17775 12434 17835
rect 12486 17775 12744 17835
rect 12796 17775 12800 17835
rect 12430 17765 12800 17775
rect 12830 17835 13200 17920
rect 12830 17775 12834 17835
rect 12886 17775 13144 17835
rect 13196 17775 13200 17835
rect 12830 17765 13200 17775
rect -330 17735 -324 17765
rect 30 17735 70 17765
rect 430 17735 470 17765
rect 830 17735 870 17765
rect 1230 17735 1270 17765
rect 1630 17735 1670 17765
rect 2030 17735 2070 17765
rect 2430 17735 2470 17765
rect 2830 17735 2870 17765
rect 3230 17735 3270 17765
rect 3630 17735 3670 17765
rect 4030 17735 4070 17765
rect 4430 17735 4470 17765
rect 4830 17735 4870 17765
rect 5230 17735 5270 17765
rect 5630 17735 5670 17765
rect 6030 17735 6070 17765
rect 6430 17735 6470 17765
rect 6830 17735 6870 17765
rect 7230 17735 7270 17765
rect 7630 17735 7670 17765
rect 8030 17735 8070 17765
rect 8430 17735 8470 17765
rect 8830 17735 8870 17765
rect 9230 17735 9270 17765
rect 9630 17735 9670 17765
rect 10030 17735 10070 17765
rect 10430 17735 10470 17765
rect 10830 17735 10870 17765
rect 11230 17735 11270 17765
rect 11630 17735 11670 17765
rect 12030 17735 12070 17765
rect 12430 17735 12470 17765
rect -330 17725 0 17735
rect -314 17665 -56 17725
rect -4 17665 0 17725
rect -330 17465 0 17665
rect -314 17405 -56 17465
rect -4 17405 0 17465
rect -330 17395 0 17405
rect 30 17725 400 17735
rect 30 17665 34 17725
rect 86 17665 344 17725
rect 396 17665 400 17725
rect 30 17590 400 17665
rect 430 17725 800 17735
rect 430 17665 434 17725
rect 486 17665 744 17725
rect 796 17665 800 17725
rect 430 17590 800 17665
rect 830 17725 1200 17735
rect 830 17665 834 17725
rect 886 17665 1144 17725
rect 1196 17665 1200 17725
rect 830 17590 1200 17665
rect 1230 17725 1600 17735
rect 1230 17665 1234 17725
rect 1286 17665 1544 17725
rect 1596 17665 1600 17725
rect 1230 17590 1600 17665
rect 1630 17725 2000 17735
rect 1630 17665 1634 17725
rect 1686 17665 1944 17725
rect 1996 17665 2000 17725
rect 1630 17590 2000 17665
rect 2030 17725 2400 17735
rect 2030 17665 2034 17725
rect 2086 17665 2344 17725
rect 2396 17665 2400 17725
rect 2030 17590 2400 17665
rect 2430 17725 2800 17735
rect 2430 17665 2434 17725
rect 2486 17665 2744 17725
rect 2796 17665 2800 17725
rect 2430 17590 2800 17665
rect 2830 17725 3200 17735
rect 2830 17665 2834 17725
rect 2886 17665 3144 17725
rect 3196 17665 3200 17725
rect 2830 17590 3200 17665
rect 30 17550 3200 17590
rect 30 17465 400 17550
rect 30 17405 34 17465
rect 86 17405 344 17465
rect 396 17405 400 17465
rect 30 17395 400 17405
rect 430 17465 800 17550
rect 430 17405 434 17465
rect 486 17405 744 17465
rect 796 17405 800 17465
rect 430 17395 800 17405
rect 830 17465 1200 17550
rect 830 17405 834 17465
rect 886 17405 1144 17465
rect 1196 17405 1200 17465
rect 830 17395 1200 17405
rect 1230 17465 1600 17550
rect 1230 17405 1234 17465
rect 1286 17405 1544 17465
rect 1596 17405 1600 17465
rect 1230 17395 1600 17405
rect 1630 17465 2000 17550
rect 1630 17405 1634 17465
rect 1686 17405 1944 17465
rect 1996 17405 2000 17465
rect 1630 17395 2000 17405
rect 2030 17465 2400 17550
rect 2030 17405 2034 17465
rect 2086 17405 2344 17465
rect 2396 17405 2400 17465
rect 2030 17395 2400 17405
rect 2430 17465 2800 17550
rect 2430 17405 2434 17465
rect 2486 17405 2744 17465
rect 2796 17405 2800 17465
rect 2430 17395 2800 17405
rect 2830 17465 3200 17550
rect 2830 17405 2834 17465
rect 2886 17405 3144 17465
rect 3196 17405 3200 17465
rect 2830 17395 3200 17405
rect 3230 17725 3600 17735
rect 3230 17665 3234 17725
rect 3286 17665 3544 17725
rect 3596 17665 3600 17725
rect 3230 17590 3600 17665
rect 3630 17725 4000 17735
rect 3630 17665 3634 17725
rect 3686 17665 3944 17725
rect 3996 17665 4000 17725
rect 3630 17590 4000 17665
rect 4030 17725 4400 17735
rect 4030 17665 4034 17725
rect 4086 17665 4344 17725
rect 4396 17665 4400 17725
rect 4030 17590 4400 17665
rect 4430 17725 4800 17735
rect 4430 17665 4434 17725
rect 4486 17665 4744 17725
rect 4796 17665 4800 17725
rect 4430 17590 4800 17665
rect 4830 17725 5200 17735
rect 4830 17665 4834 17725
rect 4886 17665 5144 17725
rect 5196 17665 5200 17725
rect 4830 17590 5200 17665
rect 5230 17725 5600 17735
rect 5230 17665 5234 17725
rect 5286 17665 5544 17725
rect 5596 17665 5600 17725
rect 5230 17590 5600 17665
rect 5630 17725 6000 17735
rect 5630 17665 5634 17725
rect 5686 17665 5944 17725
rect 5996 17665 6000 17725
rect 5630 17590 6000 17665
rect 6030 17725 6400 17735
rect 6030 17665 6034 17725
rect 6086 17665 6344 17725
rect 6396 17665 6400 17725
rect 6030 17590 6400 17665
rect 6430 17725 6800 17735
rect 6430 17665 6434 17725
rect 6486 17665 6744 17725
rect 6796 17665 6800 17725
rect 6430 17590 6800 17665
rect 6830 17725 7200 17735
rect 6830 17665 6834 17725
rect 6886 17665 7144 17725
rect 7196 17665 7200 17725
rect 6830 17590 7200 17665
rect 7230 17725 7600 17735
rect 7230 17665 7234 17725
rect 7286 17665 7544 17725
rect 7596 17665 7600 17725
rect 7230 17590 7600 17665
rect 7630 17725 8000 17735
rect 7630 17665 7634 17725
rect 7686 17665 7944 17725
rect 7996 17665 8000 17725
rect 7630 17590 8000 17665
rect 8030 17725 8400 17735
rect 8030 17665 8034 17725
rect 8086 17665 8344 17725
rect 8396 17665 8400 17725
rect 8030 17590 8400 17665
rect 8430 17725 8800 17735
rect 8430 17665 8434 17725
rect 8486 17665 8744 17725
rect 8796 17665 8800 17725
rect 8430 17590 8800 17665
rect 8830 17725 9200 17735
rect 8830 17665 8834 17725
rect 8886 17665 9144 17725
rect 9196 17665 9200 17725
rect 8830 17590 9200 17665
rect 9230 17725 9600 17735
rect 9230 17665 9234 17725
rect 9286 17665 9544 17725
rect 9596 17665 9600 17725
rect 9230 17590 9600 17665
rect 9630 17725 10000 17735
rect 9630 17665 9634 17725
rect 9686 17665 9944 17725
rect 9996 17665 10000 17725
rect 9630 17590 10000 17665
rect 10030 17725 10400 17735
rect 10030 17665 10034 17725
rect 10086 17665 10344 17725
rect 10396 17665 10400 17725
rect 10030 17590 10400 17665
rect 10430 17725 10800 17735
rect 10430 17665 10434 17725
rect 10486 17665 10744 17725
rect 10796 17665 10800 17725
rect 10430 17590 10800 17665
rect 10830 17725 11200 17735
rect 10830 17665 10834 17725
rect 10886 17665 11144 17725
rect 11196 17665 11200 17725
rect 10830 17590 11200 17665
rect 11230 17725 11600 17735
rect 11230 17665 11234 17725
rect 11286 17665 11544 17725
rect 11596 17665 11600 17725
rect 11230 17590 11600 17665
rect 11630 17725 12000 17735
rect 11630 17665 11634 17725
rect 11686 17665 11944 17725
rect 11996 17665 12000 17725
rect 11630 17590 12000 17665
rect 12030 17725 12400 17735
rect 12030 17665 12034 17725
rect 12086 17665 12344 17725
rect 12396 17665 12400 17725
rect 12030 17590 12400 17665
rect 12430 17725 12800 17735
rect 12430 17665 12434 17725
rect 12486 17665 12744 17725
rect 12796 17665 12800 17725
rect 12430 17590 12800 17665
rect 12830 17725 13200 17735
rect 12830 17665 12834 17725
rect 12886 17665 13144 17725
rect 13196 17665 13200 17725
rect 12830 17590 13200 17665
rect 3230 17550 13200 17590
rect 3230 17465 3600 17550
rect 3230 17405 3234 17465
rect 3286 17405 3544 17465
rect 3596 17405 3600 17465
rect 3230 17395 3600 17405
rect 3630 17465 4000 17550
rect 3630 17405 3634 17465
rect 3686 17405 3944 17465
rect 3996 17405 4000 17465
rect 3630 17395 4000 17405
rect 4030 17465 4400 17550
rect 4030 17405 4034 17465
rect 4086 17405 4344 17465
rect 4396 17405 4400 17465
rect 4030 17395 4400 17405
rect 4430 17465 4800 17550
rect 4430 17405 4434 17465
rect 4486 17405 4744 17465
rect 4796 17405 4800 17465
rect 4430 17395 4800 17405
rect 4830 17465 5200 17550
rect 4830 17405 4834 17465
rect 4886 17405 5144 17465
rect 5196 17405 5200 17465
rect 4830 17395 5200 17405
rect 5230 17465 5600 17550
rect 5230 17405 5234 17465
rect 5286 17405 5544 17465
rect 5596 17405 5600 17465
rect 5230 17395 5600 17405
rect 5630 17465 6000 17550
rect 5630 17405 5634 17465
rect 5686 17405 5944 17465
rect 5996 17405 6000 17465
rect 5630 17395 6000 17405
rect 6030 17465 6400 17550
rect 6030 17405 6034 17465
rect 6086 17405 6344 17465
rect 6396 17405 6400 17465
rect 6030 17395 6400 17405
rect 6430 17465 6800 17550
rect 6430 17405 6434 17465
rect 6486 17405 6744 17465
rect 6796 17405 6800 17465
rect 6430 17395 6800 17405
rect 6830 17465 7200 17550
rect 6830 17405 6834 17465
rect 6886 17405 7144 17465
rect 7196 17405 7200 17465
rect 6830 17395 7200 17405
rect 7230 17465 7600 17550
rect 7230 17405 7234 17465
rect 7286 17405 7544 17465
rect 7596 17405 7600 17465
rect 7230 17395 7600 17405
rect 7630 17465 8000 17550
rect 7630 17405 7634 17465
rect 7686 17405 7944 17465
rect 7996 17405 8000 17465
rect 7630 17395 8000 17405
rect 8030 17465 8400 17550
rect 8030 17405 8034 17465
rect 8086 17405 8344 17465
rect 8396 17405 8400 17465
rect 8030 17395 8400 17405
rect 8430 17465 8800 17550
rect 8430 17405 8434 17465
rect 8486 17405 8744 17465
rect 8796 17405 8800 17465
rect 8430 17395 8800 17405
rect 8830 17465 9200 17550
rect 8830 17405 8834 17465
rect 8886 17405 9144 17465
rect 9196 17405 9200 17465
rect 8830 17395 9200 17405
rect 9230 17465 9600 17550
rect 9230 17405 9234 17465
rect 9286 17405 9544 17465
rect 9596 17405 9600 17465
rect 9230 17395 9600 17405
rect 9630 17465 10000 17550
rect 9630 17405 9634 17465
rect 9686 17405 9944 17465
rect 9996 17405 10000 17465
rect 9630 17395 10000 17405
rect 10030 17465 10400 17550
rect 10030 17405 10034 17465
rect 10086 17405 10344 17465
rect 10396 17405 10400 17465
rect 10030 17395 10400 17405
rect 10430 17465 10800 17550
rect 10430 17405 10434 17465
rect 10486 17405 10744 17465
rect 10796 17405 10800 17465
rect 10430 17395 10800 17405
rect 10830 17465 11200 17550
rect 10830 17405 10834 17465
rect 10886 17405 11144 17465
rect 11196 17405 11200 17465
rect 10830 17395 11200 17405
rect 11230 17465 11600 17550
rect 11230 17405 11234 17465
rect 11286 17405 11544 17465
rect 11596 17405 11600 17465
rect 11230 17395 11600 17405
rect 11630 17465 12000 17550
rect 11630 17405 11634 17465
rect 11686 17405 11944 17465
rect 11996 17405 12000 17465
rect 11630 17395 12000 17405
rect 12030 17465 12400 17550
rect 12030 17405 12034 17465
rect 12086 17405 12344 17465
rect 12396 17405 12400 17465
rect 12030 17395 12400 17405
rect 12430 17465 12800 17550
rect 12430 17405 12434 17465
rect 12486 17405 12744 17465
rect 12796 17405 12800 17465
rect 12430 17395 12800 17405
rect 12830 17465 13200 17550
rect 12830 17405 12834 17465
rect 12886 17405 13144 17465
rect 13196 17405 13200 17465
rect 12830 17395 13200 17405
rect -330 17365 -324 17395
rect 30 17365 70 17395
rect 430 17365 470 17395
rect 830 17365 870 17395
rect 1230 17365 1270 17395
rect 1630 17365 1670 17395
rect 2030 17365 2070 17395
rect 2430 17365 2470 17395
rect 2830 17365 2870 17395
rect 3230 17365 3270 17395
rect 3630 17365 3670 17395
rect 4030 17365 4070 17395
rect 4430 17365 4470 17395
rect 4830 17365 4870 17395
rect 5230 17365 5270 17395
rect 5630 17365 5670 17395
rect -330 17355 0 17365
rect -314 17295 -56 17355
rect -4 17295 0 17355
rect -330 17095 0 17295
rect -314 17035 -56 17095
rect -4 17035 0 17095
rect -330 17025 0 17035
rect 30 17355 400 17365
rect 30 17295 34 17355
rect 86 17295 344 17355
rect 396 17295 400 17355
rect 30 17220 400 17295
rect 430 17355 800 17365
rect 430 17295 434 17355
rect 486 17295 744 17355
rect 796 17295 800 17355
rect 430 17220 800 17295
rect 830 17355 1200 17365
rect 830 17295 834 17355
rect 886 17295 1144 17355
rect 1196 17295 1200 17355
rect 830 17220 1200 17295
rect 1230 17355 1600 17365
rect 1230 17295 1234 17355
rect 1286 17295 1544 17355
rect 1596 17295 1600 17355
rect 1230 17220 1600 17295
rect 1630 17355 2000 17365
rect 1630 17295 1634 17355
rect 1686 17295 1944 17355
rect 1996 17295 2000 17355
rect 1630 17220 2000 17295
rect 2030 17355 2400 17365
rect 2030 17295 2034 17355
rect 2086 17295 2344 17355
rect 2396 17295 2400 17355
rect 2030 17220 2400 17295
rect 2430 17355 2800 17365
rect 2430 17295 2434 17355
rect 2486 17295 2744 17355
rect 2796 17295 2800 17355
rect 2430 17220 2800 17295
rect 2830 17355 3200 17365
rect 2830 17295 2834 17355
rect 2886 17295 3144 17355
rect 3196 17295 3200 17355
rect 2830 17220 3200 17295
rect 30 17180 3200 17220
rect 30 17095 400 17180
rect 30 17035 34 17095
rect 86 17035 344 17095
rect 396 17035 400 17095
rect 30 17025 400 17035
rect 430 17095 800 17180
rect 430 17035 434 17095
rect 486 17035 744 17095
rect 796 17035 800 17095
rect 430 17025 800 17035
rect 830 17095 1200 17180
rect 830 17035 834 17095
rect 886 17035 1144 17095
rect 1196 17035 1200 17095
rect 830 17025 1200 17035
rect 1230 17095 1600 17180
rect 1230 17035 1234 17095
rect 1286 17035 1544 17095
rect 1596 17035 1600 17095
rect 1230 17025 1600 17035
rect 1630 17095 2000 17180
rect 1630 17035 1634 17095
rect 1686 17035 1944 17095
rect 1996 17035 2000 17095
rect 1630 17025 2000 17035
rect 2030 17095 2400 17180
rect 2030 17035 2034 17095
rect 2086 17035 2344 17095
rect 2396 17035 2400 17095
rect 2030 17025 2400 17035
rect 2430 17095 2800 17180
rect 2430 17035 2434 17095
rect 2486 17035 2744 17095
rect 2796 17035 2800 17095
rect 2430 17025 2800 17035
rect 2830 17095 3200 17180
rect 2830 17035 2834 17095
rect 2886 17035 3144 17095
rect 3196 17035 3200 17095
rect 2830 17025 3200 17035
rect 3230 17355 3600 17365
rect 3230 17295 3234 17355
rect 3286 17295 3544 17355
rect 3596 17295 3600 17355
rect 3230 17220 3600 17295
rect 3630 17355 4000 17365
rect 3630 17295 3634 17355
rect 3686 17295 3944 17355
rect 3996 17295 4000 17355
rect 3630 17220 4000 17295
rect 4030 17355 4400 17365
rect 4030 17295 4034 17355
rect 4086 17295 4344 17355
rect 4396 17295 4400 17355
rect 4030 17220 4400 17295
rect 4430 17355 4800 17365
rect 4430 17295 4434 17355
rect 4486 17295 4744 17355
rect 4796 17295 4800 17355
rect 4430 17220 4800 17295
rect 4830 17355 5200 17365
rect 4830 17295 4834 17355
rect 4886 17295 5144 17355
rect 5196 17295 5200 17355
rect 4830 17220 5200 17295
rect 5230 17355 5600 17365
rect 5230 17295 5234 17355
rect 5286 17295 5544 17355
rect 5596 17295 5600 17355
rect 5230 17220 5600 17295
rect 5630 17355 6000 17365
rect 5630 17295 5634 17355
rect 5686 17295 5944 17355
rect 5996 17295 6000 17355
rect 5630 17220 6000 17295
rect 3230 17180 6000 17220
rect 3230 17095 3600 17180
rect 3230 17035 3234 17095
rect 3286 17035 3544 17095
rect 3596 17035 3600 17095
rect 3230 17025 3600 17035
rect 3630 17095 4000 17180
rect 3630 17035 3634 17095
rect 3686 17035 3944 17095
rect 3996 17035 4000 17095
rect 3630 17025 4000 17035
rect 4030 17095 4400 17180
rect 4030 17035 4034 17095
rect 4086 17035 4344 17095
rect 4396 17035 4400 17095
rect 4030 17025 4400 17035
rect 4430 17095 4800 17180
rect 4430 17035 4434 17095
rect 4486 17035 4744 17095
rect 4796 17035 4800 17095
rect 4430 17025 4800 17035
rect 4830 17095 5200 17180
rect 4830 17035 4834 17095
rect 4886 17035 5144 17095
rect 5196 17035 5200 17095
rect 4830 17025 5200 17035
rect 5230 17095 5600 17180
rect 5230 17035 5234 17095
rect 5286 17035 5544 17095
rect 5596 17035 5600 17095
rect 5230 17025 5600 17035
rect 5630 17095 6000 17180
rect 5630 17035 5634 17095
rect 5686 17035 5944 17095
rect 5996 17035 6000 17095
rect 5630 17025 6000 17035
rect 6030 17355 6400 17365
rect 6030 17295 6034 17355
rect 6086 17295 6344 17355
rect 6396 17295 6400 17355
rect 6030 17220 6400 17295
rect 6430 17355 6800 17365
rect 6430 17295 6434 17355
rect 6486 17295 6744 17355
rect 6796 17295 6800 17355
rect 6430 17220 6800 17295
rect 6830 17355 7200 17365
rect 6830 17295 6834 17355
rect 6886 17295 7144 17355
rect 7196 17295 7200 17355
rect 6830 17220 7200 17295
rect 7230 17355 7600 17365
rect 7230 17295 7234 17355
rect 7286 17295 7544 17355
rect 7596 17295 7600 17355
rect 7230 17220 7600 17295
rect 7630 17355 8000 17365
rect 7630 17295 7634 17355
rect 7686 17295 7944 17355
rect 7996 17295 8000 17355
rect 7630 17220 8000 17295
rect 8030 17355 8400 17365
rect 8030 17295 8034 17355
rect 8086 17295 8344 17355
rect 8396 17295 8400 17355
rect 8030 17220 8400 17295
rect 8430 17355 8800 17365
rect 8430 17295 8434 17355
rect 8486 17295 8744 17355
rect 8796 17295 8800 17355
rect 8430 17220 8800 17295
rect 8830 17355 9200 17365
rect 8830 17295 8834 17355
rect 8886 17295 9144 17355
rect 9196 17295 9200 17355
rect 8830 17220 9200 17295
rect 9230 17355 9600 17365
rect 9230 17295 9234 17355
rect 9286 17295 9544 17355
rect 9596 17295 9600 17355
rect 9230 17220 9600 17295
rect 9630 17355 10000 17365
rect 9630 17295 9634 17355
rect 9686 17295 9944 17355
rect 9996 17295 10000 17355
rect 9630 17220 10000 17295
rect 10030 17355 10400 17365
rect 10030 17295 10034 17355
rect 10086 17295 10344 17355
rect 10396 17295 10400 17355
rect 10030 17220 10400 17295
rect 10430 17355 10800 17365
rect 10430 17295 10434 17355
rect 10486 17295 10744 17355
rect 10796 17295 10800 17355
rect 10430 17220 10800 17295
rect 10830 17355 11200 17365
rect 10830 17295 10834 17355
rect 10886 17295 11144 17355
rect 11196 17295 11200 17355
rect 10830 17220 11200 17295
rect 11230 17355 11600 17365
rect 11230 17295 11234 17355
rect 11286 17295 11544 17355
rect 11596 17295 11600 17355
rect 11230 17220 11600 17295
rect 11630 17355 12000 17365
rect 11630 17295 11634 17355
rect 11686 17295 11944 17355
rect 11996 17295 12000 17355
rect 11630 17220 12000 17295
rect 12030 17355 12400 17365
rect 12030 17295 12034 17355
rect 12086 17295 12344 17355
rect 12396 17295 12400 17355
rect 12030 17220 12400 17295
rect 12430 17355 12800 17365
rect 12430 17295 12434 17355
rect 12486 17295 12744 17355
rect 12796 17295 12800 17355
rect 12430 17220 12800 17295
rect 12830 17355 13200 17365
rect 12830 17295 12834 17355
rect 12886 17295 13144 17355
rect 13196 17295 13200 17355
rect 12830 17220 13200 17295
rect 6030 17180 13200 17220
rect 6030 17095 6400 17180
rect 6030 17035 6034 17095
rect 6086 17035 6344 17095
rect 6396 17035 6400 17095
rect 6030 17025 6400 17035
rect 6430 17095 6800 17180
rect 6430 17035 6434 17095
rect 6486 17035 6744 17095
rect 6796 17035 6800 17095
rect 6430 17025 6800 17035
rect 6830 17095 7200 17180
rect 6830 17035 6834 17095
rect 6886 17035 7144 17095
rect 7196 17035 7200 17095
rect 6830 17025 7200 17035
rect 7230 17095 7600 17180
rect 7230 17035 7234 17095
rect 7286 17035 7544 17095
rect 7596 17035 7600 17095
rect 7230 17025 7600 17035
rect 7630 17095 8000 17180
rect 7630 17035 7634 17095
rect 7686 17035 7944 17095
rect 7996 17035 8000 17095
rect 7630 17025 8000 17035
rect 8030 17095 8400 17180
rect 8030 17035 8034 17095
rect 8086 17035 8344 17095
rect 8396 17035 8400 17095
rect 8030 17025 8400 17035
rect 8430 17095 8800 17180
rect 8430 17035 8434 17095
rect 8486 17035 8744 17095
rect 8796 17035 8800 17095
rect 8430 17025 8800 17035
rect 8830 17095 9200 17180
rect 8830 17035 8834 17095
rect 8886 17035 9144 17095
rect 9196 17035 9200 17095
rect 8830 17025 9200 17035
rect 9230 17095 9600 17180
rect 9230 17035 9234 17095
rect 9286 17035 9544 17095
rect 9596 17035 9600 17095
rect 9230 17025 9600 17035
rect 9630 17095 10000 17180
rect 9630 17035 9634 17095
rect 9686 17035 9944 17095
rect 9996 17035 10000 17095
rect 9630 17025 10000 17035
rect 10030 17095 10400 17180
rect 10030 17035 10034 17095
rect 10086 17035 10344 17095
rect 10396 17035 10400 17095
rect 10030 17025 10400 17035
rect 10430 17095 10800 17180
rect 10430 17035 10434 17095
rect 10486 17035 10744 17095
rect 10796 17035 10800 17095
rect 10430 17025 10800 17035
rect 10830 17095 11200 17180
rect 10830 17035 10834 17095
rect 10886 17035 11144 17095
rect 11196 17035 11200 17095
rect 10830 17025 11200 17035
rect 11230 17095 11600 17180
rect 11230 17035 11234 17095
rect 11286 17035 11544 17095
rect 11596 17035 11600 17095
rect 11230 17025 11600 17035
rect 11630 17095 12000 17180
rect 11630 17035 11634 17095
rect 11686 17035 11944 17095
rect 11996 17035 12000 17095
rect 11630 17025 12000 17035
rect 12030 17095 12400 17180
rect 12030 17035 12034 17095
rect 12086 17035 12344 17095
rect 12396 17035 12400 17095
rect 12030 17025 12400 17035
rect 12430 17095 12800 17180
rect 12430 17035 12434 17095
rect 12486 17035 12744 17095
rect 12796 17035 12800 17095
rect 12430 17025 12800 17035
rect 12830 17095 13200 17180
rect 12830 17035 12834 17095
rect 12886 17035 13144 17095
rect 13196 17035 13200 17095
rect 12830 17025 13200 17035
rect -330 16995 -324 17025
rect 30 16995 70 17025
rect 430 16995 470 17025
rect 830 16995 870 17025
rect 1230 16995 1270 17025
rect 1630 16995 1670 17025
rect 2030 16995 2070 17025
rect 2430 16995 2470 17025
rect 2830 16995 2870 17025
rect 3230 16995 3270 17025
rect 3630 16995 3670 17025
rect 4030 16995 4070 17025
rect 4430 16995 4470 17025
rect 4830 16995 4870 17025
rect 5230 16995 5270 17025
rect 5630 16995 5670 17025
rect 6030 16995 6070 17025
rect 6430 16995 6470 17025
rect 6830 16995 6870 17025
rect 7230 16995 7270 17025
rect 7630 16995 7670 17025
rect 8030 16995 8070 17025
rect 8430 16995 8470 17025
rect 8830 16995 8870 17025
rect 9230 16995 9270 17025
rect 9630 16995 9670 17025
rect 10030 16995 10070 17025
rect 10430 16995 10470 17025
rect 10830 16995 10870 17025
rect 11230 16995 11270 17025
rect 11630 16995 11670 17025
rect 12030 16995 12070 17025
rect 12430 16995 12470 17025
rect -330 16985 0 16995
rect -314 16925 -56 16985
rect -4 16925 0 16985
rect -330 16725 0 16925
rect -314 16665 -56 16725
rect -4 16665 0 16725
rect -330 16655 0 16665
rect 30 16985 400 16995
rect 30 16925 34 16985
rect 86 16925 344 16985
rect 396 16925 400 16985
rect 30 16850 400 16925
rect 430 16985 800 16995
rect 430 16925 434 16985
rect 486 16925 744 16985
rect 796 16925 800 16985
rect 430 16850 800 16925
rect 830 16985 1200 16995
rect 830 16925 834 16985
rect 886 16925 1144 16985
rect 1196 16925 1200 16985
rect 830 16850 1200 16925
rect 1230 16985 1600 16995
rect 1230 16925 1234 16985
rect 1286 16925 1544 16985
rect 1596 16925 1600 16985
rect 1230 16850 1600 16925
rect 1630 16985 2000 16995
rect 1630 16925 1634 16985
rect 1686 16925 1944 16985
rect 1996 16925 2000 16985
rect 1630 16850 2000 16925
rect 2030 16985 2400 16995
rect 2030 16925 2034 16985
rect 2086 16925 2344 16985
rect 2396 16925 2400 16985
rect 2030 16850 2400 16925
rect 2430 16985 2800 16995
rect 2430 16925 2434 16985
rect 2486 16925 2744 16985
rect 2796 16925 2800 16985
rect 2430 16850 2800 16925
rect 2830 16985 3200 16995
rect 2830 16925 2834 16985
rect 2886 16925 3144 16985
rect 3196 16925 3200 16985
rect 2830 16850 3200 16925
rect 30 16810 3200 16850
rect 30 16725 400 16810
rect 30 16665 34 16725
rect 86 16665 344 16725
rect 396 16665 400 16725
rect 30 16655 400 16665
rect 430 16725 800 16810
rect 430 16665 434 16725
rect 486 16665 744 16725
rect 796 16665 800 16725
rect 430 16655 800 16665
rect 830 16725 1200 16810
rect 830 16665 834 16725
rect 886 16665 1144 16725
rect 1196 16665 1200 16725
rect 830 16655 1200 16665
rect 1230 16725 1600 16810
rect 1230 16665 1234 16725
rect 1286 16665 1544 16725
rect 1596 16665 1600 16725
rect 1230 16655 1600 16665
rect 1630 16725 2000 16810
rect 1630 16665 1634 16725
rect 1686 16665 1944 16725
rect 1996 16665 2000 16725
rect 1630 16655 2000 16665
rect 2030 16725 2400 16810
rect 2030 16665 2034 16725
rect 2086 16665 2344 16725
rect 2396 16665 2400 16725
rect 2030 16655 2400 16665
rect 2430 16725 2800 16810
rect 2430 16665 2434 16725
rect 2486 16665 2744 16725
rect 2796 16665 2800 16725
rect 2430 16655 2800 16665
rect 2830 16725 3200 16810
rect 2830 16665 2834 16725
rect 2886 16665 3144 16725
rect 3196 16665 3200 16725
rect 2830 16655 3200 16665
rect 3230 16985 3600 16995
rect 3230 16925 3234 16985
rect 3286 16925 3544 16985
rect 3596 16925 3600 16985
rect 3230 16850 3600 16925
rect 3630 16985 4000 16995
rect 3630 16925 3634 16985
rect 3686 16925 3944 16985
rect 3996 16925 4000 16985
rect 3630 16850 4000 16925
rect 4030 16985 4400 16995
rect 4030 16925 4034 16985
rect 4086 16925 4344 16985
rect 4396 16925 4400 16985
rect 4030 16850 4400 16925
rect 4430 16985 4800 16995
rect 4430 16925 4434 16985
rect 4486 16925 4744 16985
rect 4796 16925 4800 16985
rect 4430 16850 4800 16925
rect 4830 16985 5200 16995
rect 4830 16925 4834 16985
rect 4886 16925 5144 16985
rect 5196 16925 5200 16985
rect 4830 16850 5200 16925
rect 5230 16985 5600 16995
rect 5230 16925 5234 16985
rect 5286 16925 5544 16985
rect 5596 16925 5600 16985
rect 5230 16850 5600 16925
rect 5630 16985 6000 16995
rect 5630 16925 5634 16985
rect 5686 16925 5944 16985
rect 5996 16925 6000 16985
rect 5630 16850 6000 16925
rect 3230 16810 6000 16850
rect 3230 16725 3600 16810
rect 3230 16665 3234 16725
rect 3286 16665 3544 16725
rect 3596 16665 3600 16725
rect 3230 16655 3600 16665
rect 3630 16725 4000 16810
rect 3630 16665 3634 16725
rect 3686 16665 3944 16725
rect 3996 16665 4000 16725
rect 3630 16655 4000 16665
rect 4030 16725 4400 16810
rect 4030 16665 4034 16725
rect 4086 16665 4344 16725
rect 4396 16665 4400 16725
rect 4030 16655 4400 16665
rect 4430 16725 4800 16810
rect 4430 16665 4434 16725
rect 4486 16665 4744 16725
rect 4796 16665 4800 16725
rect 4430 16655 4800 16665
rect 4830 16725 5200 16810
rect 4830 16665 4834 16725
rect 4886 16665 5144 16725
rect 5196 16665 5200 16725
rect 4830 16655 5200 16665
rect 5230 16725 5600 16810
rect 5230 16665 5234 16725
rect 5286 16665 5544 16725
rect 5596 16665 5600 16725
rect 5230 16655 5600 16665
rect 5630 16725 6000 16810
rect 5630 16665 5634 16725
rect 5686 16665 5944 16725
rect 5996 16665 6000 16725
rect 5630 16655 6000 16665
rect 6030 16985 6400 16995
rect 6030 16925 6034 16985
rect 6086 16925 6344 16985
rect 6396 16925 6400 16985
rect 6030 16850 6400 16925
rect 6430 16985 6800 16995
rect 6430 16925 6434 16985
rect 6486 16925 6744 16985
rect 6796 16925 6800 16985
rect 6430 16850 6800 16925
rect 6830 16985 7200 16995
rect 6830 16925 6834 16985
rect 6886 16925 7144 16985
rect 7196 16925 7200 16985
rect 6830 16850 7200 16925
rect 7230 16985 7600 16995
rect 7230 16925 7234 16985
rect 7286 16925 7544 16985
rect 7596 16925 7600 16985
rect 7230 16850 7600 16925
rect 7630 16985 8000 16995
rect 7630 16925 7634 16985
rect 7686 16925 7944 16985
rect 7996 16925 8000 16985
rect 7630 16850 8000 16925
rect 8030 16985 8400 16995
rect 8030 16925 8034 16985
rect 8086 16925 8344 16985
rect 8396 16925 8400 16985
rect 8030 16850 8400 16925
rect 8430 16985 8800 16995
rect 8430 16925 8434 16985
rect 8486 16925 8744 16985
rect 8796 16925 8800 16985
rect 8430 16850 8800 16925
rect 8830 16985 9200 16995
rect 8830 16925 8834 16985
rect 8886 16925 9144 16985
rect 9196 16925 9200 16985
rect 8830 16850 9200 16925
rect 9230 16985 9600 16995
rect 9230 16925 9234 16985
rect 9286 16925 9544 16985
rect 9596 16925 9600 16985
rect 9230 16850 9600 16925
rect 9630 16985 10000 16995
rect 9630 16925 9634 16985
rect 9686 16925 9944 16985
rect 9996 16925 10000 16985
rect 9630 16850 10000 16925
rect 10030 16985 10400 16995
rect 10030 16925 10034 16985
rect 10086 16925 10344 16985
rect 10396 16925 10400 16985
rect 10030 16850 10400 16925
rect 10430 16985 10800 16995
rect 10430 16925 10434 16985
rect 10486 16925 10744 16985
rect 10796 16925 10800 16985
rect 10430 16850 10800 16925
rect 10830 16985 11200 16995
rect 10830 16925 10834 16985
rect 10886 16925 11144 16985
rect 11196 16925 11200 16985
rect 10830 16850 11200 16925
rect 11230 16985 11600 16995
rect 11230 16925 11234 16985
rect 11286 16925 11544 16985
rect 11596 16925 11600 16985
rect 11230 16850 11600 16925
rect 11630 16985 12000 16995
rect 11630 16925 11634 16985
rect 11686 16925 11944 16985
rect 11996 16925 12000 16985
rect 11630 16850 12000 16925
rect 12030 16985 12400 16995
rect 12030 16925 12034 16985
rect 12086 16925 12344 16985
rect 12396 16925 12400 16985
rect 12030 16850 12400 16925
rect 12430 16985 12800 16995
rect 12430 16925 12434 16985
rect 12486 16925 12744 16985
rect 12796 16925 12800 16985
rect 12430 16850 12800 16925
rect 12830 16985 13200 16995
rect 12830 16925 12834 16985
rect 12886 16925 13144 16985
rect 13196 16925 13200 16985
rect 12830 16850 13200 16925
rect 6030 16810 13200 16850
rect 6030 16725 6400 16810
rect 6030 16665 6034 16725
rect 6086 16665 6344 16725
rect 6396 16665 6400 16725
rect 6030 16655 6400 16665
rect 6430 16725 6800 16810
rect 6430 16665 6434 16725
rect 6486 16665 6744 16725
rect 6796 16665 6800 16725
rect 6430 16655 6800 16665
rect 6830 16725 7200 16810
rect 6830 16665 6834 16725
rect 6886 16665 7144 16725
rect 7196 16665 7200 16725
rect 6830 16655 7200 16665
rect 7230 16725 7600 16810
rect 7230 16665 7234 16725
rect 7286 16665 7544 16725
rect 7596 16665 7600 16725
rect 7230 16655 7600 16665
rect 7630 16725 8000 16810
rect 7630 16665 7634 16725
rect 7686 16665 7944 16725
rect 7996 16665 8000 16725
rect 7630 16655 8000 16665
rect 8030 16725 8400 16810
rect 8030 16665 8034 16725
rect 8086 16665 8344 16725
rect 8396 16665 8400 16725
rect 8030 16655 8400 16665
rect 8430 16725 8800 16810
rect 8430 16665 8434 16725
rect 8486 16665 8744 16725
rect 8796 16665 8800 16725
rect 8430 16655 8800 16665
rect 8830 16725 9200 16810
rect 8830 16665 8834 16725
rect 8886 16665 9144 16725
rect 9196 16665 9200 16725
rect 8830 16655 9200 16665
rect 9230 16725 9600 16810
rect 9230 16665 9234 16725
rect 9286 16665 9544 16725
rect 9596 16665 9600 16725
rect 9230 16655 9600 16665
rect 9630 16725 10000 16810
rect 9630 16665 9634 16725
rect 9686 16665 9944 16725
rect 9996 16665 10000 16725
rect 9630 16655 10000 16665
rect 10030 16725 10400 16810
rect 10030 16665 10034 16725
rect 10086 16665 10344 16725
rect 10396 16665 10400 16725
rect 10030 16655 10400 16665
rect 10430 16725 10800 16810
rect 10430 16665 10434 16725
rect 10486 16665 10744 16725
rect 10796 16665 10800 16725
rect 10430 16655 10800 16665
rect 10830 16725 11200 16810
rect 10830 16665 10834 16725
rect 10886 16665 11144 16725
rect 11196 16665 11200 16725
rect 10830 16655 11200 16665
rect 11230 16725 11600 16810
rect 11230 16665 11234 16725
rect 11286 16665 11544 16725
rect 11596 16665 11600 16725
rect 11230 16655 11600 16665
rect 11630 16725 12000 16810
rect 11630 16665 11634 16725
rect 11686 16665 11944 16725
rect 11996 16665 12000 16725
rect 11630 16655 12000 16665
rect 12030 16725 12400 16810
rect 12030 16665 12034 16725
rect 12086 16665 12344 16725
rect 12396 16665 12400 16725
rect 12030 16655 12400 16665
rect 12430 16725 12800 16810
rect 12430 16665 12434 16725
rect 12486 16665 12744 16725
rect 12796 16665 12800 16725
rect 12430 16655 12800 16665
rect 12830 16725 13200 16810
rect 12830 16665 12834 16725
rect 12886 16665 13144 16725
rect 13196 16665 13200 16725
rect 12830 16655 13200 16665
rect -330 16625 -324 16655
rect 30 16625 70 16655
rect 430 16625 470 16655
rect 830 16625 870 16655
rect 1230 16625 1270 16655
rect 1630 16625 1670 16655
rect 2030 16625 2070 16655
rect 2430 16625 2470 16655
rect 2830 16625 2870 16655
rect 3230 16625 3270 16655
rect 3630 16625 3670 16655
rect 4030 16625 4070 16655
rect 4430 16625 4470 16655
rect 4830 16625 4870 16655
rect 5230 16625 5270 16655
rect 5630 16625 5670 16655
rect 6030 16625 6070 16655
rect 6430 16625 6470 16655
rect 6830 16625 6870 16655
rect 7230 16625 7270 16655
rect 7630 16625 7670 16655
rect 8030 16625 8070 16655
rect 8430 16625 8470 16655
rect 8830 16625 8870 16655
rect 9230 16625 9270 16655
rect 9630 16625 9670 16655
rect 10030 16625 10070 16655
rect 10430 16625 10470 16655
rect 10830 16625 10870 16655
rect 11230 16625 11270 16655
rect 11630 16625 11670 16655
rect 12030 16625 12070 16655
rect 12430 16625 12470 16655
rect -330 16615 0 16625
rect -314 16555 -56 16615
rect -4 16555 0 16615
rect -330 16355 0 16555
rect -314 16295 -56 16355
rect -4 16295 0 16355
rect -330 16285 0 16295
rect 30 16615 400 16625
rect 30 16555 34 16615
rect 86 16555 344 16615
rect 396 16555 400 16615
rect 30 16480 400 16555
rect 430 16615 800 16625
rect 430 16555 434 16615
rect 486 16555 744 16615
rect 796 16555 800 16615
rect 430 16480 800 16555
rect 830 16615 1200 16625
rect 830 16555 834 16615
rect 886 16555 1144 16615
rect 1196 16555 1200 16615
rect 830 16480 1200 16555
rect 1230 16615 1600 16625
rect 1230 16555 1234 16615
rect 1286 16555 1544 16615
rect 1596 16555 1600 16615
rect 1230 16480 1600 16555
rect 1630 16615 2000 16625
rect 1630 16555 1634 16615
rect 1686 16555 1944 16615
rect 1996 16555 2000 16615
rect 1630 16480 2000 16555
rect 2030 16615 2400 16625
rect 2030 16555 2034 16615
rect 2086 16555 2344 16615
rect 2396 16555 2400 16615
rect 2030 16480 2400 16555
rect 2430 16615 2800 16625
rect 2430 16555 2434 16615
rect 2486 16555 2744 16615
rect 2796 16555 2800 16615
rect 2430 16480 2800 16555
rect 2830 16615 3200 16625
rect 2830 16555 2834 16615
rect 2886 16555 3144 16615
rect 3196 16555 3200 16615
rect 2830 16480 3200 16555
rect 30 16440 3200 16480
rect 30 16355 400 16440
rect 30 16295 34 16355
rect 86 16295 344 16355
rect 396 16295 400 16355
rect 30 16285 400 16295
rect 430 16355 800 16440
rect 430 16295 434 16355
rect 486 16295 744 16355
rect 796 16295 800 16355
rect 430 16285 800 16295
rect 830 16355 1200 16440
rect 830 16295 834 16355
rect 886 16295 1144 16355
rect 1196 16295 1200 16355
rect 830 16285 1200 16295
rect 1230 16355 1600 16440
rect 1230 16295 1234 16355
rect 1286 16295 1544 16355
rect 1596 16295 1600 16355
rect 1230 16285 1600 16295
rect 1630 16355 2000 16440
rect 1630 16295 1634 16355
rect 1686 16295 1944 16355
rect 1996 16295 2000 16355
rect 1630 16285 2000 16295
rect 2030 16355 2400 16440
rect 2030 16295 2034 16355
rect 2086 16295 2344 16355
rect 2396 16295 2400 16355
rect 2030 16285 2400 16295
rect 2430 16355 2800 16440
rect 2430 16295 2434 16355
rect 2486 16295 2744 16355
rect 2796 16295 2800 16355
rect 2430 16285 2800 16295
rect 2830 16355 3200 16440
rect 2830 16295 2834 16355
rect 2886 16295 3144 16355
rect 3196 16295 3200 16355
rect 2830 16285 3200 16295
rect 3230 16615 3600 16625
rect 3230 16555 3234 16615
rect 3286 16555 3544 16615
rect 3596 16555 3600 16615
rect 3230 16480 3600 16555
rect 3630 16615 4000 16625
rect 3630 16555 3634 16615
rect 3686 16555 3944 16615
rect 3996 16555 4000 16615
rect 3630 16480 4000 16555
rect 4030 16615 4400 16625
rect 4030 16555 4034 16615
rect 4086 16555 4344 16615
rect 4396 16555 4400 16615
rect 4030 16480 4400 16555
rect 4430 16615 4800 16625
rect 4430 16555 4434 16615
rect 4486 16555 4744 16615
rect 4796 16555 4800 16615
rect 4430 16480 4800 16555
rect 4830 16615 5200 16625
rect 4830 16555 4834 16615
rect 4886 16555 5144 16615
rect 5196 16555 5200 16615
rect 4830 16480 5200 16555
rect 5230 16615 5600 16625
rect 5230 16555 5234 16615
rect 5286 16555 5544 16615
rect 5596 16555 5600 16615
rect 5230 16480 5600 16555
rect 5630 16615 6000 16625
rect 5630 16555 5634 16615
rect 5686 16555 5944 16615
rect 5996 16555 6000 16615
rect 5630 16480 6000 16555
rect 3230 16440 6000 16480
rect 3230 16355 3600 16440
rect 3230 16295 3234 16355
rect 3286 16295 3544 16355
rect 3596 16295 3600 16355
rect 3230 16285 3600 16295
rect 3630 16355 4000 16440
rect 3630 16295 3634 16355
rect 3686 16295 3944 16355
rect 3996 16295 4000 16355
rect 3630 16285 4000 16295
rect 4030 16355 4400 16440
rect 4030 16295 4034 16355
rect 4086 16295 4344 16355
rect 4396 16295 4400 16355
rect 4030 16285 4400 16295
rect 4430 16355 4800 16440
rect 4430 16295 4434 16355
rect 4486 16295 4744 16355
rect 4796 16295 4800 16355
rect 4430 16285 4800 16295
rect 4830 16355 5200 16440
rect 4830 16295 4834 16355
rect 4886 16295 5144 16355
rect 5196 16295 5200 16355
rect 4830 16285 5200 16295
rect 5230 16355 5600 16440
rect 5230 16295 5234 16355
rect 5286 16295 5544 16355
rect 5596 16295 5600 16355
rect 5230 16285 5600 16295
rect 5630 16355 6000 16440
rect 5630 16295 5634 16355
rect 5686 16295 5944 16355
rect 5996 16295 6000 16355
rect 5630 16285 6000 16295
rect 6030 16615 6400 16625
rect 6030 16555 6034 16615
rect 6086 16555 6344 16615
rect 6396 16555 6400 16615
rect 6030 16480 6400 16555
rect 6430 16615 6800 16625
rect 6430 16555 6434 16615
rect 6486 16555 6744 16615
rect 6796 16555 6800 16615
rect 6430 16480 6800 16555
rect 6830 16615 7200 16625
rect 6830 16555 6834 16615
rect 6886 16555 7144 16615
rect 7196 16555 7200 16615
rect 6830 16480 7200 16555
rect 7230 16615 7600 16625
rect 7230 16555 7234 16615
rect 7286 16555 7544 16615
rect 7596 16555 7600 16615
rect 7230 16480 7600 16555
rect 7630 16615 8000 16625
rect 7630 16555 7634 16615
rect 7686 16555 7944 16615
rect 7996 16555 8000 16615
rect 7630 16480 8000 16555
rect 8030 16615 8400 16625
rect 8030 16555 8034 16615
rect 8086 16555 8344 16615
rect 8396 16555 8400 16615
rect 8030 16480 8400 16555
rect 8430 16615 8800 16625
rect 8430 16555 8434 16615
rect 8486 16555 8744 16615
rect 8796 16555 8800 16615
rect 8430 16480 8800 16555
rect 8830 16615 9200 16625
rect 8830 16555 8834 16615
rect 8886 16555 9144 16615
rect 9196 16555 9200 16615
rect 8830 16480 9200 16555
rect 9230 16615 9600 16625
rect 9230 16555 9234 16615
rect 9286 16555 9544 16615
rect 9596 16555 9600 16615
rect 9230 16480 9600 16555
rect 9630 16615 10000 16625
rect 9630 16555 9634 16615
rect 9686 16555 9944 16615
rect 9996 16555 10000 16615
rect 9630 16480 10000 16555
rect 10030 16615 10400 16625
rect 10030 16555 10034 16615
rect 10086 16555 10344 16615
rect 10396 16555 10400 16615
rect 10030 16480 10400 16555
rect 10430 16615 10800 16625
rect 10430 16555 10434 16615
rect 10486 16555 10744 16615
rect 10796 16555 10800 16615
rect 10430 16480 10800 16555
rect 10830 16615 11200 16625
rect 10830 16555 10834 16615
rect 10886 16555 11144 16615
rect 11196 16555 11200 16615
rect 10830 16480 11200 16555
rect 11230 16615 11600 16625
rect 11230 16555 11234 16615
rect 11286 16555 11544 16615
rect 11596 16555 11600 16615
rect 11230 16480 11600 16555
rect 11630 16615 12000 16625
rect 11630 16555 11634 16615
rect 11686 16555 11944 16615
rect 11996 16555 12000 16615
rect 11630 16480 12000 16555
rect 12030 16615 12400 16625
rect 12030 16555 12034 16615
rect 12086 16555 12344 16615
rect 12396 16555 12400 16615
rect 12030 16480 12400 16555
rect 12430 16615 12800 16625
rect 12430 16555 12434 16615
rect 12486 16555 12744 16615
rect 12796 16555 12800 16615
rect 12430 16480 12800 16555
rect 12830 16615 13200 16625
rect 12830 16555 12834 16615
rect 12886 16555 13144 16615
rect 13196 16555 13200 16615
rect 12830 16480 13200 16555
rect 6030 16440 13200 16480
rect 6030 16355 6400 16440
rect 6030 16295 6034 16355
rect 6086 16295 6344 16355
rect 6396 16295 6400 16355
rect 6030 16285 6400 16295
rect 6430 16355 6800 16440
rect 6430 16295 6434 16355
rect 6486 16295 6744 16355
rect 6796 16295 6800 16355
rect 6430 16285 6800 16295
rect 6830 16355 7200 16440
rect 6830 16295 6834 16355
rect 6886 16295 7144 16355
rect 7196 16295 7200 16355
rect 6830 16285 7200 16295
rect 7230 16355 7600 16440
rect 7230 16295 7234 16355
rect 7286 16295 7544 16355
rect 7596 16295 7600 16355
rect 7230 16285 7600 16295
rect 7630 16355 8000 16440
rect 7630 16295 7634 16355
rect 7686 16295 7944 16355
rect 7996 16295 8000 16355
rect 7630 16285 8000 16295
rect 8030 16355 8400 16440
rect 8030 16295 8034 16355
rect 8086 16295 8344 16355
rect 8396 16295 8400 16355
rect 8030 16285 8400 16295
rect 8430 16355 8800 16440
rect 8430 16295 8434 16355
rect 8486 16295 8744 16355
rect 8796 16295 8800 16355
rect 8430 16285 8800 16295
rect 8830 16355 9200 16440
rect 8830 16295 8834 16355
rect 8886 16295 9144 16355
rect 9196 16295 9200 16355
rect 8830 16285 9200 16295
rect 9230 16355 9600 16440
rect 9230 16295 9234 16355
rect 9286 16295 9544 16355
rect 9596 16295 9600 16355
rect 9230 16285 9600 16295
rect 9630 16355 10000 16440
rect 9630 16295 9634 16355
rect 9686 16295 9944 16355
rect 9996 16295 10000 16355
rect 9630 16285 10000 16295
rect 10030 16355 10400 16440
rect 10030 16295 10034 16355
rect 10086 16295 10344 16355
rect 10396 16295 10400 16355
rect 10030 16285 10400 16295
rect 10430 16355 10800 16440
rect 10430 16295 10434 16355
rect 10486 16295 10744 16355
rect 10796 16295 10800 16355
rect 10430 16285 10800 16295
rect 10830 16355 11200 16440
rect 10830 16295 10834 16355
rect 10886 16295 11144 16355
rect 11196 16295 11200 16355
rect 10830 16285 11200 16295
rect 11230 16355 11600 16440
rect 11230 16295 11234 16355
rect 11286 16295 11544 16355
rect 11596 16295 11600 16355
rect 11230 16285 11600 16295
rect 11630 16355 12000 16440
rect 11630 16295 11634 16355
rect 11686 16295 11944 16355
rect 11996 16295 12000 16355
rect 11630 16285 12000 16295
rect 12030 16355 12400 16440
rect 12030 16295 12034 16355
rect 12086 16295 12344 16355
rect 12396 16295 12400 16355
rect 12030 16285 12400 16295
rect 12430 16355 12800 16440
rect 12430 16295 12434 16355
rect 12486 16295 12744 16355
rect 12796 16295 12800 16355
rect 12430 16285 12800 16295
rect 12830 16355 13200 16440
rect 12830 16295 12834 16355
rect 12886 16295 13144 16355
rect 13196 16295 13200 16355
rect 12830 16285 13200 16295
rect -330 16255 -324 16285
rect 30 16255 70 16285
rect 430 16255 470 16285
rect 830 16255 870 16285
rect 1230 16255 1270 16285
rect 1630 16255 1670 16285
rect 2030 16255 2070 16285
rect 2430 16255 2470 16285
rect 2830 16255 2870 16285
rect 3230 16255 3270 16285
rect 3630 16255 3670 16285
rect 4030 16255 4070 16285
rect 4430 16255 4470 16285
rect 4830 16255 4870 16285
rect 5230 16255 5270 16285
rect 5630 16255 5670 16285
rect 6030 16255 6070 16285
rect 6430 16255 6470 16285
rect 6830 16255 6870 16285
rect 7230 16255 7270 16285
rect 7630 16255 7670 16285
rect 8030 16255 8070 16285
rect 8430 16255 8470 16285
rect 8830 16255 8870 16285
rect 9230 16255 9270 16285
rect 9630 16255 9670 16285
rect 10030 16255 10070 16285
rect 10430 16255 10470 16285
rect 10830 16255 10870 16285
rect 11230 16255 11270 16285
rect 11630 16255 11670 16285
rect 12030 16255 12070 16285
rect 12430 16255 12470 16285
rect -330 16245 0 16255
rect -314 16185 -56 16245
rect -4 16185 0 16245
rect -330 15985 0 16185
rect -314 15925 -56 15985
rect -4 15925 0 15985
rect -330 15915 0 15925
rect 30 16245 400 16255
rect 30 16185 34 16245
rect 86 16185 344 16245
rect 396 16185 400 16245
rect 30 16110 400 16185
rect 430 16245 800 16255
rect 430 16185 434 16245
rect 486 16185 744 16245
rect 796 16185 800 16245
rect 430 16110 800 16185
rect 830 16245 1200 16255
rect 830 16185 834 16245
rect 886 16185 1144 16245
rect 1196 16185 1200 16245
rect 830 16110 1200 16185
rect 1230 16245 1600 16255
rect 1230 16185 1234 16245
rect 1286 16185 1544 16245
rect 1596 16185 1600 16245
rect 1230 16110 1600 16185
rect 1630 16245 2000 16255
rect 1630 16185 1634 16245
rect 1686 16185 1944 16245
rect 1996 16185 2000 16245
rect 1630 16110 2000 16185
rect 2030 16245 2400 16255
rect 2030 16185 2034 16245
rect 2086 16185 2344 16245
rect 2396 16185 2400 16245
rect 2030 16110 2400 16185
rect 2430 16245 2800 16255
rect 2430 16185 2434 16245
rect 2486 16185 2744 16245
rect 2796 16185 2800 16245
rect 2430 16110 2800 16185
rect 2830 16245 3200 16255
rect 2830 16185 2834 16245
rect 2886 16185 3144 16245
rect 3196 16185 3200 16245
rect 2830 16110 3200 16185
rect 30 16070 3200 16110
rect 30 15985 400 16070
rect 30 15925 34 15985
rect 86 15925 344 15985
rect 396 15925 400 15985
rect 30 15915 400 15925
rect 430 15985 800 16070
rect 430 15925 434 15985
rect 486 15925 744 15985
rect 796 15925 800 15985
rect 430 15915 800 15925
rect 830 15985 1200 16070
rect 830 15925 834 15985
rect 886 15925 1144 15985
rect 1196 15925 1200 15985
rect 830 15915 1200 15925
rect 1230 15985 1600 16070
rect 1230 15925 1234 15985
rect 1286 15925 1544 15985
rect 1596 15925 1600 15985
rect 1230 15915 1600 15925
rect 1630 15985 2000 16070
rect 1630 15925 1634 15985
rect 1686 15925 1944 15985
rect 1996 15925 2000 15985
rect 1630 15915 2000 15925
rect 2030 15985 2400 16070
rect 2030 15925 2034 15985
rect 2086 15925 2344 15985
rect 2396 15925 2400 15985
rect 2030 15915 2400 15925
rect 2430 15985 2800 16070
rect 2430 15925 2434 15985
rect 2486 15925 2744 15985
rect 2796 15925 2800 15985
rect 2430 15915 2800 15925
rect 2830 15985 3200 16070
rect 2830 15925 2834 15985
rect 2886 15925 3144 15985
rect 3196 15925 3200 15985
rect 2830 15915 3200 15925
rect 3230 16245 3600 16255
rect 3230 16185 3234 16245
rect 3286 16185 3544 16245
rect 3596 16185 3600 16245
rect 3230 16110 3600 16185
rect 3630 16245 4000 16255
rect 3630 16185 3634 16245
rect 3686 16185 3944 16245
rect 3996 16185 4000 16245
rect 3630 16110 4000 16185
rect 4030 16245 4400 16255
rect 4030 16185 4034 16245
rect 4086 16185 4344 16245
rect 4396 16185 4400 16245
rect 4030 16110 4400 16185
rect 4430 16245 4800 16255
rect 4430 16185 4434 16245
rect 4486 16185 4744 16245
rect 4796 16185 4800 16245
rect 4430 16110 4800 16185
rect 4830 16245 5200 16255
rect 4830 16185 4834 16245
rect 4886 16185 5144 16245
rect 5196 16185 5200 16245
rect 4830 16110 5200 16185
rect 5230 16245 5600 16255
rect 5230 16185 5234 16245
rect 5286 16185 5544 16245
rect 5596 16185 5600 16245
rect 5230 16110 5600 16185
rect 5630 16245 6000 16255
rect 5630 16185 5634 16245
rect 5686 16185 5944 16245
rect 5996 16185 6000 16245
rect 5630 16110 6000 16185
rect 3230 16070 6000 16110
rect 3230 15985 3600 16070
rect 3230 15925 3234 15985
rect 3286 15925 3544 15985
rect 3596 15925 3600 15985
rect 3230 15915 3600 15925
rect 3630 15985 4000 16070
rect 3630 15925 3634 15985
rect 3686 15925 3944 15985
rect 3996 15925 4000 15985
rect 3630 15915 4000 15925
rect 4030 15985 4400 16070
rect 4030 15925 4034 15985
rect 4086 15925 4344 15985
rect 4396 15925 4400 15985
rect 4030 15915 4400 15925
rect 4430 15985 4800 16070
rect 4430 15925 4434 15985
rect 4486 15925 4744 15985
rect 4796 15925 4800 15985
rect 4430 15915 4800 15925
rect 4830 15985 5200 16070
rect 4830 15925 4834 15985
rect 4886 15925 5144 15985
rect 5196 15925 5200 15985
rect 4830 15915 5200 15925
rect 5230 15985 5600 16070
rect 5230 15925 5234 15985
rect 5286 15925 5544 15985
rect 5596 15925 5600 15985
rect 5230 15915 5600 15925
rect 5630 15985 6000 16070
rect 5630 15925 5634 15985
rect 5686 15925 5944 15985
rect 5996 15925 6000 15985
rect 5630 15915 6000 15925
rect 6030 16245 6400 16255
rect 6030 16185 6034 16245
rect 6086 16185 6344 16245
rect 6396 16185 6400 16245
rect 6030 16110 6400 16185
rect 6430 16245 6800 16255
rect 6430 16185 6434 16245
rect 6486 16185 6744 16245
rect 6796 16185 6800 16245
rect 6430 16110 6800 16185
rect 6830 16245 7200 16255
rect 6830 16185 6834 16245
rect 6886 16185 7144 16245
rect 7196 16185 7200 16245
rect 6830 16110 7200 16185
rect 7230 16245 7600 16255
rect 7230 16185 7234 16245
rect 7286 16185 7544 16245
rect 7596 16185 7600 16245
rect 7230 16110 7600 16185
rect 7630 16245 8000 16255
rect 7630 16185 7634 16245
rect 7686 16185 7944 16245
rect 7996 16185 8000 16245
rect 7630 16110 8000 16185
rect 8030 16245 8400 16255
rect 8030 16185 8034 16245
rect 8086 16185 8344 16245
rect 8396 16185 8400 16245
rect 8030 16110 8400 16185
rect 8430 16245 8800 16255
rect 8430 16185 8434 16245
rect 8486 16185 8744 16245
rect 8796 16185 8800 16245
rect 8430 16110 8800 16185
rect 8830 16245 9200 16255
rect 8830 16185 8834 16245
rect 8886 16185 9144 16245
rect 9196 16185 9200 16245
rect 8830 16110 9200 16185
rect 9230 16245 9600 16255
rect 9230 16185 9234 16245
rect 9286 16185 9544 16245
rect 9596 16185 9600 16245
rect 9230 16110 9600 16185
rect 9630 16245 10000 16255
rect 9630 16185 9634 16245
rect 9686 16185 9944 16245
rect 9996 16185 10000 16245
rect 9630 16110 10000 16185
rect 10030 16245 10400 16255
rect 10030 16185 10034 16245
rect 10086 16185 10344 16245
rect 10396 16185 10400 16245
rect 10030 16110 10400 16185
rect 10430 16245 10800 16255
rect 10430 16185 10434 16245
rect 10486 16185 10744 16245
rect 10796 16185 10800 16245
rect 10430 16110 10800 16185
rect 10830 16245 11200 16255
rect 10830 16185 10834 16245
rect 10886 16185 11144 16245
rect 11196 16185 11200 16245
rect 10830 16110 11200 16185
rect 11230 16245 11600 16255
rect 11230 16185 11234 16245
rect 11286 16185 11544 16245
rect 11596 16185 11600 16245
rect 11230 16110 11600 16185
rect 11630 16245 12000 16255
rect 11630 16185 11634 16245
rect 11686 16185 11944 16245
rect 11996 16185 12000 16245
rect 11630 16110 12000 16185
rect 12030 16245 12400 16255
rect 12030 16185 12034 16245
rect 12086 16185 12344 16245
rect 12396 16185 12400 16245
rect 12030 16110 12400 16185
rect 12430 16245 12800 16255
rect 12430 16185 12434 16245
rect 12486 16185 12744 16245
rect 12796 16185 12800 16245
rect 12430 16110 12800 16185
rect 12830 16245 13200 16255
rect 12830 16185 12834 16245
rect 12886 16185 13144 16245
rect 13196 16185 13200 16245
rect 12830 16110 13200 16185
rect 6030 16070 13200 16110
rect 6030 15985 6400 16070
rect 6030 15925 6034 15985
rect 6086 15925 6344 15985
rect 6396 15925 6400 15985
rect 6030 15915 6400 15925
rect 6430 15985 6800 16070
rect 6430 15925 6434 15985
rect 6486 15925 6744 15985
rect 6796 15925 6800 15985
rect 6430 15915 6800 15925
rect 6830 15985 7200 16070
rect 6830 15925 6834 15985
rect 6886 15925 7144 15985
rect 7196 15925 7200 15985
rect 6830 15915 7200 15925
rect 7230 15985 7600 16070
rect 7230 15925 7234 15985
rect 7286 15925 7544 15985
rect 7596 15925 7600 15985
rect 7230 15915 7600 15925
rect 7630 15985 8000 16070
rect 7630 15925 7634 15985
rect 7686 15925 7944 15985
rect 7996 15925 8000 15985
rect 7630 15915 8000 15925
rect 8030 15985 8400 16070
rect 8030 15925 8034 15985
rect 8086 15925 8344 15985
rect 8396 15925 8400 15985
rect 8030 15915 8400 15925
rect 8430 15985 8800 16070
rect 8430 15925 8434 15985
rect 8486 15925 8744 15985
rect 8796 15925 8800 15985
rect 8430 15915 8800 15925
rect 8830 15985 9200 16070
rect 8830 15925 8834 15985
rect 8886 15925 9144 15985
rect 9196 15925 9200 15985
rect 8830 15915 9200 15925
rect 9230 15985 9600 16070
rect 9230 15925 9234 15985
rect 9286 15925 9544 15985
rect 9596 15925 9600 15985
rect 9230 15915 9600 15925
rect 9630 15985 10000 16070
rect 9630 15925 9634 15985
rect 9686 15925 9944 15985
rect 9996 15925 10000 15985
rect 9630 15915 10000 15925
rect 10030 15985 10400 16070
rect 10030 15925 10034 15985
rect 10086 15925 10344 15985
rect 10396 15925 10400 15985
rect 10030 15915 10400 15925
rect 10430 15985 10800 16070
rect 10430 15925 10434 15985
rect 10486 15925 10744 15985
rect 10796 15925 10800 15985
rect 10430 15915 10800 15925
rect 10830 15985 11200 16070
rect 10830 15925 10834 15985
rect 10886 15925 11144 15985
rect 11196 15925 11200 15985
rect 10830 15915 11200 15925
rect 11230 15985 11600 16070
rect 11230 15925 11234 15985
rect 11286 15925 11544 15985
rect 11596 15925 11600 15985
rect 11230 15915 11600 15925
rect 11630 15985 12000 16070
rect 11630 15925 11634 15985
rect 11686 15925 11944 15985
rect 11996 15925 12000 15985
rect 11630 15915 12000 15925
rect 12030 15985 12400 16070
rect 12030 15925 12034 15985
rect 12086 15925 12344 15985
rect 12396 15925 12400 15985
rect 12030 15915 12400 15925
rect 12430 15985 12800 16070
rect 12430 15925 12434 15985
rect 12486 15925 12744 15985
rect 12796 15925 12800 15985
rect 12430 15915 12800 15925
rect 12830 15985 13200 16070
rect 12830 15925 12834 15985
rect 12886 15925 13144 15985
rect 13196 15925 13200 15985
rect 12830 15915 13200 15925
rect -330 15885 -324 15915
rect 30 15885 70 15915
rect 430 15885 470 15915
rect 830 15885 870 15915
rect 1230 15885 1270 15915
rect 1630 15885 1670 15915
rect 2030 15885 2070 15915
rect 2430 15885 2470 15915
rect 2830 15885 2870 15915
rect 3230 15885 3270 15915
rect 3630 15885 3670 15915
rect 4030 15885 4070 15915
rect 4430 15885 4470 15915
rect 4830 15885 4870 15915
rect 5230 15885 5270 15915
rect 5630 15885 5670 15915
rect 6030 15885 6070 15915
rect 6430 15885 6470 15915
rect 6830 15885 6870 15915
rect 7230 15885 7270 15915
rect 7630 15885 7670 15915
rect 8030 15885 8070 15915
rect 8430 15885 8470 15915
rect 8830 15885 8870 15915
rect 9230 15885 9270 15915
rect 9630 15885 9670 15915
rect 10030 15885 10070 15915
rect 10430 15885 10470 15915
rect 10830 15885 10870 15915
rect 11230 15885 11270 15915
rect 11630 15885 11670 15915
rect 12030 15885 12070 15915
rect 12430 15885 12470 15915
rect -330 15875 0 15885
rect -314 15815 -56 15875
rect -4 15815 0 15875
rect -330 15615 0 15815
rect -314 15555 -56 15615
rect -4 15555 0 15615
rect -330 15545 0 15555
rect 30 15875 400 15885
rect 30 15815 34 15875
rect 86 15815 344 15875
rect 396 15815 400 15875
rect 30 15740 400 15815
rect 430 15875 800 15885
rect 430 15815 434 15875
rect 486 15815 744 15875
rect 796 15815 800 15875
rect 430 15740 800 15815
rect 830 15875 1200 15885
rect 830 15815 834 15875
rect 886 15815 1144 15875
rect 1196 15815 1200 15875
rect 830 15740 1200 15815
rect 1230 15875 1600 15885
rect 1230 15815 1234 15875
rect 1286 15815 1544 15875
rect 1596 15815 1600 15875
rect 1230 15740 1600 15815
rect 1630 15875 2000 15885
rect 1630 15815 1634 15875
rect 1686 15815 1944 15875
rect 1996 15815 2000 15875
rect 1630 15740 2000 15815
rect 2030 15875 2400 15885
rect 2030 15815 2034 15875
rect 2086 15815 2344 15875
rect 2396 15815 2400 15875
rect 2030 15740 2400 15815
rect 2430 15875 2800 15885
rect 2430 15815 2434 15875
rect 2486 15815 2744 15875
rect 2796 15815 2800 15875
rect 2430 15740 2800 15815
rect 2830 15875 3200 15885
rect 2830 15815 2834 15875
rect 2886 15815 3144 15875
rect 3196 15815 3200 15875
rect 2830 15740 3200 15815
rect 30 15700 3200 15740
rect 30 15615 400 15700
rect 30 15555 34 15615
rect 86 15555 344 15615
rect 396 15555 400 15615
rect 30 15545 400 15555
rect 430 15615 800 15700
rect 430 15555 434 15615
rect 486 15555 744 15615
rect 796 15555 800 15615
rect 430 15545 800 15555
rect 830 15615 1200 15700
rect 830 15555 834 15615
rect 886 15555 1144 15615
rect 1196 15555 1200 15615
rect 830 15545 1200 15555
rect 1230 15615 1600 15700
rect 1230 15555 1234 15615
rect 1286 15555 1544 15615
rect 1596 15555 1600 15615
rect 1230 15545 1600 15555
rect 1630 15615 2000 15700
rect 1630 15555 1634 15615
rect 1686 15555 1944 15615
rect 1996 15555 2000 15615
rect 1630 15545 2000 15555
rect 2030 15615 2400 15700
rect 2030 15555 2034 15615
rect 2086 15555 2344 15615
rect 2396 15555 2400 15615
rect 2030 15545 2400 15555
rect 2430 15615 2800 15700
rect 2430 15555 2434 15615
rect 2486 15555 2744 15615
rect 2796 15555 2800 15615
rect 2430 15545 2800 15555
rect 2830 15615 3200 15700
rect 2830 15555 2834 15615
rect 2886 15555 3144 15615
rect 3196 15555 3200 15615
rect 2830 15545 3200 15555
rect 3230 15875 3600 15885
rect 3230 15815 3234 15875
rect 3286 15815 3544 15875
rect 3596 15815 3600 15875
rect 3230 15740 3600 15815
rect 3630 15875 4000 15885
rect 3630 15815 3634 15875
rect 3686 15815 3944 15875
rect 3996 15815 4000 15875
rect 3630 15740 4000 15815
rect 4030 15875 4400 15885
rect 4030 15815 4034 15875
rect 4086 15815 4344 15875
rect 4396 15815 4400 15875
rect 4030 15740 4400 15815
rect 4430 15875 4800 15885
rect 4430 15815 4434 15875
rect 4486 15815 4744 15875
rect 4796 15815 4800 15875
rect 4430 15740 4800 15815
rect 4830 15875 5200 15885
rect 4830 15815 4834 15875
rect 4886 15815 5144 15875
rect 5196 15815 5200 15875
rect 4830 15740 5200 15815
rect 5230 15875 5600 15885
rect 5230 15815 5234 15875
rect 5286 15815 5544 15875
rect 5596 15815 5600 15875
rect 5230 15740 5600 15815
rect 5630 15875 6000 15885
rect 5630 15815 5634 15875
rect 5686 15815 5944 15875
rect 5996 15815 6000 15875
rect 5630 15740 6000 15815
rect 3230 15700 6000 15740
rect 3230 15615 3600 15700
rect 3230 15555 3234 15615
rect 3286 15555 3544 15615
rect 3596 15555 3600 15615
rect 3230 15545 3600 15555
rect 3630 15615 4000 15700
rect 3630 15555 3634 15615
rect 3686 15555 3944 15615
rect 3996 15555 4000 15615
rect 3630 15545 4000 15555
rect 4030 15615 4400 15700
rect 4030 15555 4034 15615
rect 4086 15555 4344 15615
rect 4396 15555 4400 15615
rect 4030 15545 4400 15555
rect 4430 15615 4800 15700
rect 4430 15555 4434 15615
rect 4486 15555 4744 15615
rect 4796 15555 4800 15615
rect 4430 15545 4800 15555
rect 4830 15615 5200 15700
rect 4830 15555 4834 15615
rect 4886 15555 5144 15615
rect 5196 15555 5200 15615
rect 4830 15545 5200 15555
rect 5230 15615 5600 15700
rect 5230 15555 5234 15615
rect 5286 15555 5544 15615
rect 5596 15555 5600 15615
rect 5230 15545 5600 15555
rect 5630 15615 6000 15700
rect 5630 15555 5634 15615
rect 5686 15555 5944 15615
rect 5996 15555 6000 15615
rect 5630 15545 6000 15555
rect 6030 15875 6400 15885
rect 6030 15815 6034 15875
rect 6086 15815 6344 15875
rect 6396 15815 6400 15875
rect 6030 15740 6400 15815
rect 6430 15875 6800 15885
rect 6430 15815 6434 15875
rect 6486 15815 6744 15875
rect 6796 15815 6800 15875
rect 6430 15740 6800 15815
rect 6830 15875 7200 15885
rect 6830 15815 6834 15875
rect 6886 15815 7144 15875
rect 7196 15815 7200 15875
rect 6830 15740 7200 15815
rect 7230 15875 7600 15885
rect 7230 15815 7234 15875
rect 7286 15815 7544 15875
rect 7596 15815 7600 15875
rect 7230 15740 7600 15815
rect 7630 15875 8000 15885
rect 7630 15815 7634 15875
rect 7686 15815 7944 15875
rect 7996 15815 8000 15875
rect 7630 15740 8000 15815
rect 8030 15875 8400 15885
rect 8030 15815 8034 15875
rect 8086 15815 8344 15875
rect 8396 15815 8400 15875
rect 8030 15740 8400 15815
rect 8430 15875 8800 15885
rect 8430 15815 8434 15875
rect 8486 15815 8744 15875
rect 8796 15815 8800 15875
rect 8430 15740 8800 15815
rect 8830 15875 9200 15885
rect 8830 15815 8834 15875
rect 8886 15815 9144 15875
rect 9196 15815 9200 15875
rect 8830 15740 9200 15815
rect 9230 15875 9600 15885
rect 9230 15815 9234 15875
rect 9286 15815 9544 15875
rect 9596 15815 9600 15875
rect 9230 15740 9600 15815
rect 9630 15875 10000 15885
rect 9630 15815 9634 15875
rect 9686 15815 9944 15875
rect 9996 15815 10000 15875
rect 9630 15740 10000 15815
rect 10030 15875 10400 15885
rect 10030 15815 10034 15875
rect 10086 15815 10344 15875
rect 10396 15815 10400 15875
rect 10030 15740 10400 15815
rect 10430 15875 10800 15885
rect 10430 15815 10434 15875
rect 10486 15815 10744 15875
rect 10796 15815 10800 15875
rect 10430 15740 10800 15815
rect 10830 15875 11200 15885
rect 10830 15815 10834 15875
rect 10886 15815 11144 15875
rect 11196 15815 11200 15875
rect 10830 15740 11200 15815
rect 11230 15875 11600 15885
rect 11230 15815 11234 15875
rect 11286 15815 11544 15875
rect 11596 15815 11600 15875
rect 11230 15740 11600 15815
rect 11630 15875 12000 15885
rect 11630 15815 11634 15875
rect 11686 15815 11944 15875
rect 11996 15815 12000 15875
rect 11630 15740 12000 15815
rect 12030 15875 12400 15885
rect 12030 15815 12034 15875
rect 12086 15815 12344 15875
rect 12396 15815 12400 15875
rect 12030 15740 12400 15815
rect 12430 15875 12800 15885
rect 12430 15815 12434 15875
rect 12486 15815 12744 15875
rect 12796 15815 12800 15875
rect 12430 15740 12800 15815
rect 12830 15875 13200 15885
rect 12830 15815 12834 15875
rect 12886 15815 13144 15875
rect 13196 15815 13200 15875
rect 12830 15740 13200 15815
rect 6030 15700 13200 15740
rect 6030 15615 6400 15700
rect 6030 15555 6034 15615
rect 6086 15555 6344 15615
rect 6396 15555 6400 15615
rect 6030 15545 6400 15555
rect 6430 15615 6800 15700
rect 6430 15555 6434 15615
rect 6486 15555 6744 15615
rect 6796 15555 6800 15615
rect 6430 15545 6800 15555
rect 6830 15615 7200 15700
rect 6830 15555 6834 15615
rect 6886 15555 7144 15615
rect 7196 15555 7200 15615
rect 6830 15545 7200 15555
rect 7230 15615 7600 15700
rect 7230 15555 7234 15615
rect 7286 15555 7544 15615
rect 7596 15555 7600 15615
rect 7230 15545 7600 15555
rect 7630 15615 8000 15700
rect 7630 15555 7634 15615
rect 7686 15555 7944 15615
rect 7996 15555 8000 15615
rect 7630 15545 8000 15555
rect 8030 15615 8400 15700
rect 8030 15555 8034 15615
rect 8086 15555 8344 15615
rect 8396 15555 8400 15615
rect 8030 15545 8400 15555
rect 8430 15615 8800 15700
rect 8430 15555 8434 15615
rect 8486 15555 8744 15615
rect 8796 15555 8800 15615
rect 8430 15545 8800 15555
rect 8830 15615 9200 15700
rect 8830 15555 8834 15615
rect 8886 15555 9144 15615
rect 9196 15555 9200 15615
rect 8830 15545 9200 15555
rect 9230 15615 9600 15700
rect 9230 15555 9234 15615
rect 9286 15555 9544 15615
rect 9596 15555 9600 15615
rect 9230 15545 9600 15555
rect 9630 15615 10000 15700
rect 9630 15555 9634 15615
rect 9686 15555 9944 15615
rect 9996 15555 10000 15615
rect 9630 15545 10000 15555
rect 10030 15615 10400 15700
rect 10030 15555 10034 15615
rect 10086 15555 10344 15615
rect 10396 15555 10400 15615
rect 10030 15545 10400 15555
rect 10430 15615 10800 15700
rect 10430 15555 10434 15615
rect 10486 15555 10744 15615
rect 10796 15555 10800 15615
rect 10430 15545 10800 15555
rect 10830 15615 11200 15700
rect 10830 15555 10834 15615
rect 10886 15555 11144 15615
rect 11196 15555 11200 15615
rect 10830 15545 11200 15555
rect 11230 15615 11600 15700
rect 11230 15555 11234 15615
rect 11286 15555 11544 15615
rect 11596 15555 11600 15615
rect 11230 15545 11600 15555
rect 11630 15615 12000 15700
rect 11630 15555 11634 15615
rect 11686 15555 11944 15615
rect 11996 15555 12000 15615
rect 11630 15545 12000 15555
rect 12030 15615 12400 15700
rect 12030 15555 12034 15615
rect 12086 15555 12344 15615
rect 12396 15555 12400 15615
rect 12030 15545 12400 15555
rect 12430 15615 12800 15700
rect 12430 15555 12434 15615
rect 12486 15555 12744 15615
rect 12796 15555 12800 15615
rect 12430 15545 12800 15555
rect 12830 15615 13200 15700
rect 12830 15555 12834 15615
rect 12886 15555 13144 15615
rect 13196 15555 13200 15615
rect 12830 15545 13200 15555
rect -330 15515 -324 15545
rect 30 15515 70 15545
rect 430 15515 470 15545
rect 830 15515 870 15545
rect 1230 15515 1270 15545
rect 1630 15515 1670 15545
rect 2030 15515 2070 15545
rect 2430 15515 2470 15545
rect 2830 15515 2870 15545
rect 3230 15515 3270 15545
rect 3630 15515 3670 15545
rect 4030 15515 4070 15545
rect 4430 15515 4470 15545
rect 4830 15515 4870 15545
rect 5230 15515 5270 15545
rect 5630 15515 5670 15545
rect 6030 15515 6070 15545
rect 6430 15515 6470 15545
rect 6830 15515 6870 15545
rect 7230 15515 7270 15545
rect 7630 15515 7670 15545
rect -330 15505 0 15515
rect -314 15445 -56 15505
rect -4 15445 0 15505
rect -330 15245 0 15445
rect -314 15185 -56 15245
rect -4 15185 0 15245
rect -330 15175 0 15185
rect 30 15505 400 15515
rect 30 15445 34 15505
rect 86 15445 344 15505
rect 396 15445 400 15505
rect 30 15370 400 15445
rect 430 15505 800 15515
rect 430 15445 434 15505
rect 486 15445 744 15505
rect 796 15445 800 15505
rect 430 15370 800 15445
rect 830 15505 1200 15515
rect 830 15445 834 15505
rect 886 15445 1144 15505
rect 1196 15445 1200 15505
rect 830 15370 1200 15445
rect 1230 15505 1600 15515
rect 1230 15445 1234 15505
rect 1286 15445 1544 15505
rect 1596 15445 1600 15505
rect 1230 15370 1600 15445
rect 1630 15505 2000 15515
rect 1630 15445 1634 15505
rect 1686 15445 1944 15505
rect 1996 15445 2000 15505
rect 1630 15370 2000 15445
rect 2030 15505 2400 15515
rect 2030 15445 2034 15505
rect 2086 15445 2344 15505
rect 2396 15445 2400 15505
rect 2030 15370 2400 15445
rect 2430 15505 2800 15515
rect 2430 15445 2434 15505
rect 2486 15445 2744 15505
rect 2796 15445 2800 15505
rect 2430 15370 2800 15445
rect 2830 15505 3200 15515
rect 2830 15445 2834 15505
rect 2886 15445 3144 15505
rect 3196 15445 3200 15505
rect 2830 15370 3200 15445
rect 30 15330 3200 15370
rect 30 15245 400 15330
rect 30 15185 34 15245
rect 86 15185 344 15245
rect 396 15185 400 15245
rect 30 15175 400 15185
rect 430 15245 800 15330
rect 430 15185 434 15245
rect 486 15185 744 15245
rect 796 15185 800 15245
rect 430 15175 800 15185
rect 830 15245 1200 15330
rect 830 15185 834 15245
rect 886 15185 1144 15245
rect 1196 15185 1200 15245
rect 830 15175 1200 15185
rect 1230 15245 1600 15330
rect 1230 15185 1234 15245
rect 1286 15185 1544 15245
rect 1596 15185 1600 15245
rect 1230 15175 1600 15185
rect 1630 15245 2000 15330
rect 1630 15185 1634 15245
rect 1686 15185 1944 15245
rect 1996 15185 2000 15245
rect 1630 15175 2000 15185
rect 2030 15245 2400 15330
rect 2030 15185 2034 15245
rect 2086 15185 2344 15245
rect 2396 15185 2400 15245
rect 2030 15175 2400 15185
rect 2430 15245 2800 15330
rect 2430 15185 2434 15245
rect 2486 15185 2744 15245
rect 2796 15185 2800 15245
rect 2430 15175 2800 15185
rect 2830 15245 3200 15330
rect 2830 15185 2834 15245
rect 2886 15185 3144 15245
rect 3196 15185 3200 15245
rect 2830 15175 3200 15185
rect 3230 15505 3600 15515
rect 3230 15445 3234 15505
rect 3286 15445 3544 15505
rect 3596 15445 3600 15505
rect 3230 15370 3600 15445
rect 3630 15505 4000 15515
rect 3630 15445 3634 15505
rect 3686 15445 3944 15505
rect 3996 15445 4000 15505
rect 3630 15370 4000 15445
rect 4030 15505 4400 15515
rect 4030 15445 4034 15505
rect 4086 15445 4344 15505
rect 4396 15445 4400 15505
rect 4030 15370 4400 15445
rect 4430 15505 4800 15515
rect 4430 15445 4434 15505
rect 4486 15445 4744 15505
rect 4796 15445 4800 15505
rect 4430 15370 4800 15445
rect 4830 15505 5200 15515
rect 4830 15445 4834 15505
rect 4886 15445 5144 15505
rect 5196 15445 5200 15505
rect 4830 15370 5200 15445
rect 5230 15505 5600 15515
rect 5230 15445 5234 15505
rect 5286 15445 5544 15505
rect 5596 15445 5600 15505
rect 5230 15370 5600 15445
rect 5630 15505 6000 15515
rect 5630 15445 5634 15505
rect 5686 15445 5944 15505
rect 5996 15445 6000 15505
rect 5630 15370 6000 15445
rect 3230 15330 6000 15370
rect 3230 15245 3600 15330
rect 3230 15185 3234 15245
rect 3286 15185 3544 15245
rect 3596 15185 3600 15245
rect 3230 15175 3600 15185
rect 3630 15245 4000 15330
rect 3630 15185 3634 15245
rect 3686 15185 3944 15245
rect 3996 15185 4000 15245
rect 3630 15175 4000 15185
rect 4030 15245 4400 15330
rect 4030 15185 4034 15245
rect 4086 15185 4344 15245
rect 4396 15185 4400 15245
rect 4030 15175 4400 15185
rect 4430 15245 4800 15330
rect 4430 15185 4434 15245
rect 4486 15185 4744 15245
rect 4796 15185 4800 15245
rect 4430 15175 4800 15185
rect 4830 15245 5200 15330
rect 4830 15185 4834 15245
rect 4886 15185 5144 15245
rect 5196 15185 5200 15245
rect 4830 15175 5200 15185
rect 5230 15245 5600 15330
rect 5230 15185 5234 15245
rect 5286 15185 5544 15245
rect 5596 15185 5600 15245
rect 5230 15175 5600 15185
rect 5630 15245 6000 15330
rect 5630 15185 5634 15245
rect 5686 15185 5944 15245
rect 5996 15185 6000 15245
rect 5630 15175 6000 15185
rect 6030 15505 6400 15515
rect 6030 15445 6034 15505
rect 6086 15445 6344 15505
rect 6396 15445 6400 15505
rect 6030 15370 6400 15445
rect 6430 15505 6800 15515
rect 6430 15445 6434 15505
rect 6486 15445 6744 15505
rect 6796 15445 6800 15505
rect 6430 15370 6800 15445
rect 6830 15505 7200 15515
rect 6830 15445 6834 15505
rect 6886 15445 7144 15505
rect 7196 15445 7200 15505
rect 6830 15370 7200 15445
rect 7230 15505 7600 15515
rect 7230 15445 7234 15505
rect 7286 15445 7544 15505
rect 7596 15445 7600 15505
rect 7230 15370 7600 15445
rect 7630 15505 8000 15515
rect 7630 15445 7634 15505
rect 7686 15445 7944 15505
rect 7996 15445 8000 15505
rect 7630 15370 8000 15445
rect 6030 15330 8000 15370
rect 6030 15245 6400 15330
rect 6030 15185 6034 15245
rect 6086 15185 6344 15245
rect 6396 15185 6400 15245
rect 6030 15175 6400 15185
rect 6430 15245 6800 15330
rect 6430 15185 6434 15245
rect 6486 15185 6744 15245
rect 6796 15185 6800 15245
rect 6430 15175 6800 15185
rect 6830 15245 7200 15330
rect 6830 15185 6834 15245
rect 6886 15185 7144 15245
rect 7196 15185 7200 15245
rect 6830 15175 7200 15185
rect 7230 15245 7600 15330
rect 7230 15185 7234 15245
rect 7286 15185 7544 15245
rect 7596 15185 7600 15245
rect 7230 15175 7600 15185
rect 7630 15245 8000 15330
rect 7630 15185 7634 15245
rect 7686 15185 7944 15245
rect 7996 15185 8000 15245
rect 7630 15175 8000 15185
rect 8030 15505 8400 15515
rect 8030 15445 8034 15505
rect 8086 15445 8344 15505
rect 8396 15445 8400 15505
rect 8030 15370 8400 15445
rect 8430 15505 8800 15515
rect 8430 15445 8434 15505
rect 8486 15445 8744 15505
rect 8796 15445 8800 15505
rect 8430 15370 8800 15445
rect 8830 15505 9200 15515
rect 8830 15445 8834 15505
rect 8886 15445 9144 15505
rect 9196 15445 9200 15505
rect 8830 15370 9200 15445
rect 9230 15505 9600 15515
rect 9230 15445 9234 15505
rect 9286 15445 9544 15505
rect 9596 15445 9600 15505
rect 9230 15370 9600 15445
rect 9630 15505 10000 15515
rect 9630 15445 9634 15505
rect 9686 15445 9944 15505
rect 9996 15445 10000 15505
rect 9630 15370 10000 15445
rect 10030 15505 10400 15515
rect 10030 15445 10034 15505
rect 10086 15445 10344 15505
rect 10396 15445 10400 15505
rect 10030 15370 10400 15445
rect 10430 15505 10800 15515
rect 10430 15445 10434 15505
rect 10486 15445 10744 15505
rect 10796 15445 10800 15505
rect 10430 15370 10800 15445
rect 10830 15505 11200 15515
rect 10830 15445 10834 15505
rect 10886 15445 11144 15505
rect 11196 15445 11200 15505
rect 10830 15370 11200 15445
rect 11230 15505 11600 15515
rect 11230 15445 11234 15505
rect 11286 15445 11544 15505
rect 11596 15445 11600 15505
rect 11230 15370 11600 15445
rect 11630 15505 12000 15515
rect 11630 15445 11634 15505
rect 11686 15445 11944 15505
rect 11996 15445 12000 15505
rect 11630 15370 12000 15445
rect 12030 15505 12400 15515
rect 12030 15445 12034 15505
rect 12086 15445 12344 15505
rect 12396 15445 12400 15505
rect 12030 15370 12400 15445
rect 12430 15505 12800 15515
rect 12430 15445 12434 15505
rect 12486 15445 12744 15505
rect 12796 15445 12800 15505
rect 12430 15370 12800 15445
rect 12830 15505 13200 15515
rect 12830 15445 12834 15505
rect 12886 15445 13144 15505
rect 13196 15445 13200 15505
rect 12830 15370 13200 15445
rect 8030 15330 13200 15370
rect 8030 15245 8400 15330
rect 8030 15185 8034 15245
rect 8086 15185 8344 15245
rect 8396 15185 8400 15245
rect 8030 15175 8400 15185
rect 8430 15245 8800 15330
rect 8430 15185 8434 15245
rect 8486 15185 8744 15245
rect 8796 15185 8800 15245
rect 8430 15175 8800 15185
rect 8830 15245 9200 15330
rect 8830 15185 8834 15245
rect 8886 15185 9144 15245
rect 9196 15185 9200 15245
rect 8830 15175 9200 15185
rect 9230 15245 9600 15330
rect 9230 15185 9234 15245
rect 9286 15185 9544 15245
rect 9596 15185 9600 15245
rect 9230 15175 9600 15185
rect 9630 15245 10000 15330
rect 9630 15185 9634 15245
rect 9686 15185 9944 15245
rect 9996 15185 10000 15245
rect 9630 15175 10000 15185
rect 10030 15245 10400 15330
rect 10030 15185 10034 15245
rect 10086 15185 10344 15245
rect 10396 15185 10400 15245
rect 10030 15175 10400 15185
rect 10430 15245 10800 15330
rect 10430 15185 10434 15245
rect 10486 15185 10744 15245
rect 10796 15185 10800 15245
rect 10430 15175 10800 15185
rect 10830 15245 11200 15330
rect 10830 15185 10834 15245
rect 10886 15185 11144 15245
rect 11196 15185 11200 15245
rect 10830 15175 11200 15185
rect 11230 15245 11600 15330
rect 11230 15185 11234 15245
rect 11286 15185 11544 15245
rect 11596 15185 11600 15245
rect 11230 15175 11600 15185
rect 11630 15245 12000 15330
rect 11630 15185 11634 15245
rect 11686 15185 11944 15245
rect 11996 15185 12000 15245
rect 11630 15175 12000 15185
rect 12030 15245 12400 15330
rect 12030 15185 12034 15245
rect 12086 15185 12344 15245
rect 12396 15185 12400 15245
rect 12030 15175 12400 15185
rect 12430 15245 12800 15330
rect 12430 15185 12434 15245
rect 12486 15185 12744 15245
rect 12796 15185 12800 15245
rect 12430 15175 12800 15185
rect 12830 15245 13200 15330
rect 12830 15185 12834 15245
rect 12886 15185 13144 15245
rect 13196 15185 13200 15245
rect 12830 15175 13200 15185
rect -330 15145 -324 15175
rect 30 15145 70 15175
rect 430 15145 470 15175
rect 830 15145 870 15175
rect 1230 15145 1270 15175
rect 1630 15145 1670 15175
rect 2030 15145 2070 15175
rect 2430 15145 2470 15175
rect 2830 15145 2870 15175
rect 3230 15145 3270 15175
rect 3630 15145 3670 15175
rect 4030 15145 4070 15175
rect 4430 15145 4470 15175
rect 4830 15145 4870 15175
rect 5230 15145 5270 15175
rect 5630 15145 5670 15175
rect 6030 15145 6070 15175
rect 6430 15145 6470 15175
rect 6830 15145 6870 15175
rect 7230 15145 7270 15175
rect 7630 15145 7670 15175
rect 8030 15145 8070 15175
rect 8430 15145 8470 15175
rect 8830 15145 8870 15175
rect 9230 15145 9270 15175
rect 9630 15145 9670 15175
rect 10030 15145 10070 15175
rect 10430 15145 10470 15175
rect 10830 15145 10870 15175
rect 11230 15145 11270 15175
rect 11630 15145 11670 15175
rect 12030 15145 12070 15175
rect 12430 15145 12470 15175
rect -330 15135 0 15145
rect -314 15075 -56 15135
rect -4 15075 0 15135
rect -330 14875 0 15075
rect -314 14815 -56 14875
rect -4 14815 0 14875
rect -330 14805 0 14815
rect 30 15135 400 15145
rect 30 15075 34 15135
rect 86 15075 344 15135
rect 396 15075 400 15135
rect 30 15000 400 15075
rect 430 15135 800 15145
rect 430 15075 434 15135
rect 486 15075 744 15135
rect 796 15075 800 15135
rect 430 15000 800 15075
rect 830 15135 1200 15145
rect 830 15075 834 15135
rect 886 15075 1144 15135
rect 1196 15075 1200 15135
rect 830 15000 1200 15075
rect 1230 15135 1600 15145
rect 1230 15075 1234 15135
rect 1286 15075 1544 15135
rect 1596 15075 1600 15135
rect 1230 15000 1600 15075
rect 1630 15135 2000 15145
rect 1630 15075 1634 15135
rect 1686 15075 1944 15135
rect 1996 15075 2000 15135
rect 1630 15000 2000 15075
rect 2030 15135 2400 15145
rect 2030 15075 2034 15135
rect 2086 15075 2344 15135
rect 2396 15075 2400 15135
rect 2030 15000 2400 15075
rect 2430 15135 2800 15145
rect 2430 15075 2434 15135
rect 2486 15075 2744 15135
rect 2796 15075 2800 15135
rect 2430 15000 2800 15075
rect 2830 15135 3200 15145
rect 2830 15075 2834 15135
rect 2886 15075 3144 15135
rect 3196 15075 3200 15135
rect 2830 15000 3200 15075
rect 30 14960 3200 15000
rect 30 14875 400 14960
rect 30 14815 34 14875
rect 86 14815 344 14875
rect 396 14815 400 14875
rect 30 14805 400 14815
rect 430 14875 800 14960
rect 430 14815 434 14875
rect 486 14815 744 14875
rect 796 14815 800 14875
rect 430 14805 800 14815
rect 830 14875 1200 14960
rect 830 14815 834 14875
rect 886 14815 1144 14875
rect 1196 14815 1200 14875
rect 830 14805 1200 14815
rect 1230 14875 1600 14960
rect 1230 14815 1234 14875
rect 1286 14815 1544 14875
rect 1596 14815 1600 14875
rect 1230 14805 1600 14815
rect 1630 14875 2000 14960
rect 1630 14815 1634 14875
rect 1686 14815 1944 14875
rect 1996 14815 2000 14875
rect 1630 14805 2000 14815
rect 2030 14875 2400 14960
rect 2030 14815 2034 14875
rect 2086 14815 2344 14875
rect 2396 14815 2400 14875
rect 2030 14805 2400 14815
rect 2430 14875 2800 14960
rect 2430 14815 2434 14875
rect 2486 14815 2744 14875
rect 2796 14815 2800 14875
rect 2430 14805 2800 14815
rect 2830 14875 3200 14960
rect 2830 14815 2834 14875
rect 2886 14815 3144 14875
rect 3196 14815 3200 14875
rect 2830 14805 3200 14815
rect 3230 15135 3600 15145
rect 3230 15075 3234 15135
rect 3286 15075 3544 15135
rect 3596 15075 3600 15135
rect 3230 15000 3600 15075
rect 3630 15135 4000 15145
rect 3630 15075 3634 15135
rect 3686 15075 3944 15135
rect 3996 15075 4000 15135
rect 3630 15000 4000 15075
rect 4030 15135 4400 15145
rect 4030 15075 4034 15135
rect 4086 15075 4344 15135
rect 4396 15075 4400 15135
rect 4030 15000 4400 15075
rect 4430 15135 4800 15145
rect 4430 15075 4434 15135
rect 4486 15075 4744 15135
rect 4796 15075 4800 15135
rect 4430 15000 4800 15075
rect 4830 15135 5200 15145
rect 4830 15075 4834 15135
rect 4886 15075 5144 15135
rect 5196 15075 5200 15135
rect 4830 15000 5200 15075
rect 5230 15135 5600 15145
rect 5230 15075 5234 15135
rect 5286 15075 5544 15135
rect 5596 15075 5600 15135
rect 5230 15000 5600 15075
rect 5630 15135 6000 15145
rect 5630 15075 5634 15135
rect 5686 15075 5944 15135
rect 5996 15075 6000 15135
rect 5630 15000 6000 15075
rect 3230 14960 6000 15000
rect 3230 14875 3600 14960
rect 3230 14815 3234 14875
rect 3286 14815 3544 14875
rect 3596 14815 3600 14875
rect 3230 14805 3600 14815
rect 3630 14875 4000 14960
rect 3630 14815 3634 14875
rect 3686 14815 3944 14875
rect 3996 14815 4000 14875
rect 3630 14805 4000 14815
rect 4030 14875 4400 14960
rect 4030 14815 4034 14875
rect 4086 14815 4344 14875
rect 4396 14815 4400 14875
rect 4030 14805 4400 14815
rect 4430 14875 4800 14960
rect 4430 14815 4434 14875
rect 4486 14815 4744 14875
rect 4796 14815 4800 14875
rect 4430 14805 4800 14815
rect 4830 14875 5200 14960
rect 4830 14815 4834 14875
rect 4886 14815 5144 14875
rect 5196 14815 5200 14875
rect 4830 14805 5200 14815
rect 5230 14875 5600 14960
rect 5230 14815 5234 14875
rect 5286 14815 5544 14875
rect 5596 14815 5600 14875
rect 5230 14805 5600 14815
rect 5630 14875 6000 14960
rect 5630 14815 5634 14875
rect 5686 14815 5944 14875
rect 5996 14815 6000 14875
rect 5630 14805 6000 14815
rect 6030 15135 6400 15145
rect 6030 15075 6034 15135
rect 6086 15075 6344 15135
rect 6396 15075 6400 15135
rect 6030 15000 6400 15075
rect 6430 15135 6800 15145
rect 6430 15075 6434 15135
rect 6486 15075 6744 15135
rect 6796 15075 6800 15135
rect 6430 15000 6800 15075
rect 6830 15135 7200 15145
rect 6830 15075 6834 15135
rect 6886 15075 7144 15135
rect 7196 15075 7200 15135
rect 6830 15000 7200 15075
rect 7230 15135 7600 15145
rect 7230 15075 7234 15135
rect 7286 15075 7544 15135
rect 7596 15075 7600 15135
rect 7230 15000 7600 15075
rect 7630 15135 8000 15145
rect 7630 15075 7634 15135
rect 7686 15075 7944 15135
rect 7996 15075 8000 15135
rect 7630 15000 8000 15075
rect 6030 14960 8000 15000
rect 6030 14875 6400 14960
rect 6030 14815 6034 14875
rect 6086 14815 6344 14875
rect 6396 14815 6400 14875
rect 6030 14805 6400 14815
rect 6430 14875 6800 14960
rect 6430 14815 6434 14875
rect 6486 14815 6744 14875
rect 6796 14815 6800 14875
rect 6430 14805 6800 14815
rect 6830 14875 7200 14960
rect 6830 14815 6834 14875
rect 6886 14815 7144 14875
rect 7196 14815 7200 14875
rect 6830 14805 7200 14815
rect 7230 14875 7600 14960
rect 7230 14815 7234 14875
rect 7286 14815 7544 14875
rect 7596 14815 7600 14875
rect 7230 14805 7600 14815
rect 7630 14875 8000 14960
rect 7630 14815 7634 14875
rect 7686 14815 7944 14875
rect 7996 14815 8000 14875
rect 7630 14805 8000 14815
rect 8030 15135 8400 15145
rect 8030 15075 8034 15135
rect 8086 15075 8344 15135
rect 8396 15075 8400 15135
rect 8030 15000 8400 15075
rect 8430 15135 8800 15145
rect 8430 15075 8434 15135
rect 8486 15075 8744 15135
rect 8796 15075 8800 15135
rect 8430 15000 8800 15075
rect 8830 15135 9200 15145
rect 8830 15075 8834 15135
rect 8886 15075 9144 15135
rect 9196 15075 9200 15135
rect 8830 15000 9200 15075
rect 9230 15135 9600 15145
rect 9230 15075 9234 15135
rect 9286 15075 9544 15135
rect 9596 15075 9600 15135
rect 9230 15000 9600 15075
rect 9630 15135 10000 15145
rect 9630 15075 9634 15135
rect 9686 15075 9944 15135
rect 9996 15075 10000 15135
rect 9630 15000 10000 15075
rect 10030 15135 10400 15145
rect 10030 15075 10034 15135
rect 10086 15075 10344 15135
rect 10396 15075 10400 15135
rect 10030 15000 10400 15075
rect 10430 15135 10800 15145
rect 10430 15075 10434 15135
rect 10486 15075 10744 15135
rect 10796 15075 10800 15135
rect 10430 15000 10800 15075
rect 10830 15135 11200 15145
rect 10830 15075 10834 15135
rect 10886 15075 11144 15135
rect 11196 15075 11200 15135
rect 10830 15000 11200 15075
rect 11230 15135 11600 15145
rect 11230 15075 11234 15135
rect 11286 15075 11544 15135
rect 11596 15075 11600 15135
rect 11230 15000 11600 15075
rect 11630 15135 12000 15145
rect 11630 15075 11634 15135
rect 11686 15075 11944 15135
rect 11996 15075 12000 15135
rect 11630 15000 12000 15075
rect 12030 15135 12400 15145
rect 12030 15075 12034 15135
rect 12086 15075 12344 15135
rect 12396 15075 12400 15135
rect 12030 15000 12400 15075
rect 12430 15135 12800 15145
rect 12430 15075 12434 15135
rect 12486 15075 12744 15135
rect 12796 15075 12800 15135
rect 12430 15000 12800 15075
rect 12830 15135 13200 15145
rect 12830 15075 12834 15135
rect 12886 15075 13144 15135
rect 13196 15075 13200 15135
rect 12830 15000 13200 15075
rect 8030 14960 13200 15000
rect 8030 14875 8400 14960
rect 8030 14815 8034 14875
rect 8086 14815 8344 14875
rect 8396 14815 8400 14875
rect 8030 14805 8400 14815
rect 8430 14875 8800 14960
rect 8430 14815 8434 14875
rect 8486 14815 8744 14875
rect 8796 14815 8800 14875
rect 8430 14805 8800 14815
rect 8830 14875 9200 14960
rect 8830 14815 8834 14875
rect 8886 14815 9144 14875
rect 9196 14815 9200 14875
rect 8830 14805 9200 14815
rect 9230 14875 9600 14960
rect 9230 14815 9234 14875
rect 9286 14815 9544 14875
rect 9596 14815 9600 14875
rect 9230 14805 9600 14815
rect 9630 14875 10000 14960
rect 9630 14815 9634 14875
rect 9686 14815 9944 14875
rect 9996 14815 10000 14875
rect 9630 14805 10000 14815
rect 10030 14875 10400 14960
rect 10030 14815 10034 14875
rect 10086 14815 10344 14875
rect 10396 14815 10400 14875
rect 10030 14805 10400 14815
rect 10430 14875 10800 14960
rect 10430 14815 10434 14875
rect 10486 14815 10744 14875
rect 10796 14815 10800 14875
rect 10430 14805 10800 14815
rect 10830 14875 11200 14960
rect 10830 14815 10834 14875
rect 10886 14815 11144 14875
rect 11196 14815 11200 14875
rect 10830 14805 11200 14815
rect 11230 14875 11600 14960
rect 11230 14815 11234 14875
rect 11286 14815 11544 14875
rect 11596 14815 11600 14875
rect 11230 14805 11600 14815
rect 11630 14875 12000 14960
rect 11630 14815 11634 14875
rect 11686 14815 11944 14875
rect 11996 14815 12000 14875
rect 11630 14805 12000 14815
rect 12030 14875 12400 14960
rect 12030 14815 12034 14875
rect 12086 14815 12344 14875
rect 12396 14815 12400 14875
rect 12030 14805 12400 14815
rect 12430 14875 12800 14960
rect 12430 14815 12434 14875
rect 12486 14815 12744 14875
rect 12796 14815 12800 14875
rect 12430 14805 12800 14815
rect 12830 14875 13200 14960
rect 12830 14815 12834 14875
rect 12886 14815 13144 14875
rect 13196 14815 13200 14875
rect 12830 14805 13200 14815
rect -330 14775 -324 14805
rect 30 14775 70 14805
rect 430 14775 470 14805
rect 830 14775 870 14805
rect 1230 14775 1270 14805
rect 1630 14775 1670 14805
rect 2030 14775 2070 14805
rect 2430 14775 2470 14805
rect 3230 14775 3270 14805
rect 3630 14775 3670 14805
rect 4030 14775 4070 14805
rect 4430 14775 4470 14805
rect 4830 14775 4870 14805
rect 5230 14775 5270 14805
rect 5630 14775 5670 14805
rect 6030 14775 6070 14805
rect 6430 14775 6470 14805
rect 6830 14775 6870 14805
rect 7230 14775 7270 14805
rect 8030 14775 8070 14805
rect 8430 14775 8470 14805
rect 8830 14775 8870 14805
rect 9230 14775 9270 14805
rect 9630 14775 9670 14805
rect 10030 14775 10070 14805
rect 10430 14775 10470 14805
rect 10830 14775 10870 14805
rect 11230 14775 11270 14805
rect 11630 14775 11670 14805
rect 12030 14775 12070 14805
rect 12430 14775 12470 14805
rect -330 14765 0 14775
rect -314 14705 -56 14765
rect -4 14705 0 14765
rect -330 14505 0 14705
rect -314 14445 -56 14505
rect -4 14445 0 14505
rect -330 14435 0 14445
rect 30 14765 400 14775
rect 30 14705 34 14765
rect 86 14705 344 14765
rect 396 14705 400 14765
rect 30 14630 400 14705
rect 430 14765 800 14775
rect 430 14705 434 14765
rect 486 14705 744 14765
rect 796 14705 800 14765
rect 430 14630 800 14705
rect 830 14765 1200 14775
rect 830 14705 834 14765
rect 886 14705 1144 14765
rect 1196 14705 1200 14765
rect 830 14630 1200 14705
rect 1230 14765 1600 14775
rect 1230 14705 1234 14765
rect 1286 14705 1544 14765
rect 1596 14705 1600 14765
rect 1230 14630 1600 14705
rect 1630 14765 2000 14775
rect 1630 14705 1634 14765
rect 1686 14705 1944 14765
rect 1996 14705 2000 14765
rect 1630 14630 2000 14705
rect 2030 14765 2400 14775
rect 2030 14705 2034 14765
rect 2086 14705 2344 14765
rect 2396 14705 2400 14765
rect 2030 14630 2400 14705
rect 2430 14765 2800 14775
rect 2430 14705 2434 14765
rect 2486 14705 2744 14765
rect 2796 14705 2800 14765
rect 2430 14630 2800 14705
rect 30 14590 2800 14630
rect 30 14505 400 14590
rect 30 14445 34 14505
rect 86 14445 344 14505
rect 396 14445 400 14505
rect 30 14435 400 14445
rect 430 14505 800 14590
rect 430 14445 434 14505
rect 486 14445 744 14505
rect 796 14445 800 14505
rect 430 14435 800 14445
rect 830 14505 1200 14590
rect 830 14445 834 14505
rect 886 14445 1144 14505
rect 1196 14445 1200 14505
rect 830 14435 1200 14445
rect 1230 14505 1600 14590
rect 1230 14445 1234 14505
rect 1286 14445 1544 14505
rect 1596 14445 1600 14505
rect 1230 14435 1600 14445
rect 1630 14505 2000 14590
rect 1630 14445 1634 14505
rect 1686 14445 1944 14505
rect 1996 14445 2000 14505
rect 1630 14435 2000 14445
rect 2030 14505 2400 14590
rect 2030 14445 2034 14505
rect 2086 14445 2344 14505
rect 2396 14445 2400 14505
rect 2030 14435 2400 14445
rect 2430 14505 2800 14590
rect 2430 14445 2434 14505
rect 2486 14445 2744 14505
rect 2796 14445 2800 14505
rect 2430 14435 2800 14445
rect 2830 14765 3200 14775
rect 2830 14705 2834 14765
rect 2886 14705 3144 14765
rect 3196 14705 3200 14765
rect 2830 14630 3200 14705
rect 3230 14765 3600 14775
rect 3230 14705 3234 14765
rect 3286 14705 3544 14765
rect 3596 14705 3600 14765
rect 3230 14630 3600 14705
rect 3630 14765 4000 14775
rect 3630 14705 3634 14765
rect 3686 14705 3944 14765
rect 3996 14705 4000 14765
rect 3630 14630 4000 14705
rect 4030 14765 4400 14775
rect 4030 14705 4034 14765
rect 4086 14705 4344 14765
rect 4396 14705 4400 14765
rect 4030 14630 4400 14705
rect 4430 14765 4800 14775
rect 4430 14705 4434 14765
rect 4486 14705 4744 14765
rect 4796 14705 4800 14765
rect 4430 14630 4800 14705
rect 4830 14765 5200 14775
rect 4830 14705 4834 14765
rect 4886 14705 5144 14765
rect 5196 14705 5200 14765
rect 4830 14630 5200 14705
rect 5230 14765 5600 14775
rect 5230 14705 5234 14765
rect 5286 14705 5544 14765
rect 5596 14705 5600 14765
rect 5230 14630 5600 14705
rect 5630 14765 6000 14775
rect 5630 14705 5634 14765
rect 5686 14705 5944 14765
rect 5996 14705 6000 14765
rect 5630 14630 6000 14705
rect 2830 14590 6000 14630
rect 2830 14505 3200 14590
rect 2830 14445 2834 14505
rect 2886 14445 3144 14505
rect 3196 14445 3200 14505
rect 2830 14435 3200 14445
rect 3230 14505 3600 14590
rect 3230 14445 3234 14505
rect 3286 14445 3544 14505
rect 3596 14445 3600 14505
rect 3230 14435 3600 14445
rect 3630 14505 4000 14590
rect 3630 14445 3634 14505
rect 3686 14445 3944 14505
rect 3996 14445 4000 14505
rect 3630 14435 4000 14445
rect 4030 14505 4400 14590
rect 4030 14445 4034 14505
rect 4086 14445 4344 14505
rect 4396 14445 4400 14505
rect 4030 14435 4400 14445
rect 4430 14505 4800 14590
rect 4430 14445 4434 14505
rect 4486 14445 4744 14505
rect 4796 14445 4800 14505
rect 4430 14435 4800 14445
rect 4830 14505 5200 14590
rect 4830 14445 4834 14505
rect 4886 14445 5144 14505
rect 5196 14445 5200 14505
rect 4830 14435 5200 14445
rect 5230 14505 5600 14590
rect 5230 14445 5234 14505
rect 5286 14445 5544 14505
rect 5596 14445 5600 14505
rect 5230 14435 5600 14445
rect 5630 14505 6000 14590
rect 5630 14445 5634 14505
rect 5686 14445 5944 14505
rect 5996 14445 6000 14505
rect 5630 14435 6000 14445
rect 6030 14765 6400 14775
rect 6030 14705 6034 14765
rect 6086 14705 6344 14765
rect 6396 14705 6400 14765
rect 6030 14630 6400 14705
rect 6430 14765 6800 14775
rect 6430 14705 6434 14765
rect 6486 14705 6744 14765
rect 6796 14705 6800 14765
rect 6430 14630 6800 14705
rect 6830 14765 7200 14775
rect 6830 14705 6834 14765
rect 6886 14705 7144 14765
rect 7196 14705 7200 14765
rect 6830 14630 7200 14705
rect 7230 14765 7600 14775
rect 7230 14705 7234 14765
rect 7286 14705 7544 14765
rect 7596 14705 7600 14765
rect 7230 14630 7600 14705
rect 6030 14590 7600 14630
rect 6030 14505 6400 14590
rect 6030 14445 6034 14505
rect 6086 14445 6344 14505
rect 6396 14445 6400 14505
rect 6030 14435 6400 14445
rect 6430 14505 6800 14590
rect 6430 14445 6434 14505
rect 6486 14445 6744 14505
rect 6796 14445 6800 14505
rect 6430 14435 6800 14445
rect 6830 14505 7200 14590
rect 6830 14445 6834 14505
rect 6886 14445 7144 14505
rect 7196 14445 7200 14505
rect 6830 14435 7200 14445
rect 7230 14505 7600 14590
rect 7230 14445 7234 14505
rect 7286 14445 7544 14505
rect 7596 14445 7600 14505
rect 7230 14435 7600 14445
rect 7630 14765 8000 14775
rect 7630 14705 7634 14765
rect 7686 14705 7944 14765
rect 7996 14705 8000 14765
rect 7630 14630 8000 14705
rect 8030 14765 8400 14775
rect 8030 14705 8034 14765
rect 8086 14705 8344 14765
rect 8396 14705 8400 14765
rect 8030 14630 8400 14705
rect 8430 14765 8800 14775
rect 8430 14705 8434 14765
rect 8486 14705 8744 14765
rect 8796 14705 8800 14765
rect 8430 14630 8800 14705
rect 8830 14765 9200 14775
rect 8830 14705 8834 14765
rect 8886 14705 9144 14765
rect 9196 14705 9200 14765
rect 8830 14630 9200 14705
rect 9230 14765 9600 14775
rect 9230 14705 9234 14765
rect 9286 14705 9544 14765
rect 9596 14705 9600 14765
rect 9230 14630 9600 14705
rect 9630 14765 10000 14775
rect 9630 14705 9634 14765
rect 9686 14705 9944 14765
rect 9996 14705 10000 14765
rect 9630 14630 10000 14705
rect 10030 14765 10400 14775
rect 10030 14705 10034 14765
rect 10086 14705 10344 14765
rect 10396 14705 10400 14765
rect 10030 14630 10400 14705
rect 10430 14765 10800 14775
rect 10430 14705 10434 14765
rect 10486 14705 10744 14765
rect 10796 14705 10800 14765
rect 10430 14630 10800 14705
rect 10830 14765 11200 14775
rect 10830 14705 10834 14765
rect 10886 14705 11144 14765
rect 11196 14705 11200 14765
rect 10830 14630 11200 14705
rect 11230 14765 11600 14775
rect 11230 14705 11234 14765
rect 11286 14705 11544 14765
rect 11596 14705 11600 14765
rect 11230 14630 11600 14705
rect 11630 14765 12000 14775
rect 11630 14705 11634 14765
rect 11686 14705 11944 14765
rect 11996 14705 12000 14765
rect 11630 14630 12000 14705
rect 12030 14765 12400 14775
rect 12030 14705 12034 14765
rect 12086 14705 12344 14765
rect 12396 14705 12400 14765
rect 12030 14630 12400 14705
rect 12430 14765 12800 14775
rect 12430 14705 12434 14765
rect 12486 14705 12744 14765
rect 12796 14705 12800 14765
rect 12430 14630 12800 14705
rect 12830 14765 13200 14775
rect 12830 14705 12834 14765
rect 12886 14705 13144 14765
rect 13196 14705 13200 14765
rect 12830 14630 13200 14705
rect 7630 14590 13200 14630
rect 7630 14505 8000 14590
rect 7630 14445 7634 14505
rect 7686 14445 7944 14505
rect 7996 14445 8000 14505
rect 7630 14435 8000 14445
rect 8030 14505 8400 14590
rect 8030 14445 8034 14505
rect 8086 14445 8344 14505
rect 8396 14445 8400 14505
rect 8030 14435 8400 14445
rect 8430 14505 8800 14590
rect 8430 14445 8434 14505
rect 8486 14445 8744 14505
rect 8796 14445 8800 14505
rect 8430 14435 8800 14445
rect 8830 14505 9200 14590
rect 8830 14445 8834 14505
rect 8886 14445 9144 14505
rect 9196 14445 9200 14505
rect 8830 14435 9200 14445
rect 9230 14505 9600 14590
rect 9230 14445 9234 14505
rect 9286 14445 9544 14505
rect 9596 14445 9600 14505
rect 9230 14435 9600 14445
rect 9630 14505 10000 14590
rect 9630 14445 9634 14505
rect 9686 14445 9944 14505
rect 9996 14445 10000 14505
rect 9630 14435 10000 14445
rect 10030 14505 10400 14590
rect 10030 14445 10034 14505
rect 10086 14445 10344 14505
rect 10396 14445 10400 14505
rect 10030 14435 10400 14445
rect 10430 14505 10800 14590
rect 10430 14445 10434 14505
rect 10486 14445 10744 14505
rect 10796 14445 10800 14505
rect 10430 14435 10800 14445
rect 10830 14505 11200 14590
rect 10830 14445 10834 14505
rect 10886 14445 11144 14505
rect 11196 14445 11200 14505
rect 10830 14435 11200 14445
rect 11230 14505 11600 14590
rect 11230 14445 11234 14505
rect 11286 14445 11544 14505
rect 11596 14445 11600 14505
rect 11230 14435 11600 14445
rect 11630 14505 12000 14590
rect 11630 14445 11634 14505
rect 11686 14445 11944 14505
rect 11996 14445 12000 14505
rect 11630 14435 12000 14445
rect 12030 14505 12400 14590
rect 12030 14445 12034 14505
rect 12086 14445 12344 14505
rect 12396 14445 12400 14505
rect 12030 14435 12400 14445
rect 12430 14505 12800 14590
rect 12430 14445 12434 14505
rect 12486 14445 12744 14505
rect 12796 14445 12800 14505
rect 12430 14435 12800 14445
rect 12830 14505 13200 14590
rect 12830 14445 12834 14505
rect 12886 14445 13144 14505
rect 13196 14445 13200 14505
rect 12830 14435 13200 14445
rect -330 14405 -324 14435
rect 30 14405 70 14435
rect 430 14405 470 14435
rect 830 14405 870 14435
rect 1230 14405 1270 14435
rect 1630 14405 1670 14435
rect 2030 14405 2070 14435
rect 2430 14405 2470 14435
rect 2830 14405 2870 14435
rect 3230 14405 3270 14435
rect 3630 14405 3670 14435
rect 4030 14405 4070 14435
rect 4430 14405 4470 14435
rect 4830 14405 4870 14435
rect 5230 14405 5270 14435
rect 5630 14405 5670 14435
rect 6030 14405 6070 14435
rect 6430 14405 6470 14435
rect 6830 14405 6870 14435
rect 7230 14405 7270 14435
rect 7630 14405 7670 14435
rect 8030 14405 8070 14435
rect 8430 14405 8470 14435
rect 8830 14405 8870 14435
rect -330 14395 0 14405
rect -314 14335 -56 14395
rect -4 14335 0 14395
rect -330 14135 0 14335
rect -314 14075 -56 14135
rect -4 14075 0 14135
rect -330 14065 0 14075
rect 30 14395 400 14405
rect 30 14335 34 14395
rect 86 14335 344 14395
rect 396 14335 400 14395
rect 30 14260 400 14335
rect 430 14395 800 14405
rect 430 14335 434 14395
rect 486 14335 744 14395
rect 796 14335 800 14395
rect 430 14260 800 14335
rect 830 14395 1200 14405
rect 830 14335 834 14395
rect 886 14335 1144 14395
rect 1196 14335 1200 14395
rect 830 14260 1200 14335
rect 1230 14395 1600 14405
rect 1230 14335 1234 14395
rect 1286 14335 1544 14395
rect 1596 14335 1600 14395
rect 1230 14260 1600 14335
rect 1630 14395 2000 14405
rect 1630 14335 1634 14395
rect 1686 14335 1944 14395
rect 1996 14335 2000 14395
rect 1630 14260 2000 14335
rect 2030 14395 2400 14405
rect 2030 14335 2034 14395
rect 2086 14335 2344 14395
rect 2396 14335 2400 14395
rect 2030 14260 2400 14335
rect 2430 14395 2800 14405
rect 2430 14335 2434 14395
rect 2486 14335 2744 14395
rect 2796 14335 2800 14395
rect 2430 14260 2800 14335
rect 30 14220 2800 14260
rect 30 14135 400 14220
rect 30 14075 34 14135
rect 86 14075 344 14135
rect 396 14075 400 14135
rect 30 14065 400 14075
rect 430 14135 800 14220
rect 430 14075 434 14135
rect 486 14075 744 14135
rect 796 14075 800 14135
rect 430 14065 800 14075
rect 830 14135 1200 14220
rect 830 14075 834 14135
rect 886 14075 1144 14135
rect 1196 14075 1200 14135
rect 830 14065 1200 14075
rect 1230 14135 1600 14220
rect 1230 14075 1234 14135
rect 1286 14075 1544 14135
rect 1596 14075 1600 14135
rect 1230 14065 1600 14075
rect 1630 14135 2000 14220
rect 1630 14075 1634 14135
rect 1686 14075 1944 14135
rect 1996 14075 2000 14135
rect 1630 14065 2000 14075
rect 2030 14135 2400 14220
rect 2030 14075 2034 14135
rect 2086 14075 2344 14135
rect 2396 14075 2400 14135
rect 2030 14065 2400 14075
rect 2430 14135 2800 14220
rect 2430 14075 2434 14135
rect 2486 14075 2744 14135
rect 2796 14075 2800 14135
rect 2430 14065 2800 14075
rect 2830 14395 3200 14405
rect 2830 14335 2834 14395
rect 2886 14335 3144 14395
rect 3196 14335 3200 14395
rect 2830 14260 3200 14335
rect 3230 14395 3600 14405
rect 3230 14335 3234 14395
rect 3286 14335 3544 14395
rect 3596 14335 3600 14395
rect 3230 14260 3600 14335
rect 3630 14395 4000 14405
rect 3630 14335 3634 14395
rect 3686 14335 3944 14395
rect 3996 14335 4000 14395
rect 3630 14260 4000 14335
rect 4030 14395 4400 14405
rect 4030 14335 4034 14395
rect 4086 14335 4344 14395
rect 4396 14335 4400 14395
rect 4030 14260 4400 14335
rect 4430 14395 4800 14405
rect 4430 14335 4434 14395
rect 4486 14335 4744 14395
rect 4796 14335 4800 14395
rect 4430 14260 4800 14335
rect 4830 14395 5200 14405
rect 4830 14335 4834 14395
rect 4886 14335 5144 14395
rect 5196 14335 5200 14395
rect 4830 14260 5200 14335
rect 5230 14395 5600 14405
rect 5230 14335 5234 14395
rect 5286 14335 5544 14395
rect 5596 14335 5600 14395
rect 5230 14260 5600 14335
rect 5630 14395 6000 14405
rect 5630 14335 5634 14395
rect 5686 14335 5944 14395
rect 5996 14335 6000 14395
rect 5630 14260 6000 14335
rect 2830 14220 6000 14260
rect 2830 14135 3200 14220
rect 2830 14075 2834 14135
rect 2886 14075 3144 14135
rect 3196 14075 3200 14135
rect 2830 14065 3200 14075
rect 3230 14135 3600 14220
rect 3230 14075 3234 14135
rect 3286 14075 3544 14135
rect 3596 14075 3600 14135
rect 3230 14065 3600 14075
rect 3630 14135 4000 14220
rect 3630 14075 3634 14135
rect 3686 14075 3944 14135
rect 3996 14075 4000 14135
rect 3630 14065 4000 14075
rect 4030 14135 4400 14220
rect 4030 14075 4034 14135
rect 4086 14075 4344 14135
rect 4396 14075 4400 14135
rect 4030 14065 4400 14075
rect 4430 14135 4800 14220
rect 4430 14075 4434 14135
rect 4486 14075 4744 14135
rect 4796 14075 4800 14135
rect 4430 14065 4800 14075
rect 4830 14135 5200 14220
rect 4830 14075 4834 14135
rect 4886 14075 5144 14135
rect 5196 14075 5200 14135
rect 4830 14065 5200 14075
rect 5230 14135 5600 14220
rect 5230 14075 5234 14135
rect 5286 14075 5544 14135
rect 5596 14075 5600 14135
rect 5230 14065 5600 14075
rect 5630 14135 6000 14220
rect 5630 14075 5634 14135
rect 5686 14075 5944 14135
rect 5996 14075 6000 14135
rect 5630 14065 6000 14075
rect 6030 14395 6400 14405
rect 6030 14335 6034 14395
rect 6086 14335 6344 14395
rect 6396 14335 6400 14395
rect 6030 14260 6400 14335
rect 6430 14395 6800 14405
rect 6430 14335 6434 14395
rect 6486 14335 6744 14395
rect 6796 14335 6800 14395
rect 6430 14260 6800 14335
rect 6830 14395 7200 14405
rect 6830 14335 6834 14395
rect 6886 14335 7144 14395
rect 7196 14335 7200 14395
rect 6830 14260 7200 14335
rect 7230 14395 7600 14405
rect 7230 14335 7234 14395
rect 7286 14335 7544 14395
rect 7596 14335 7600 14395
rect 7230 14260 7600 14335
rect 6030 14220 7600 14260
rect 6030 14135 6400 14220
rect 6030 14075 6034 14135
rect 6086 14075 6344 14135
rect 6396 14075 6400 14135
rect 6030 14065 6400 14075
rect 6430 14135 6800 14220
rect 6430 14075 6434 14135
rect 6486 14075 6744 14135
rect 6796 14075 6800 14135
rect 6430 14065 6800 14075
rect 6830 14135 7200 14220
rect 6830 14075 6834 14135
rect 6886 14075 7144 14135
rect 7196 14075 7200 14135
rect 6830 14065 7200 14075
rect 7230 14135 7600 14220
rect 7230 14075 7234 14135
rect 7286 14075 7544 14135
rect 7596 14075 7600 14135
rect 7230 14065 7600 14075
rect 7630 14395 8000 14405
rect 7630 14335 7634 14395
rect 7686 14335 7944 14395
rect 7996 14335 8000 14395
rect 7630 14260 8000 14335
rect 8030 14395 8400 14405
rect 8030 14335 8034 14395
rect 8086 14335 8344 14395
rect 8396 14335 8400 14395
rect 8030 14260 8400 14335
rect 7630 14220 8400 14260
rect 7630 14135 8000 14220
rect 7630 14075 7634 14135
rect 7686 14075 7944 14135
rect 7996 14075 8000 14135
rect 7630 14065 8000 14075
rect 8030 14135 8400 14220
rect 8030 14075 8034 14135
rect 8086 14075 8344 14135
rect 8396 14075 8400 14135
rect 8030 14065 8400 14075
rect 8430 14395 8800 14405
rect 8430 14335 8434 14395
rect 8486 14335 8744 14395
rect 8796 14335 8800 14395
rect 8430 14135 8800 14335
rect 8430 14075 8434 14135
rect 8486 14075 8744 14135
rect 8796 14075 8800 14135
rect 8430 14065 8800 14075
rect 8830 14395 9200 14405
rect 8830 14335 8834 14395
rect 8886 14335 9144 14395
rect 9196 14335 9200 14395
rect 8830 14135 9200 14335
rect 8830 14075 8834 14135
rect 8886 14075 9144 14135
rect 9196 14075 9200 14135
rect 8830 14065 9200 14075
rect 9230 14395 9600 14405
rect 9230 14335 9234 14395
rect 9286 14335 9544 14395
rect 9596 14335 9600 14395
rect 9230 14260 9600 14335
rect 9630 14395 10000 14405
rect 9630 14335 9634 14395
rect 9686 14335 9944 14395
rect 9996 14335 10000 14395
rect 9630 14260 10000 14335
rect 10030 14395 10400 14405
rect 10030 14335 10034 14395
rect 10086 14335 10344 14395
rect 10396 14335 10400 14395
rect 10030 14260 10400 14335
rect 10430 14395 10800 14405
rect 10430 14335 10434 14395
rect 10486 14335 10744 14395
rect 10796 14335 10800 14395
rect 10430 14260 10800 14335
rect 10830 14395 11200 14405
rect 10830 14335 10834 14395
rect 10886 14335 11144 14395
rect 11196 14335 11200 14395
rect 10830 14260 11200 14335
rect 11230 14395 11600 14405
rect 11230 14335 11234 14395
rect 11286 14335 11544 14395
rect 11596 14335 11600 14395
rect 11230 14260 11600 14335
rect 11630 14395 12000 14405
rect 11630 14335 11634 14395
rect 11686 14335 11944 14395
rect 11996 14335 12000 14395
rect 11630 14260 12000 14335
rect 12030 14395 12400 14405
rect 12030 14335 12034 14395
rect 12086 14335 12344 14395
rect 12396 14335 12400 14395
rect 12030 14260 12400 14335
rect 12430 14395 12800 14405
rect 12430 14335 12434 14395
rect 12486 14335 12744 14395
rect 12796 14335 12800 14395
rect 12430 14260 12800 14335
rect 12830 14395 13200 14405
rect 12830 14335 12834 14395
rect 12886 14335 13144 14395
rect 13196 14335 13200 14395
rect 12830 14260 13200 14335
rect 9230 14220 13200 14260
rect 9230 14135 9600 14220
rect 9230 14075 9234 14135
rect 9286 14075 9544 14135
rect 9596 14075 9600 14135
rect 9230 14065 9600 14075
rect 9630 14135 10000 14220
rect 9630 14075 9634 14135
rect 9686 14075 9944 14135
rect 9996 14075 10000 14135
rect 9630 14065 10000 14075
rect 10030 14135 10400 14220
rect 10030 14075 10034 14135
rect 10086 14075 10344 14135
rect 10396 14075 10400 14135
rect 10030 14065 10400 14075
rect 10430 14135 10800 14220
rect 10430 14075 10434 14135
rect 10486 14075 10744 14135
rect 10796 14075 10800 14135
rect 10430 14065 10800 14075
rect 10830 14135 11200 14220
rect 10830 14075 10834 14135
rect 10886 14075 11144 14135
rect 11196 14075 11200 14135
rect 10830 14065 11200 14075
rect 11230 14135 11600 14220
rect 11230 14075 11234 14135
rect 11286 14075 11544 14135
rect 11596 14075 11600 14135
rect 11230 14065 11600 14075
rect 11630 14135 12000 14220
rect 11630 14075 11634 14135
rect 11686 14075 11944 14135
rect 11996 14075 12000 14135
rect 11630 14065 12000 14075
rect 12030 14135 12400 14220
rect 12030 14075 12034 14135
rect 12086 14075 12344 14135
rect 12396 14075 12400 14135
rect 12030 14065 12400 14075
rect 12430 14135 12800 14220
rect 12430 14075 12434 14135
rect 12486 14075 12744 14135
rect 12796 14075 12800 14135
rect 12430 14065 12800 14075
rect 12830 14135 13200 14220
rect 12830 14075 12834 14135
rect 12886 14075 13144 14135
rect 13196 14075 13200 14135
rect 12830 14065 13200 14075
rect -330 14035 -324 14065
rect 30 14035 70 14065
rect 430 14035 470 14065
rect 830 14035 870 14065
rect 1230 14035 1270 14065
rect 1630 14035 1670 14065
rect 2030 14035 2070 14065
rect 2430 14035 2470 14065
rect 2830 14035 2870 14065
rect 3230 14035 3270 14065
rect 3630 14035 3670 14065
rect 4030 14035 4070 14065
rect 4430 14035 4470 14065
rect 4830 14035 4870 14065
rect 5230 14035 5270 14065
rect 5630 14035 5670 14065
rect 6030 14035 6070 14065
rect 6430 14035 6470 14065
rect 6830 14035 6870 14065
rect 7230 14035 7270 14065
rect 7630 14035 7670 14065
rect 8030 14035 8070 14065
rect 8430 14035 8470 14065
rect 8830 14035 8870 14065
rect 9230 14035 9270 14065
rect 9630 14035 9670 14065
rect 10030 14035 10070 14065
rect 10430 14035 10470 14065
rect 10830 14035 10870 14065
rect 11230 14035 11270 14065
rect 11630 14035 11670 14065
rect 12030 14035 12070 14065
rect 12430 14035 12470 14065
rect -330 14025 0 14035
rect -314 13965 -56 14025
rect -4 13965 0 14025
rect -330 13765 0 13965
rect -314 13705 -56 13765
rect -4 13705 0 13765
rect -330 13695 0 13705
rect 30 14025 400 14035
rect 30 13965 34 14025
rect 86 13965 344 14025
rect 396 13965 400 14025
rect 30 13890 400 13965
rect 430 14025 800 14035
rect 430 13965 434 14025
rect 486 13965 744 14025
rect 796 13965 800 14025
rect 430 13890 800 13965
rect 830 14025 1200 14035
rect 830 13965 834 14025
rect 886 13965 1144 14025
rect 1196 13965 1200 14025
rect 830 13890 1200 13965
rect 1230 14025 1600 14035
rect 1230 13965 1234 14025
rect 1286 13965 1544 14025
rect 1596 13965 1600 14025
rect 1230 13890 1600 13965
rect 1630 14025 2000 14035
rect 1630 13965 1634 14025
rect 1686 13965 1944 14025
rect 1996 13965 2000 14025
rect 1630 13890 2000 13965
rect 2030 14025 2400 14035
rect 2030 13965 2034 14025
rect 2086 13965 2344 14025
rect 2396 13965 2400 14025
rect 2030 13890 2400 13965
rect 2430 14025 2800 14035
rect 2430 13965 2434 14025
rect 2486 13965 2744 14025
rect 2796 13965 2800 14025
rect 2430 13890 2800 13965
rect 30 13850 2800 13890
rect 30 13765 400 13850
rect 30 13705 34 13765
rect 86 13705 344 13765
rect 396 13705 400 13765
rect 30 13695 400 13705
rect 430 13765 800 13850
rect 430 13705 434 13765
rect 486 13705 744 13765
rect 796 13705 800 13765
rect 430 13695 800 13705
rect 830 13765 1200 13850
rect 830 13705 834 13765
rect 886 13705 1144 13765
rect 1196 13705 1200 13765
rect 830 13695 1200 13705
rect 1230 13765 1600 13850
rect 1230 13705 1234 13765
rect 1286 13705 1544 13765
rect 1596 13705 1600 13765
rect 1230 13695 1600 13705
rect 1630 13765 2000 13850
rect 1630 13705 1634 13765
rect 1686 13705 1944 13765
rect 1996 13705 2000 13765
rect 1630 13695 2000 13705
rect 2030 13765 2400 13850
rect 2030 13705 2034 13765
rect 2086 13705 2344 13765
rect 2396 13705 2400 13765
rect 2030 13695 2400 13705
rect 2430 13765 2800 13850
rect 2430 13705 2434 13765
rect 2486 13705 2744 13765
rect 2796 13705 2800 13765
rect 2430 13695 2800 13705
rect 2830 14025 3200 14035
rect 2830 13965 2834 14025
rect 2886 13965 3144 14025
rect 3196 13965 3200 14025
rect 2830 13890 3200 13965
rect 3230 14025 3600 14035
rect 3230 13965 3234 14025
rect 3286 13965 3544 14025
rect 3596 13965 3600 14025
rect 3230 13890 3600 13965
rect 3630 14025 4000 14035
rect 3630 13965 3634 14025
rect 3686 13965 3944 14025
rect 3996 13965 4000 14025
rect 3630 13890 4000 13965
rect 4030 14025 4400 14035
rect 4030 13965 4034 14025
rect 4086 13965 4344 14025
rect 4396 13965 4400 14025
rect 4030 13890 4400 13965
rect 4430 14025 4800 14035
rect 4430 13965 4434 14025
rect 4486 13965 4744 14025
rect 4796 13965 4800 14025
rect 4430 13890 4800 13965
rect 4830 14025 5200 14035
rect 4830 13965 4834 14025
rect 4886 13965 5144 14025
rect 5196 13965 5200 14025
rect 4830 13890 5200 13965
rect 5230 14025 5600 14035
rect 5230 13965 5234 14025
rect 5286 13965 5544 14025
rect 5596 13965 5600 14025
rect 5230 13890 5600 13965
rect 5630 14025 6000 14035
rect 5630 13965 5634 14025
rect 5686 13965 5944 14025
rect 5996 13965 6000 14025
rect 5630 13890 6000 13965
rect 2830 13850 6000 13890
rect 2830 13765 3200 13850
rect 2830 13705 2834 13765
rect 2886 13705 3144 13765
rect 3196 13705 3200 13765
rect 2830 13695 3200 13705
rect 3230 13765 3600 13850
rect 3230 13705 3234 13765
rect 3286 13705 3544 13765
rect 3596 13705 3600 13765
rect 3230 13695 3600 13705
rect 3630 13765 4000 13850
rect 3630 13705 3634 13765
rect 3686 13705 3944 13765
rect 3996 13705 4000 13765
rect 3630 13695 4000 13705
rect 4030 13765 4400 13850
rect 4030 13705 4034 13765
rect 4086 13705 4344 13765
rect 4396 13705 4400 13765
rect 4030 13695 4400 13705
rect 4430 13765 4800 13850
rect 4430 13705 4434 13765
rect 4486 13705 4744 13765
rect 4796 13705 4800 13765
rect 4430 13695 4800 13705
rect 4830 13765 5200 13850
rect 4830 13705 4834 13765
rect 4886 13705 5144 13765
rect 5196 13705 5200 13765
rect 4830 13695 5200 13705
rect 5230 13765 5600 13850
rect 5230 13705 5234 13765
rect 5286 13705 5544 13765
rect 5596 13705 5600 13765
rect 5230 13695 5600 13705
rect 5630 13765 6000 13850
rect 5630 13705 5634 13765
rect 5686 13705 5944 13765
rect 5996 13705 6000 13765
rect 5630 13695 6000 13705
rect 6030 14025 6400 14035
rect 6030 13965 6034 14025
rect 6086 13965 6344 14025
rect 6396 13965 6400 14025
rect 6030 13890 6400 13965
rect 6430 14025 6800 14035
rect 6430 13965 6434 14025
rect 6486 13965 6744 14025
rect 6796 13965 6800 14025
rect 6430 13890 6800 13965
rect 6830 14025 7200 14035
rect 6830 13965 6834 14025
rect 6886 13965 7144 14025
rect 7196 13965 7200 14025
rect 6830 13890 7200 13965
rect 7230 14025 7600 14035
rect 7230 13965 7234 14025
rect 7286 13965 7544 14025
rect 7596 13965 7600 14025
rect 7230 13890 7600 13965
rect 6030 13850 7600 13890
rect 6030 13765 6400 13850
rect 6030 13705 6034 13765
rect 6086 13705 6344 13765
rect 6396 13705 6400 13765
rect 6030 13695 6400 13705
rect 6430 13765 6800 13850
rect 6430 13705 6434 13765
rect 6486 13705 6744 13765
rect 6796 13705 6800 13765
rect 6430 13695 6800 13705
rect 6830 13765 7200 13850
rect 6830 13705 6834 13765
rect 6886 13705 7144 13765
rect 7196 13705 7200 13765
rect 6830 13695 7200 13705
rect 7230 13765 7600 13850
rect 7230 13705 7234 13765
rect 7286 13705 7544 13765
rect 7596 13705 7600 13765
rect 7230 13695 7600 13705
rect 7630 14025 8000 14035
rect 7630 13965 7634 14025
rect 7686 13965 7944 14025
rect 7996 13965 8000 14025
rect 7630 13890 8000 13965
rect 8030 14025 8400 14035
rect 8030 13965 8034 14025
rect 8086 13965 8344 14025
rect 8396 13965 8400 14025
rect 8030 13890 8400 13965
rect 7630 13850 8400 13890
rect 7630 13765 8000 13850
rect 7630 13705 7634 13765
rect 7686 13705 7944 13765
rect 7996 13705 8000 13765
rect 7630 13695 8000 13705
rect 8030 13765 8400 13850
rect 8030 13705 8034 13765
rect 8086 13705 8344 13765
rect 8396 13705 8400 13765
rect 8030 13695 8400 13705
rect 8430 14025 8800 14035
rect 8430 13965 8434 14025
rect 8486 13965 8744 14025
rect 8796 13965 8800 14025
rect 8430 13765 8800 13965
rect 8430 13705 8434 13765
rect 8486 13705 8744 13765
rect 8796 13705 8800 13765
rect 8430 13695 8800 13705
rect 8830 14025 9200 14035
rect 8830 13965 8834 14025
rect 8886 13965 9144 14025
rect 9196 13965 9200 14025
rect 8830 13765 9200 13965
rect 8830 13705 8834 13765
rect 8886 13705 9144 13765
rect 9196 13705 9200 13765
rect 8830 13695 9200 13705
rect 9230 14025 9600 14035
rect 9230 13965 9234 14025
rect 9286 13965 9544 14025
rect 9596 13965 9600 14025
rect 9230 13890 9600 13965
rect 9630 14025 10000 14035
rect 9630 13965 9634 14025
rect 9686 13965 9944 14025
rect 9996 13965 10000 14025
rect 9630 13890 10000 13965
rect 10030 14025 10400 14035
rect 10030 13965 10034 14025
rect 10086 13965 10344 14025
rect 10396 13965 10400 14025
rect 10030 13890 10400 13965
rect 10430 14025 10800 14035
rect 10430 13965 10434 14025
rect 10486 13965 10744 14025
rect 10796 13965 10800 14025
rect 10430 13890 10800 13965
rect 10830 14025 11200 14035
rect 10830 13965 10834 14025
rect 10886 13965 11144 14025
rect 11196 13965 11200 14025
rect 10830 13890 11200 13965
rect 11230 14025 11600 14035
rect 11230 13965 11234 14025
rect 11286 13965 11544 14025
rect 11596 13965 11600 14025
rect 11230 13890 11600 13965
rect 11630 14025 12000 14035
rect 11630 13965 11634 14025
rect 11686 13965 11944 14025
rect 11996 13965 12000 14025
rect 11630 13890 12000 13965
rect 12030 14025 12400 14035
rect 12030 13965 12034 14025
rect 12086 13965 12344 14025
rect 12396 13965 12400 14025
rect 12030 13890 12400 13965
rect 12430 14025 12800 14035
rect 12430 13965 12434 14025
rect 12486 13965 12744 14025
rect 12796 13965 12800 14025
rect 12430 13890 12800 13965
rect 12830 14025 13200 14035
rect 12830 13965 12834 14025
rect 12886 13965 13144 14025
rect 13196 13965 13200 14025
rect 12830 13890 13200 13965
rect 9230 13850 13200 13890
rect 9230 13765 9600 13850
rect 9230 13705 9234 13765
rect 9286 13705 9544 13765
rect 9596 13705 9600 13765
rect 9230 13695 9600 13705
rect 9630 13765 10000 13850
rect 9630 13705 9634 13765
rect 9686 13705 9944 13765
rect 9996 13705 10000 13765
rect 9630 13695 10000 13705
rect 10030 13765 10400 13850
rect 10030 13705 10034 13765
rect 10086 13705 10344 13765
rect 10396 13705 10400 13765
rect 10030 13695 10400 13705
rect 10430 13765 10800 13850
rect 10430 13705 10434 13765
rect 10486 13705 10744 13765
rect 10796 13705 10800 13765
rect 10430 13695 10800 13705
rect 10830 13765 11200 13850
rect 10830 13705 10834 13765
rect 10886 13705 11144 13765
rect 11196 13705 11200 13765
rect 10830 13695 11200 13705
rect 11230 13765 11600 13850
rect 11230 13705 11234 13765
rect 11286 13705 11544 13765
rect 11596 13705 11600 13765
rect 11230 13695 11600 13705
rect 11630 13765 12000 13850
rect 11630 13705 11634 13765
rect 11686 13705 11944 13765
rect 11996 13705 12000 13765
rect 11630 13695 12000 13705
rect 12030 13765 12400 13850
rect 12030 13705 12034 13765
rect 12086 13705 12344 13765
rect 12396 13705 12400 13765
rect 12030 13695 12400 13705
rect 12430 13765 12800 13850
rect 12430 13705 12434 13765
rect 12486 13705 12744 13765
rect 12796 13705 12800 13765
rect 12430 13695 12800 13705
rect 12830 13765 13200 13850
rect 12830 13705 12834 13765
rect 12886 13705 13144 13765
rect 13196 13705 13200 13765
rect 12830 13695 13200 13705
rect -330 13665 -324 13695
rect 30 13665 70 13695
rect 430 13665 470 13695
rect 830 13665 870 13695
rect 1230 13665 1270 13695
rect 1630 13665 1670 13695
rect 2030 13665 2070 13695
rect 2430 13665 2470 13695
rect 2830 13665 2870 13695
rect 3230 13665 3270 13695
rect 3630 13665 3670 13695
rect 4030 13665 4070 13695
rect 4430 13665 4470 13695
rect 4830 13665 4870 13695
rect 5230 13665 5270 13695
rect 5630 13665 5670 13695
rect 6030 13665 6070 13695
rect 6430 13665 6470 13695
rect 6830 13665 6870 13695
rect 7230 13665 7270 13695
rect 7630 13665 7670 13695
rect 8030 13665 8070 13695
rect 8430 13665 8470 13695
rect 8830 13665 8870 13695
rect 9230 13665 9270 13695
rect 9630 13665 9670 13695
rect 10030 13665 10070 13695
rect -330 13655 0 13665
rect -314 13595 -56 13655
rect -4 13595 0 13655
rect -330 13395 0 13595
rect -314 13335 -56 13395
rect -4 13335 0 13395
rect -330 13325 0 13335
rect 30 13655 400 13665
rect 30 13595 34 13655
rect 86 13595 344 13655
rect 396 13595 400 13655
rect 30 13520 400 13595
rect 430 13655 800 13665
rect 430 13595 434 13655
rect 486 13595 744 13655
rect 796 13595 800 13655
rect 430 13520 800 13595
rect 830 13655 1200 13665
rect 830 13595 834 13655
rect 886 13595 1144 13655
rect 1196 13595 1200 13655
rect 830 13520 1200 13595
rect 1230 13655 1600 13665
rect 1230 13595 1234 13655
rect 1286 13595 1544 13655
rect 1596 13595 1600 13655
rect 1230 13520 1600 13595
rect 1630 13655 2000 13665
rect 1630 13595 1634 13655
rect 1686 13595 1944 13655
rect 1996 13595 2000 13655
rect 1630 13520 2000 13595
rect 2030 13655 2400 13665
rect 2030 13595 2034 13655
rect 2086 13595 2344 13655
rect 2396 13595 2400 13655
rect 2030 13520 2400 13595
rect 2430 13655 2800 13665
rect 2430 13595 2434 13655
rect 2486 13595 2744 13655
rect 2796 13595 2800 13655
rect 2430 13520 2800 13595
rect 30 13480 2800 13520
rect 30 13395 400 13480
rect 30 13335 34 13395
rect 86 13335 344 13395
rect 396 13335 400 13395
rect 30 13325 400 13335
rect 430 13395 800 13480
rect 430 13335 434 13395
rect 486 13335 744 13395
rect 796 13335 800 13395
rect 430 13325 800 13335
rect 830 13395 1200 13480
rect 830 13335 834 13395
rect 886 13335 1144 13395
rect 1196 13335 1200 13395
rect 830 13325 1200 13335
rect 1230 13395 1600 13480
rect 1230 13335 1234 13395
rect 1286 13335 1544 13395
rect 1596 13335 1600 13395
rect 1230 13325 1600 13335
rect 1630 13395 2000 13480
rect 1630 13335 1634 13395
rect 1686 13335 1944 13395
rect 1996 13335 2000 13395
rect 1630 13325 2000 13335
rect 2030 13395 2400 13480
rect 2030 13335 2034 13395
rect 2086 13335 2344 13395
rect 2396 13335 2400 13395
rect 2030 13325 2400 13335
rect 2430 13395 2800 13480
rect 2430 13335 2434 13395
rect 2486 13335 2744 13395
rect 2796 13335 2800 13395
rect 2430 13325 2800 13335
rect 2830 13655 3200 13665
rect 2830 13595 2834 13655
rect 2886 13595 3144 13655
rect 3196 13595 3200 13655
rect 2830 13520 3200 13595
rect 3230 13655 3600 13665
rect 3230 13595 3234 13655
rect 3286 13595 3544 13655
rect 3596 13595 3600 13655
rect 3230 13520 3600 13595
rect 3630 13655 4000 13665
rect 3630 13595 3634 13655
rect 3686 13595 3944 13655
rect 3996 13595 4000 13655
rect 3630 13520 4000 13595
rect 4030 13655 4400 13665
rect 4030 13595 4034 13655
rect 4086 13595 4344 13655
rect 4396 13595 4400 13655
rect 4030 13520 4400 13595
rect 4430 13655 4800 13665
rect 4430 13595 4434 13655
rect 4486 13595 4744 13655
rect 4796 13595 4800 13655
rect 4430 13520 4800 13595
rect 4830 13655 5200 13665
rect 4830 13595 4834 13655
rect 4886 13595 5144 13655
rect 5196 13595 5200 13655
rect 4830 13520 5200 13595
rect 5230 13655 5600 13665
rect 5230 13595 5234 13655
rect 5286 13595 5544 13655
rect 5596 13595 5600 13655
rect 5230 13520 5600 13595
rect 5630 13655 6000 13665
rect 5630 13595 5634 13655
rect 5686 13595 5944 13655
rect 5996 13595 6000 13655
rect 5630 13520 6000 13595
rect 2830 13480 6000 13520
rect 2830 13395 3200 13480
rect 2830 13335 2834 13395
rect 2886 13335 3144 13395
rect 3196 13335 3200 13395
rect 2830 13325 3200 13335
rect 3230 13395 3600 13480
rect 3230 13335 3234 13395
rect 3286 13335 3544 13395
rect 3596 13335 3600 13395
rect 3230 13325 3600 13335
rect 3630 13395 4000 13480
rect 3630 13335 3634 13395
rect 3686 13335 3944 13395
rect 3996 13335 4000 13395
rect 3630 13325 4000 13335
rect 4030 13395 4400 13480
rect 4030 13335 4034 13395
rect 4086 13335 4344 13395
rect 4396 13335 4400 13395
rect 4030 13325 4400 13335
rect 4430 13395 4800 13480
rect 4430 13335 4434 13395
rect 4486 13335 4744 13395
rect 4796 13335 4800 13395
rect 4430 13325 4800 13335
rect 4830 13395 5200 13480
rect 4830 13335 4834 13395
rect 4886 13335 5144 13395
rect 5196 13335 5200 13395
rect 4830 13325 5200 13335
rect 5230 13395 5600 13480
rect 5230 13335 5234 13395
rect 5286 13335 5544 13395
rect 5596 13335 5600 13395
rect 5230 13325 5600 13335
rect 5630 13395 6000 13480
rect 5630 13335 5634 13395
rect 5686 13335 5944 13395
rect 5996 13335 6000 13395
rect 5630 13325 6000 13335
rect 6030 13655 6400 13665
rect 6030 13595 6034 13655
rect 6086 13595 6344 13655
rect 6396 13595 6400 13655
rect 6030 13520 6400 13595
rect 6430 13655 6800 13665
rect 6430 13595 6434 13655
rect 6486 13595 6744 13655
rect 6796 13595 6800 13655
rect 6430 13520 6800 13595
rect 6830 13655 7200 13665
rect 6830 13595 6834 13655
rect 6886 13595 7144 13655
rect 7196 13595 7200 13655
rect 6830 13520 7200 13595
rect 7230 13655 7600 13665
rect 7230 13595 7234 13655
rect 7286 13595 7544 13655
rect 7596 13595 7600 13655
rect 7230 13520 7600 13595
rect 6030 13480 7600 13520
rect 6030 13395 6400 13480
rect 6030 13335 6034 13395
rect 6086 13335 6344 13395
rect 6396 13335 6400 13395
rect 6030 13325 6400 13335
rect 6430 13395 6800 13480
rect 6430 13335 6434 13395
rect 6486 13335 6744 13395
rect 6796 13335 6800 13395
rect 6430 13325 6800 13335
rect 6830 13395 7200 13480
rect 6830 13335 6834 13395
rect 6886 13335 7144 13395
rect 7196 13335 7200 13395
rect 6830 13325 7200 13335
rect 7230 13395 7600 13480
rect 7230 13335 7234 13395
rect 7286 13335 7544 13395
rect 7596 13335 7600 13395
rect 7230 13325 7600 13335
rect 7630 13655 8000 13665
rect 7630 13595 7634 13655
rect 7686 13595 7944 13655
rect 7996 13595 8000 13655
rect 7630 13520 8000 13595
rect 8030 13655 8400 13665
rect 8030 13595 8034 13655
rect 8086 13595 8344 13655
rect 8396 13595 8400 13655
rect 8030 13520 8400 13595
rect 7630 13480 8400 13520
rect 7630 13395 8000 13480
rect 7630 13335 7634 13395
rect 7686 13335 7944 13395
rect 7996 13335 8000 13395
rect 7630 13325 8000 13335
rect 8030 13395 8400 13480
rect 8030 13335 8034 13395
rect 8086 13335 8344 13395
rect 8396 13335 8400 13395
rect 8030 13325 8400 13335
rect 8430 13655 8800 13665
rect 8430 13595 8434 13655
rect 8486 13595 8744 13655
rect 8796 13595 8800 13655
rect 8430 13395 8800 13595
rect 8430 13335 8434 13395
rect 8486 13335 8744 13395
rect 8796 13335 8800 13395
rect 8430 13325 8800 13335
rect 8830 13655 9200 13665
rect 8830 13595 8834 13655
rect 8886 13595 9144 13655
rect 9196 13595 9200 13655
rect 8830 13395 9200 13595
rect 8830 13335 8834 13395
rect 8886 13335 9144 13395
rect 9196 13335 9200 13395
rect 8830 13325 9200 13335
rect 9230 13655 9600 13665
rect 9230 13595 9234 13655
rect 9286 13595 9544 13655
rect 9596 13595 9600 13655
rect 9230 13520 9600 13595
rect 9630 13655 10000 13665
rect 9630 13595 9634 13655
rect 9686 13595 9944 13655
rect 9996 13595 10000 13655
rect 9630 13520 10000 13595
rect 10030 13655 10400 13665
rect 10030 13595 10034 13655
rect 10086 13595 10344 13655
rect 10396 13595 10400 13655
rect 10030 13520 10400 13595
rect 9230 13480 10400 13520
rect 9230 13395 9600 13480
rect 9230 13335 9234 13395
rect 9286 13335 9544 13395
rect 9596 13335 9600 13395
rect 9230 13325 9600 13335
rect 9630 13395 10000 13480
rect 9630 13335 9634 13395
rect 9686 13335 9944 13395
rect 9996 13335 10000 13395
rect 9630 13325 10000 13335
rect 10030 13395 10400 13480
rect 10030 13335 10034 13395
rect 10086 13335 10344 13395
rect 10396 13335 10400 13395
rect 10030 13325 10400 13335
rect 10430 13655 10800 13665
rect 10430 13595 10434 13655
rect 10486 13595 10744 13655
rect 10796 13595 10800 13655
rect 10430 13520 10800 13595
rect 10830 13655 11200 13665
rect 10830 13595 10834 13655
rect 10886 13595 11144 13655
rect 11196 13595 11200 13655
rect 10830 13520 11200 13595
rect 11230 13655 11600 13665
rect 11230 13595 11234 13655
rect 11286 13595 11544 13655
rect 11596 13595 11600 13655
rect 11230 13520 11600 13595
rect 11630 13655 12000 13665
rect 11630 13595 11634 13655
rect 11686 13595 11944 13655
rect 11996 13595 12000 13655
rect 11630 13520 12000 13595
rect 12030 13655 12400 13665
rect 12030 13595 12034 13655
rect 12086 13595 12344 13655
rect 12396 13595 12400 13655
rect 12030 13520 12400 13595
rect 12430 13655 12800 13665
rect 12430 13595 12434 13655
rect 12486 13595 12744 13655
rect 12796 13595 12800 13655
rect 12430 13520 12800 13595
rect 12830 13655 13200 13665
rect 12830 13595 12834 13655
rect 12886 13595 13144 13655
rect 13196 13595 13200 13655
rect 12830 13520 13200 13595
rect 10430 13480 13200 13520
rect 10430 13395 10800 13480
rect 10430 13335 10434 13395
rect 10486 13335 10744 13395
rect 10796 13335 10800 13395
rect 10430 13325 10800 13335
rect 10830 13395 11200 13480
rect 10830 13335 10834 13395
rect 10886 13335 11144 13395
rect 11196 13335 11200 13395
rect 10830 13325 11200 13335
rect 11230 13395 11600 13480
rect 11230 13335 11234 13395
rect 11286 13335 11544 13395
rect 11596 13335 11600 13395
rect 11230 13325 11600 13335
rect 11630 13395 12000 13480
rect 11630 13335 11634 13395
rect 11686 13335 11944 13395
rect 11996 13335 12000 13395
rect 11630 13325 12000 13335
rect 12030 13395 12400 13480
rect 12030 13335 12034 13395
rect 12086 13335 12344 13395
rect 12396 13335 12400 13395
rect 12030 13325 12400 13335
rect 12430 13395 12800 13480
rect 12430 13335 12434 13395
rect 12486 13335 12744 13395
rect 12796 13335 12800 13395
rect 12430 13325 12800 13335
rect 12830 13395 13200 13480
rect 12830 13335 12834 13395
rect 12886 13335 13144 13395
rect 13196 13335 13200 13395
rect 12830 13325 13200 13335
rect -330 13295 -324 13325
rect 30 13295 70 13325
rect 430 13295 470 13325
rect 830 13295 870 13325
rect 1230 13295 1270 13325
rect 1630 13295 1670 13325
rect 2030 13295 2070 13325
rect 2430 13295 2470 13325
rect 2830 13295 2870 13325
rect 3230 13295 3270 13325
rect 3630 13295 3670 13325
rect 4030 13295 4070 13325
rect 4430 13295 4470 13325
rect 4830 13295 4870 13325
rect 5230 13295 5270 13325
rect 5630 13295 5670 13325
rect 6030 13295 6070 13325
rect 6430 13295 6470 13325
rect 6830 13295 6870 13325
rect 7230 13295 7270 13325
rect 7630 13295 7670 13325
rect 8030 13295 8070 13325
rect 8430 13295 8470 13325
rect 8830 13295 8870 13325
rect 9230 13295 9270 13325
rect 9630 13295 9670 13325
rect 10030 13295 10070 13325
rect 10430 13295 10470 13325
rect 10830 13295 10870 13325
rect -330 13285 0 13295
rect -314 13225 -56 13285
rect -4 13225 0 13285
rect -330 13025 0 13225
rect -314 12965 -56 13025
rect -4 12965 0 13025
rect -330 12955 0 12965
rect 30 13285 400 13295
rect 30 13225 34 13285
rect 86 13225 344 13285
rect 396 13225 400 13285
rect 30 13150 400 13225
rect 430 13285 800 13295
rect 430 13225 434 13285
rect 486 13225 744 13285
rect 796 13225 800 13285
rect 430 13150 800 13225
rect 830 13285 1200 13295
rect 830 13225 834 13285
rect 886 13225 1144 13285
rect 1196 13225 1200 13285
rect 830 13150 1200 13225
rect 1230 13285 1600 13295
rect 1230 13225 1234 13285
rect 1286 13225 1544 13285
rect 1596 13225 1600 13285
rect 1230 13150 1600 13225
rect 1630 13285 2000 13295
rect 1630 13225 1634 13285
rect 1686 13225 1944 13285
rect 1996 13225 2000 13285
rect 1630 13150 2000 13225
rect 2030 13285 2400 13295
rect 2030 13225 2034 13285
rect 2086 13225 2344 13285
rect 2396 13225 2400 13285
rect 2030 13150 2400 13225
rect 2430 13285 2800 13295
rect 2430 13225 2434 13285
rect 2486 13225 2744 13285
rect 2796 13225 2800 13285
rect 2430 13150 2800 13225
rect 30 13110 2800 13150
rect 30 13025 400 13110
rect 30 12965 34 13025
rect 86 12965 344 13025
rect 396 12965 400 13025
rect 30 12955 400 12965
rect 430 13025 800 13110
rect 430 12965 434 13025
rect 486 12965 744 13025
rect 796 12965 800 13025
rect 430 12955 800 12965
rect 830 13025 1200 13110
rect 830 12965 834 13025
rect 886 12965 1144 13025
rect 1196 12965 1200 13025
rect 830 12955 1200 12965
rect 1230 13025 1600 13110
rect 1230 12965 1234 13025
rect 1286 12965 1544 13025
rect 1596 12965 1600 13025
rect 1230 12955 1600 12965
rect 1630 13025 2000 13110
rect 1630 12965 1634 13025
rect 1686 12965 1944 13025
rect 1996 12965 2000 13025
rect 1630 12955 2000 12965
rect 2030 13025 2400 13110
rect 2030 12965 2034 13025
rect 2086 12965 2344 13025
rect 2396 12965 2400 13025
rect 2030 12955 2400 12965
rect 2430 13025 2800 13110
rect 2430 12965 2434 13025
rect 2486 12965 2744 13025
rect 2796 12965 2800 13025
rect 2430 12955 2800 12965
rect 2830 13285 3200 13295
rect 2830 13225 2834 13285
rect 2886 13225 3144 13285
rect 3196 13225 3200 13285
rect 2830 13150 3200 13225
rect 3230 13285 3600 13295
rect 3230 13225 3234 13285
rect 3286 13225 3544 13285
rect 3596 13225 3600 13285
rect 3230 13150 3600 13225
rect 3630 13285 4000 13295
rect 3630 13225 3634 13285
rect 3686 13225 3944 13285
rect 3996 13225 4000 13285
rect 3630 13150 4000 13225
rect 4030 13285 4400 13295
rect 4030 13225 4034 13285
rect 4086 13225 4344 13285
rect 4396 13225 4400 13285
rect 4030 13150 4400 13225
rect 4430 13285 4800 13295
rect 4430 13225 4434 13285
rect 4486 13225 4744 13285
rect 4796 13225 4800 13285
rect 4430 13150 4800 13225
rect 4830 13285 5200 13295
rect 4830 13225 4834 13285
rect 4886 13225 5144 13285
rect 5196 13225 5200 13285
rect 4830 13150 5200 13225
rect 5230 13285 5600 13295
rect 5230 13225 5234 13285
rect 5286 13225 5544 13285
rect 5596 13225 5600 13285
rect 5230 13150 5600 13225
rect 5630 13285 6000 13295
rect 5630 13225 5634 13285
rect 5686 13225 5944 13285
rect 5996 13225 6000 13285
rect 5630 13150 6000 13225
rect 2830 13110 6000 13150
rect 2830 13025 3200 13110
rect 2830 12965 2834 13025
rect 2886 12965 3144 13025
rect 3196 12965 3200 13025
rect 2830 12955 3200 12965
rect 3230 13025 3600 13110
rect 3230 12965 3234 13025
rect 3286 12965 3544 13025
rect 3596 12965 3600 13025
rect 3230 12955 3600 12965
rect 3630 13025 4000 13110
rect 3630 12965 3634 13025
rect 3686 12965 3944 13025
rect 3996 12965 4000 13025
rect 3630 12955 4000 12965
rect 4030 13025 4400 13110
rect 4030 12965 4034 13025
rect 4086 12965 4344 13025
rect 4396 12965 4400 13025
rect 4030 12955 4400 12965
rect 4430 13025 4800 13110
rect 4430 12965 4434 13025
rect 4486 12965 4744 13025
rect 4796 12965 4800 13025
rect 4430 12955 4800 12965
rect 4830 13025 5200 13110
rect 4830 12965 4834 13025
rect 4886 12965 5144 13025
rect 5196 12965 5200 13025
rect 4830 12955 5200 12965
rect 5230 13025 5600 13110
rect 5230 12965 5234 13025
rect 5286 12965 5544 13025
rect 5596 12965 5600 13025
rect 5230 12955 5600 12965
rect 5630 13025 6000 13110
rect 5630 12965 5634 13025
rect 5686 12965 5944 13025
rect 5996 12965 6000 13025
rect 5630 12955 6000 12965
rect 6030 13285 6400 13295
rect 6030 13225 6034 13285
rect 6086 13225 6344 13285
rect 6396 13225 6400 13285
rect 6030 13150 6400 13225
rect 6430 13285 6800 13295
rect 6430 13225 6434 13285
rect 6486 13225 6744 13285
rect 6796 13225 6800 13285
rect 6430 13150 6800 13225
rect 6830 13285 7200 13295
rect 6830 13225 6834 13285
rect 6886 13225 7144 13285
rect 7196 13225 7200 13285
rect 6830 13150 7200 13225
rect 7230 13285 7600 13295
rect 7230 13225 7234 13285
rect 7286 13225 7544 13285
rect 7596 13225 7600 13285
rect 7230 13150 7600 13225
rect 6030 13110 7600 13150
rect 6030 13025 6400 13110
rect 6030 12965 6034 13025
rect 6086 12965 6344 13025
rect 6396 12965 6400 13025
rect 6030 12955 6400 12965
rect 6430 13025 6800 13110
rect 6430 12965 6434 13025
rect 6486 12965 6744 13025
rect 6796 12965 6800 13025
rect 6430 12955 6800 12965
rect 6830 13025 7200 13110
rect 6830 12965 6834 13025
rect 6886 12965 7144 13025
rect 7196 12965 7200 13025
rect 6830 12955 7200 12965
rect 7230 13025 7600 13110
rect 7230 12965 7234 13025
rect 7286 12965 7544 13025
rect 7596 12965 7600 13025
rect 7230 12955 7600 12965
rect 7630 13285 8000 13295
rect 7630 13225 7634 13285
rect 7686 13225 7944 13285
rect 7996 13225 8000 13285
rect 7630 13150 8000 13225
rect 8030 13285 8400 13295
rect 8030 13225 8034 13285
rect 8086 13225 8344 13285
rect 8396 13225 8400 13285
rect 8030 13150 8400 13225
rect 7630 13110 8400 13150
rect 7630 13025 8000 13110
rect 7630 12965 7634 13025
rect 7686 12965 7944 13025
rect 7996 12965 8000 13025
rect 7630 12955 8000 12965
rect 8030 13025 8400 13110
rect 8030 12965 8034 13025
rect 8086 12965 8344 13025
rect 8396 12965 8400 13025
rect 8030 12955 8400 12965
rect 8430 13285 8800 13295
rect 8430 13225 8434 13285
rect 8486 13225 8744 13285
rect 8796 13225 8800 13285
rect 8430 13025 8800 13225
rect 8430 12965 8434 13025
rect 8486 12965 8744 13025
rect 8796 12965 8800 13025
rect 8430 12955 8800 12965
rect 8830 13285 9200 13295
rect 8830 13225 8834 13285
rect 8886 13225 9144 13285
rect 9196 13225 9200 13285
rect 8830 13025 9200 13225
rect 8830 12965 8834 13025
rect 8886 12965 9144 13025
rect 9196 12965 9200 13025
rect 8830 12955 9200 12965
rect 9230 13285 9600 13295
rect 9230 13225 9234 13285
rect 9286 13225 9544 13285
rect 9596 13225 9600 13285
rect 9230 13150 9600 13225
rect 9630 13285 10000 13295
rect 9630 13225 9634 13285
rect 9686 13225 9944 13285
rect 9996 13225 10000 13285
rect 9630 13150 10000 13225
rect 10030 13285 10400 13295
rect 10030 13225 10034 13285
rect 10086 13225 10344 13285
rect 10396 13225 10400 13285
rect 10030 13150 10400 13225
rect 9230 13110 10400 13150
rect 9230 13025 9600 13110
rect 9230 12965 9234 13025
rect 9286 12965 9544 13025
rect 9596 12965 9600 13025
rect 9230 12955 9600 12965
rect 9630 13025 10000 13110
rect 9630 12965 9634 13025
rect 9686 12965 9944 13025
rect 9996 12965 10000 13025
rect 9630 12955 10000 12965
rect 10030 13025 10400 13110
rect 10030 12965 10034 13025
rect 10086 12965 10344 13025
rect 10396 12965 10400 13025
rect 10030 12955 10400 12965
rect 10430 13285 10800 13295
rect 10430 13225 10434 13285
rect 10486 13225 10744 13285
rect 10796 13225 10800 13285
rect 10430 13150 10800 13225
rect 10830 13285 11200 13295
rect 10830 13225 10834 13285
rect 10886 13225 11144 13285
rect 11196 13225 11200 13285
rect 10830 13150 11200 13225
rect 10430 13110 11200 13150
rect 10430 13025 10800 13110
rect 10430 12965 10434 13025
rect 10486 12965 10744 13025
rect 10796 12965 10800 13025
rect 10430 12955 10800 12965
rect 10830 13025 11200 13110
rect 10830 12965 10834 13025
rect 10886 12965 11144 13025
rect 11196 12965 11200 13025
rect 10830 12955 11200 12965
rect 11230 13285 11600 13295
rect 11230 13225 11234 13285
rect 11286 13225 11544 13285
rect 11596 13225 11600 13285
rect 11230 13150 11600 13225
rect 11630 13285 12000 13295
rect 11630 13225 11634 13285
rect 11686 13225 11944 13285
rect 11996 13225 12000 13285
rect 11630 13150 12000 13225
rect 12030 13285 12400 13295
rect 12030 13225 12034 13285
rect 12086 13225 12344 13285
rect 12396 13225 12400 13285
rect 12030 13150 12400 13225
rect 12430 13285 12800 13295
rect 12430 13225 12434 13285
rect 12486 13225 12744 13285
rect 12796 13225 12800 13285
rect 12430 13150 12800 13225
rect 12830 13285 13200 13295
rect 12830 13225 12834 13285
rect 12886 13225 13144 13285
rect 13196 13225 13200 13285
rect 12830 13150 13200 13225
rect 11230 13110 13200 13150
rect 11230 13025 11600 13110
rect 11230 12965 11234 13025
rect 11286 12965 11544 13025
rect 11596 12965 11600 13025
rect 11230 12955 11600 12965
rect 11630 13025 12000 13110
rect 11630 12965 11634 13025
rect 11686 12965 11944 13025
rect 11996 12965 12000 13025
rect 11630 12955 12000 12965
rect 12030 13025 12400 13110
rect 12030 12965 12034 13025
rect 12086 12965 12344 13025
rect 12396 12965 12400 13025
rect 12030 12955 12400 12965
rect 12430 13025 12800 13110
rect 12430 12965 12434 13025
rect 12486 12965 12744 13025
rect 12796 12965 12800 13025
rect 12430 12955 12800 12965
rect 12830 13025 13200 13110
rect 12830 12965 12834 13025
rect 12886 12965 13144 13025
rect 13196 12965 13200 13025
rect 12830 12955 13200 12965
rect -330 12925 -324 12955
rect 30 12925 70 12955
rect 430 12925 470 12955
rect 830 12925 870 12955
rect 1230 12925 1270 12955
rect 1630 12925 1670 12955
rect 2030 12925 2070 12955
rect 2430 12925 2470 12955
rect 2830 12925 2870 12955
rect 3230 12925 3270 12955
rect 3630 12925 3670 12955
rect 4030 12925 4070 12955
rect 4430 12925 4470 12955
rect 4830 12925 4870 12955
rect 5230 12925 5270 12955
rect 5630 12925 5670 12955
rect 6030 12925 6070 12955
rect 6430 12925 6470 12955
rect 6830 12925 6870 12955
rect 7230 12925 7270 12955
rect 7630 12925 7670 12955
rect 8030 12925 8070 12955
rect 8430 12925 8470 12955
rect 8830 12925 8870 12955
rect 9230 12925 9270 12955
rect 9630 12925 9670 12955
rect 10030 12925 10070 12955
rect 10430 12925 10470 12955
rect 10830 12925 10870 12955
rect 11230 12925 11270 12955
rect -330 12915 0 12925
rect -314 12855 -56 12915
rect -4 12855 0 12915
rect -330 12655 0 12855
rect -314 12595 -56 12655
rect -4 12595 0 12655
rect -330 12585 0 12595
rect 30 12915 400 12925
rect 30 12855 34 12915
rect 86 12855 344 12915
rect 396 12855 400 12915
rect 30 12780 400 12855
rect 430 12915 800 12925
rect 430 12855 434 12915
rect 486 12855 744 12915
rect 796 12855 800 12915
rect 430 12780 800 12855
rect 830 12915 1200 12925
rect 830 12855 834 12915
rect 886 12855 1144 12915
rect 1196 12855 1200 12915
rect 830 12780 1200 12855
rect 1230 12915 1600 12925
rect 1230 12855 1234 12915
rect 1286 12855 1544 12915
rect 1596 12855 1600 12915
rect 1230 12780 1600 12855
rect 1630 12915 2000 12925
rect 1630 12855 1634 12915
rect 1686 12855 1944 12915
rect 1996 12855 2000 12915
rect 1630 12780 2000 12855
rect 2030 12915 2400 12925
rect 2030 12855 2034 12915
rect 2086 12855 2344 12915
rect 2396 12855 2400 12915
rect 2030 12780 2400 12855
rect 2430 12915 2800 12925
rect 2430 12855 2434 12915
rect 2486 12855 2744 12915
rect 2796 12855 2800 12915
rect 2430 12780 2800 12855
rect 30 12740 2800 12780
rect 30 12655 400 12740
rect 30 12595 34 12655
rect 86 12595 344 12655
rect 396 12595 400 12655
rect 30 12585 400 12595
rect 430 12655 800 12740
rect 430 12595 434 12655
rect 486 12595 744 12655
rect 796 12595 800 12655
rect 430 12585 800 12595
rect 830 12655 1200 12740
rect 830 12595 834 12655
rect 886 12595 1144 12655
rect 1196 12595 1200 12655
rect 830 12585 1200 12595
rect 1230 12655 1600 12740
rect 1230 12595 1234 12655
rect 1286 12595 1544 12655
rect 1596 12595 1600 12655
rect 1230 12585 1600 12595
rect 1630 12655 2000 12740
rect 1630 12595 1634 12655
rect 1686 12595 1944 12655
rect 1996 12595 2000 12655
rect 1630 12585 2000 12595
rect 2030 12655 2400 12740
rect 2030 12595 2034 12655
rect 2086 12595 2344 12655
rect 2396 12595 2400 12655
rect 2030 12585 2400 12595
rect 2430 12655 2800 12740
rect 2430 12595 2434 12655
rect 2486 12595 2744 12655
rect 2796 12595 2800 12655
rect 2430 12585 2800 12595
rect 2830 12915 3200 12925
rect 2830 12855 2834 12915
rect 2886 12855 3144 12915
rect 3196 12855 3200 12915
rect 2830 12780 3200 12855
rect 3230 12915 3600 12925
rect 3230 12855 3234 12915
rect 3286 12855 3544 12915
rect 3596 12855 3600 12915
rect 3230 12780 3600 12855
rect 3630 12915 4000 12925
rect 3630 12855 3634 12915
rect 3686 12855 3944 12915
rect 3996 12855 4000 12915
rect 3630 12780 4000 12855
rect 4030 12915 4400 12925
rect 4030 12855 4034 12915
rect 4086 12855 4344 12915
rect 4396 12855 4400 12915
rect 4030 12780 4400 12855
rect 4430 12915 4800 12925
rect 4430 12855 4434 12915
rect 4486 12855 4744 12915
rect 4796 12855 4800 12915
rect 4430 12780 4800 12855
rect 4830 12915 5200 12925
rect 4830 12855 4834 12915
rect 4886 12855 5144 12915
rect 5196 12855 5200 12915
rect 4830 12780 5200 12855
rect 5230 12915 5600 12925
rect 5230 12855 5234 12915
rect 5286 12855 5544 12915
rect 5596 12855 5600 12915
rect 5230 12780 5600 12855
rect 5630 12915 6000 12925
rect 5630 12855 5634 12915
rect 5686 12855 5944 12915
rect 5996 12855 6000 12915
rect 5630 12780 6000 12855
rect 2830 12740 6000 12780
rect 2830 12655 3200 12740
rect 2830 12595 2834 12655
rect 2886 12595 3144 12655
rect 3196 12595 3200 12655
rect 2830 12585 3200 12595
rect 3230 12655 3600 12740
rect 3230 12595 3234 12655
rect 3286 12595 3544 12655
rect 3596 12595 3600 12655
rect 3230 12585 3600 12595
rect 3630 12655 4000 12740
rect 3630 12595 3634 12655
rect 3686 12595 3944 12655
rect 3996 12595 4000 12655
rect 3630 12585 4000 12595
rect 4030 12655 4400 12740
rect 4030 12595 4034 12655
rect 4086 12595 4344 12655
rect 4396 12595 4400 12655
rect 4030 12585 4400 12595
rect 4430 12655 4800 12740
rect 4430 12595 4434 12655
rect 4486 12595 4744 12655
rect 4796 12595 4800 12655
rect 4430 12585 4800 12595
rect 4830 12655 5200 12740
rect 4830 12595 4834 12655
rect 4886 12595 5144 12655
rect 5196 12595 5200 12655
rect 4830 12585 5200 12595
rect 5230 12655 5600 12740
rect 5230 12595 5234 12655
rect 5286 12595 5544 12655
rect 5596 12595 5600 12655
rect 5230 12585 5600 12595
rect 5630 12655 6000 12740
rect 5630 12595 5634 12655
rect 5686 12595 5944 12655
rect 5996 12595 6000 12655
rect 5630 12585 6000 12595
rect 6030 12915 6400 12925
rect 6030 12855 6034 12915
rect 6086 12855 6344 12915
rect 6396 12855 6400 12915
rect 6030 12780 6400 12855
rect 6430 12915 6800 12925
rect 6430 12855 6434 12915
rect 6486 12855 6744 12915
rect 6796 12855 6800 12915
rect 6430 12780 6800 12855
rect 6830 12915 7200 12925
rect 6830 12855 6834 12915
rect 6886 12855 7144 12915
rect 7196 12855 7200 12915
rect 6830 12780 7200 12855
rect 7230 12915 7600 12925
rect 7230 12855 7234 12915
rect 7286 12855 7544 12915
rect 7596 12855 7600 12915
rect 7230 12780 7600 12855
rect 6030 12740 7600 12780
rect 6030 12655 6400 12740
rect 6030 12595 6034 12655
rect 6086 12595 6344 12655
rect 6396 12595 6400 12655
rect 6030 12585 6400 12595
rect 6430 12655 6800 12740
rect 6430 12595 6434 12655
rect 6486 12595 6744 12655
rect 6796 12595 6800 12655
rect 6430 12585 6800 12595
rect 6830 12655 7200 12740
rect 6830 12595 6834 12655
rect 6886 12595 7144 12655
rect 7196 12595 7200 12655
rect 6830 12585 7200 12595
rect 7230 12655 7600 12740
rect 7230 12595 7234 12655
rect 7286 12595 7544 12655
rect 7596 12595 7600 12655
rect 7230 12585 7600 12595
rect 7630 12915 8000 12925
rect 7630 12855 7634 12915
rect 7686 12855 7944 12915
rect 7996 12855 8000 12915
rect 7630 12780 8000 12855
rect 8030 12915 8400 12925
rect 8030 12855 8034 12915
rect 8086 12855 8344 12915
rect 8396 12855 8400 12915
rect 8030 12780 8400 12855
rect 7630 12740 8400 12780
rect 7630 12655 8000 12740
rect 7630 12595 7634 12655
rect 7686 12595 7944 12655
rect 7996 12595 8000 12655
rect 7630 12585 8000 12595
rect 8030 12655 8400 12740
rect 8030 12595 8034 12655
rect 8086 12595 8344 12655
rect 8396 12595 8400 12655
rect 8030 12585 8400 12595
rect 8430 12915 8800 12925
rect 8430 12855 8434 12915
rect 8486 12855 8744 12915
rect 8796 12855 8800 12915
rect 8430 12655 8800 12855
rect 8430 12595 8434 12655
rect 8486 12595 8744 12655
rect 8796 12595 8800 12655
rect 8430 12585 8800 12595
rect 8830 12915 9200 12925
rect 8830 12855 8834 12915
rect 8886 12855 9144 12915
rect 9196 12855 9200 12915
rect 8830 12655 9200 12855
rect 8830 12595 8834 12655
rect 8886 12595 9144 12655
rect 9196 12595 9200 12655
rect 8830 12585 9200 12595
rect 9230 12915 9600 12925
rect 9230 12855 9234 12915
rect 9286 12855 9544 12915
rect 9596 12855 9600 12915
rect 9230 12780 9600 12855
rect 9630 12915 10000 12925
rect 9630 12855 9634 12915
rect 9686 12855 9944 12915
rect 9996 12855 10000 12915
rect 9630 12780 10000 12855
rect 10030 12915 10400 12925
rect 10030 12855 10034 12915
rect 10086 12855 10344 12915
rect 10396 12855 10400 12915
rect 10030 12780 10400 12855
rect 9230 12740 10400 12780
rect 9230 12655 9600 12740
rect 9230 12595 9234 12655
rect 9286 12595 9544 12655
rect 9596 12595 9600 12655
rect 9230 12585 9600 12595
rect 9630 12655 10000 12740
rect 9630 12595 9634 12655
rect 9686 12595 9944 12655
rect 9996 12595 10000 12655
rect 9630 12585 10000 12595
rect 10030 12655 10400 12740
rect 10030 12595 10034 12655
rect 10086 12595 10344 12655
rect 10396 12595 10400 12655
rect 10030 12585 10400 12595
rect 10430 12915 10800 12925
rect 10430 12855 10434 12915
rect 10486 12855 10744 12915
rect 10796 12855 10800 12915
rect 10430 12780 10800 12855
rect 10830 12915 11200 12925
rect 10830 12855 10834 12915
rect 10886 12855 11144 12915
rect 11196 12855 11200 12915
rect 10830 12780 11200 12855
rect 10430 12740 11200 12780
rect 10430 12655 10800 12740
rect 10430 12595 10434 12655
rect 10486 12595 10744 12655
rect 10796 12595 10800 12655
rect 10430 12585 10800 12595
rect 10830 12655 11200 12740
rect 10830 12595 10834 12655
rect 10886 12595 11144 12655
rect 11196 12595 11200 12655
rect 10830 12585 11200 12595
rect 11230 12915 11600 12925
rect 11230 12855 11234 12915
rect 11286 12855 11544 12915
rect 11596 12855 11600 12915
rect 11230 12655 11600 12855
rect 11230 12595 11234 12655
rect 11286 12595 11544 12655
rect 11596 12595 11600 12655
rect 11230 12585 11600 12595
rect 11630 12915 12000 12925
rect 11630 12855 11634 12915
rect 11686 12855 11944 12915
rect 11996 12855 12000 12915
rect 11630 12780 12000 12855
rect 12030 12915 12400 12925
rect 12030 12855 12034 12915
rect 12086 12855 12344 12915
rect 12396 12855 12400 12915
rect 12030 12780 12400 12855
rect 12430 12915 12800 12925
rect 12430 12855 12434 12915
rect 12486 12855 12744 12915
rect 12796 12855 12800 12915
rect 12430 12780 12800 12855
rect 12830 12915 13200 12925
rect 12830 12855 12834 12915
rect 12886 12855 13144 12915
rect 13196 12855 13200 12915
rect 12830 12780 13200 12855
rect 11630 12740 13390 12780
rect 11630 12655 12000 12740
rect 11630 12595 11634 12655
rect 11686 12595 11944 12655
rect 11996 12595 12000 12655
rect 11630 12585 12000 12595
rect 12030 12655 12400 12740
rect 12030 12595 12034 12655
rect 12086 12595 12344 12655
rect 12396 12595 12400 12655
rect 12030 12585 12400 12595
rect 12430 12655 12800 12740
rect 12430 12595 12434 12655
rect 12486 12595 12744 12655
rect 12796 12595 12800 12655
rect 12430 12585 12800 12595
rect 12830 12655 13200 12740
rect 12830 12595 12834 12655
rect 12886 12595 13144 12655
rect 13196 12595 13200 12655
rect 12830 12585 13200 12595
rect -330 12555 -324 12585
rect 30 12555 70 12585
rect 430 12555 470 12585
rect 830 12555 870 12585
rect 1230 12555 1270 12585
rect 1630 12555 1670 12585
rect 2030 12555 2070 12585
rect 2430 12555 2470 12585
rect 2830 12555 2870 12585
rect 3230 12555 3270 12585
rect 3630 12555 3670 12585
rect 4030 12555 4070 12585
rect 4430 12555 4470 12585
rect 4830 12555 4870 12585
rect 5230 12555 5270 12585
rect 5630 12555 5670 12585
rect 6030 12555 6070 12585
rect 6430 12555 6470 12585
rect 6830 12555 6870 12585
rect 7230 12555 7270 12585
rect 7630 12555 7670 12585
rect 8030 12555 8070 12585
rect 8430 12555 8470 12585
rect 8830 12555 8870 12585
rect 9230 12555 9270 12585
rect 9630 12555 9670 12585
rect 10430 12555 10470 12585
rect 10830 12555 10870 12585
rect 11230 12555 11270 12585
rect 11630 12555 11670 12585
rect -330 12545 0 12555
rect -314 12485 -56 12545
rect -4 12485 0 12545
rect -330 12285 0 12485
rect -314 12225 -56 12285
rect -4 12225 0 12285
rect -330 12215 0 12225
rect 30 12545 400 12555
rect 30 12485 34 12545
rect 86 12485 344 12545
rect 396 12485 400 12545
rect 30 12410 400 12485
rect 430 12545 800 12555
rect 430 12485 434 12545
rect 486 12485 744 12545
rect 796 12485 800 12545
rect 430 12410 800 12485
rect 830 12545 1200 12555
rect 830 12485 834 12545
rect 886 12485 1144 12545
rect 1196 12485 1200 12545
rect 830 12410 1200 12485
rect 1230 12545 1600 12555
rect 1230 12485 1234 12545
rect 1286 12485 1544 12545
rect 1596 12485 1600 12545
rect 1230 12410 1600 12485
rect 1630 12545 2000 12555
rect 1630 12485 1634 12545
rect 1686 12485 1944 12545
rect 1996 12485 2000 12545
rect 1630 12410 2000 12485
rect 2030 12545 2400 12555
rect 2030 12485 2034 12545
rect 2086 12485 2344 12545
rect 2396 12485 2400 12545
rect 2030 12410 2400 12485
rect 2430 12545 2800 12555
rect 2430 12485 2434 12545
rect 2486 12485 2744 12545
rect 2796 12485 2800 12545
rect 2430 12410 2800 12485
rect 30 12370 2800 12410
rect 30 12285 400 12370
rect 30 12225 34 12285
rect 86 12225 344 12285
rect 396 12225 400 12285
rect 30 12215 400 12225
rect 430 12285 800 12370
rect 430 12225 434 12285
rect 486 12225 744 12285
rect 796 12225 800 12285
rect 430 12215 800 12225
rect 830 12285 1200 12370
rect 830 12225 834 12285
rect 886 12225 1144 12285
rect 1196 12225 1200 12285
rect 830 12215 1200 12225
rect 1230 12285 1600 12370
rect 1230 12225 1234 12285
rect 1286 12225 1544 12285
rect 1596 12225 1600 12285
rect 1230 12215 1600 12225
rect 1630 12285 2000 12370
rect 1630 12225 1634 12285
rect 1686 12225 1944 12285
rect 1996 12225 2000 12285
rect 1630 12215 2000 12225
rect 2030 12285 2400 12370
rect 2030 12225 2034 12285
rect 2086 12225 2344 12285
rect 2396 12225 2400 12285
rect 2030 12215 2400 12225
rect 2430 12285 2800 12370
rect 2430 12225 2434 12285
rect 2486 12225 2744 12285
rect 2796 12225 2800 12285
rect 2430 12215 2800 12225
rect 2830 12545 3200 12555
rect 2830 12485 2834 12545
rect 2886 12485 3144 12545
rect 3196 12485 3200 12545
rect 2830 12410 3200 12485
rect 3230 12545 3600 12555
rect 3230 12485 3234 12545
rect 3286 12485 3544 12545
rect 3596 12485 3600 12545
rect 3230 12410 3600 12485
rect 3630 12545 4000 12555
rect 3630 12485 3634 12545
rect 3686 12485 3944 12545
rect 3996 12485 4000 12545
rect 3630 12410 4000 12485
rect 4030 12545 4400 12555
rect 4030 12485 4034 12545
rect 4086 12485 4344 12545
rect 4396 12485 4400 12545
rect 4030 12410 4400 12485
rect 4430 12545 4800 12555
rect 4430 12485 4434 12545
rect 4486 12485 4744 12545
rect 4796 12485 4800 12545
rect 4430 12410 4800 12485
rect 4830 12545 5200 12555
rect 4830 12485 4834 12545
rect 4886 12485 5144 12545
rect 5196 12485 5200 12545
rect 4830 12410 5200 12485
rect 5230 12545 5600 12555
rect 5230 12485 5234 12545
rect 5286 12485 5544 12545
rect 5596 12485 5600 12545
rect 5230 12410 5600 12485
rect 5630 12545 6000 12555
rect 5630 12485 5634 12545
rect 5686 12485 5944 12545
rect 5996 12485 6000 12545
rect 5630 12410 6000 12485
rect 2830 12370 6000 12410
rect 2830 12285 3200 12370
rect 2830 12225 2834 12285
rect 2886 12225 3144 12285
rect 3196 12225 3200 12285
rect 2830 12215 3200 12225
rect 3230 12285 3600 12370
rect 3230 12225 3234 12285
rect 3286 12225 3544 12285
rect 3596 12225 3600 12285
rect 3230 12215 3600 12225
rect 3630 12285 4000 12370
rect 3630 12225 3634 12285
rect 3686 12225 3944 12285
rect 3996 12225 4000 12285
rect 3630 12215 4000 12225
rect 4030 12285 4400 12370
rect 4030 12225 4034 12285
rect 4086 12225 4344 12285
rect 4396 12225 4400 12285
rect 4030 12215 4400 12225
rect 4430 12285 4800 12370
rect 4430 12225 4434 12285
rect 4486 12225 4744 12285
rect 4796 12225 4800 12285
rect 4430 12215 4800 12225
rect 4830 12285 5200 12370
rect 4830 12225 4834 12285
rect 4886 12225 5144 12285
rect 5196 12225 5200 12285
rect 4830 12215 5200 12225
rect 5230 12285 5600 12370
rect 5230 12225 5234 12285
rect 5286 12225 5544 12285
rect 5596 12225 5600 12285
rect 5230 12215 5600 12225
rect 5630 12285 6000 12370
rect 5630 12225 5634 12285
rect 5686 12225 5944 12285
rect 5996 12225 6000 12285
rect 5630 12215 6000 12225
rect 6030 12545 6400 12555
rect 6030 12485 6034 12545
rect 6086 12485 6344 12545
rect 6396 12485 6400 12545
rect 6030 12410 6400 12485
rect 6430 12545 6800 12555
rect 6430 12485 6434 12545
rect 6486 12485 6744 12545
rect 6796 12485 6800 12545
rect 6430 12410 6800 12485
rect 6830 12545 7200 12555
rect 6830 12485 6834 12545
rect 6886 12485 7144 12545
rect 7196 12485 7200 12545
rect 6830 12410 7200 12485
rect 7230 12545 7600 12555
rect 7230 12485 7234 12545
rect 7286 12485 7544 12545
rect 7596 12485 7600 12545
rect 7230 12410 7600 12485
rect 6030 12370 7600 12410
rect 6030 12285 6400 12370
rect 6030 12225 6034 12285
rect 6086 12225 6344 12285
rect 6396 12225 6400 12285
rect 6030 12215 6400 12225
rect 6430 12285 6800 12370
rect 6430 12225 6434 12285
rect 6486 12225 6744 12285
rect 6796 12225 6800 12285
rect 6430 12215 6800 12225
rect 6830 12285 7200 12370
rect 6830 12225 6834 12285
rect 6886 12225 7144 12285
rect 7196 12225 7200 12285
rect 6830 12215 7200 12225
rect 7230 12285 7600 12370
rect 7230 12225 7234 12285
rect 7286 12225 7544 12285
rect 7596 12225 7600 12285
rect 7230 12215 7600 12225
rect 7630 12545 8000 12555
rect 7630 12485 7634 12545
rect 7686 12485 7944 12545
rect 7996 12485 8000 12545
rect 7630 12410 8000 12485
rect 8030 12545 8400 12555
rect 8030 12485 8034 12545
rect 8086 12485 8344 12545
rect 8396 12485 8400 12545
rect 8030 12410 8400 12485
rect 7630 12370 8400 12410
rect 7630 12285 8000 12370
rect 7630 12225 7634 12285
rect 7686 12225 7944 12285
rect 7996 12225 8000 12285
rect 7630 12215 8000 12225
rect 8030 12285 8400 12370
rect 8030 12225 8034 12285
rect 8086 12225 8344 12285
rect 8396 12225 8400 12285
rect 8030 12215 8400 12225
rect 8430 12545 8800 12555
rect 8430 12485 8434 12545
rect 8486 12485 8744 12545
rect 8796 12485 8800 12545
rect 8430 12285 8800 12485
rect 8430 12225 8434 12285
rect 8486 12225 8744 12285
rect 8796 12225 8800 12285
rect 8430 12215 8800 12225
rect 8830 12545 9200 12555
rect 8830 12485 8834 12545
rect 8886 12485 9144 12545
rect 9196 12485 9200 12545
rect 8830 12285 9200 12485
rect 8830 12225 8834 12285
rect 8886 12225 9144 12285
rect 9196 12225 9200 12285
rect 8830 12215 9200 12225
rect 9230 12545 9600 12555
rect 9230 12485 9234 12545
rect 9286 12485 9544 12545
rect 9596 12485 9600 12545
rect 9230 12410 9600 12485
rect 9630 12545 10000 12555
rect 9630 12485 9634 12545
rect 9686 12485 9944 12545
rect 9996 12485 10000 12545
rect 9630 12410 10000 12485
rect 9230 12370 10000 12410
rect 9230 12285 9600 12370
rect 9230 12225 9234 12285
rect 9286 12225 9544 12285
rect 9596 12225 9600 12285
rect 9230 12215 9600 12225
rect 9630 12285 10000 12370
rect 9630 12225 9634 12285
rect 9686 12225 9944 12285
rect 9996 12225 10000 12285
rect 9630 12215 10000 12225
rect 10030 12545 10400 12555
rect 10030 12485 10034 12545
rect 10086 12485 10344 12545
rect 10396 12485 10400 12545
rect 10030 12410 10400 12485
rect 10430 12545 10800 12555
rect 10430 12485 10434 12545
rect 10486 12485 10744 12545
rect 10796 12485 10800 12545
rect 10430 12410 10800 12485
rect 10830 12545 11200 12555
rect 10830 12485 10834 12545
rect 10886 12485 11144 12545
rect 11196 12485 11200 12545
rect 10830 12410 11200 12485
rect 10030 12370 11200 12410
rect 10030 12285 10400 12370
rect 10030 12225 10034 12285
rect 10086 12225 10344 12285
rect 10396 12225 10400 12285
rect 10030 12215 10400 12225
rect 10430 12285 10800 12370
rect 10430 12225 10434 12285
rect 10486 12225 10744 12285
rect 10796 12225 10800 12285
rect 10430 12215 10800 12225
rect 10830 12285 11200 12370
rect 10830 12225 10834 12285
rect 10886 12225 11144 12285
rect 11196 12225 11200 12285
rect 10830 12215 11200 12225
rect 11230 12545 11600 12555
rect 11230 12485 11234 12545
rect 11286 12485 11544 12545
rect 11596 12485 11600 12545
rect 11230 12285 11600 12485
rect 11230 12225 11234 12285
rect 11286 12225 11544 12285
rect 11596 12225 11600 12285
rect 11230 12215 11600 12225
rect 11630 12545 12000 12555
rect 11630 12485 11634 12545
rect 11686 12485 11944 12545
rect 11996 12485 12000 12545
rect 11630 12285 12000 12485
rect 11630 12225 11634 12285
rect 11686 12225 11944 12285
rect 11996 12225 12000 12285
rect 11630 12215 12000 12225
rect 12030 12545 12400 12555
rect 12030 12485 12034 12545
rect 12086 12485 12344 12545
rect 12396 12485 12400 12545
rect 12030 12410 12400 12485
rect 12430 12545 12800 12555
rect 12430 12485 12434 12545
rect 12486 12485 12744 12545
rect 12796 12485 12800 12545
rect 12430 12410 12800 12485
rect 12830 12545 13200 12555
rect 12830 12485 12834 12545
rect 12886 12485 13144 12545
rect 13196 12485 13200 12545
rect 12830 12410 13200 12485
rect 12030 12370 13390 12410
rect 12030 12285 12400 12370
rect 12030 12225 12034 12285
rect 12086 12225 12344 12285
rect 12396 12225 12400 12285
rect 12030 12215 12400 12225
rect 12430 12285 12800 12370
rect 12430 12225 12434 12285
rect 12486 12225 12744 12285
rect 12796 12225 12800 12285
rect 12430 12215 12800 12225
rect 12830 12285 13200 12370
rect 12830 12225 12834 12285
rect 12886 12225 13144 12285
rect 13196 12225 13200 12285
rect 12830 12215 13200 12225
rect -330 12185 -324 12215
rect 30 12185 70 12215
rect 430 12185 470 12215
rect 830 12185 870 12215
rect 1230 12185 1270 12215
rect 1630 12185 1670 12215
rect 2030 12185 2070 12215
rect 2430 12185 2470 12215
rect 2830 12185 2870 12215
rect 3230 12185 3270 12215
rect 3630 12185 3670 12215
rect 4030 12185 4070 12215
rect 4430 12185 4470 12215
rect 4830 12185 4870 12215
rect 5230 12185 5270 12215
rect 6030 12185 6070 12215
rect 6430 12185 6470 12215
rect 6830 12185 6870 12215
rect 7230 12185 7270 12215
rect 7630 12185 7670 12215
rect 8030 12185 8070 12215
rect 8430 12185 8470 12215
rect 9230 12185 9270 12215
rect 9630 12185 9670 12215
rect 10030 12185 10070 12215
rect 10430 12185 10470 12215
rect 10830 12185 10870 12215
rect 11230 12185 11270 12215
rect 11630 12185 11670 12215
rect -330 12175 0 12185
rect -314 12115 -56 12175
rect -4 12115 0 12175
rect -330 11915 0 12115
rect -314 11855 -56 11915
rect -4 11855 0 11915
rect -330 11845 0 11855
rect 30 12175 400 12185
rect 30 12115 34 12175
rect 86 12115 344 12175
rect 396 12115 400 12175
rect 30 12040 400 12115
rect 430 12175 800 12185
rect 430 12115 434 12175
rect 486 12115 744 12175
rect 796 12115 800 12175
rect 430 12040 800 12115
rect 830 12175 1200 12185
rect 830 12115 834 12175
rect 886 12115 1144 12175
rect 1196 12115 1200 12175
rect 830 12040 1200 12115
rect 1230 12175 1600 12185
rect 1230 12115 1234 12175
rect 1286 12115 1544 12175
rect 1596 12115 1600 12175
rect 1230 12040 1600 12115
rect 1630 12175 2000 12185
rect 1630 12115 1634 12175
rect 1686 12115 1944 12175
rect 1996 12115 2000 12175
rect 1630 12040 2000 12115
rect 2030 12175 2400 12185
rect 2030 12115 2034 12175
rect 2086 12115 2344 12175
rect 2396 12115 2400 12175
rect 2030 12040 2400 12115
rect 2430 12175 2800 12185
rect 2430 12115 2434 12175
rect 2486 12115 2744 12175
rect 2796 12115 2800 12175
rect 2430 12040 2800 12115
rect 30 12000 2800 12040
rect 30 11915 400 12000
rect 30 11855 34 11915
rect 86 11855 344 11915
rect 396 11855 400 11915
rect 30 11845 400 11855
rect 430 11915 800 12000
rect 430 11855 434 11915
rect 486 11855 744 11915
rect 796 11855 800 11915
rect 430 11845 800 11855
rect 830 11915 1200 12000
rect 830 11855 834 11915
rect 886 11855 1144 11915
rect 1196 11855 1200 11915
rect 830 11845 1200 11855
rect 1230 11915 1600 12000
rect 1230 11855 1234 11915
rect 1286 11855 1544 11915
rect 1596 11855 1600 11915
rect 1230 11845 1600 11855
rect 1630 11915 2000 12000
rect 1630 11855 1634 11915
rect 1686 11855 1944 11915
rect 1996 11855 2000 11915
rect 1630 11845 2000 11855
rect 2030 11915 2400 12000
rect 2030 11855 2034 11915
rect 2086 11855 2344 11915
rect 2396 11855 2400 11915
rect 2030 11845 2400 11855
rect 2430 11915 2800 12000
rect 2430 11855 2434 11915
rect 2486 11855 2744 11915
rect 2796 11855 2800 11915
rect 2430 11845 2800 11855
rect 2830 12175 3200 12185
rect 2830 12115 2834 12175
rect 2886 12115 3144 12175
rect 3196 12115 3200 12175
rect 2830 12040 3200 12115
rect 3230 12175 3600 12185
rect 3230 12115 3234 12175
rect 3286 12115 3544 12175
rect 3596 12115 3600 12175
rect 3230 12040 3600 12115
rect 3630 12175 4000 12185
rect 3630 12115 3634 12175
rect 3686 12115 3944 12175
rect 3996 12115 4000 12175
rect 3630 12040 4000 12115
rect 4030 12175 4400 12185
rect 4030 12115 4034 12175
rect 4086 12115 4344 12175
rect 4396 12115 4400 12175
rect 4030 12040 4400 12115
rect 4430 12175 4800 12185
rect 4430 12115 4434 12175
rect 4486 12115 4744 12175
rect 4796 12115 4800 12175
rect 4430 12040 4800 12115
rect 4830 12175 5200 12185
rect 4830 12115 4834 12175
rect 4886 12115 5144 12175
rect 5196 12115 5200 12175
rect 4830 12040 5200 12115
rect 5230 12175 5600 12185
rect 5230 12115 5234 12175
rect 5286 12115 5544 12175
rect 5596 12115 5600 12175
rect 5230 12040 5600 12115
rect 2830 12000 5600 12040
rect 2830 11915 3200 12000
rect 2830 11855 2834 11915
rect 2886 11855 3144 11915
rect 3196 11855 3200 11915
rect 2830 11845 3200 11855
rect 3230 11915 3600 12000
rect 3230 11855 3234 11915
rect 3286 11855 3544 11915
rect 3596 11855 3600 11915
rect 3230 11845 3600 11855
rect 3630 11915 4000 12000
rect 3630 11855 3634 11915
rect 3686 11855 3944 11915
rect 3996 11855 4000 11915
rect 3630 11845 4000 11855
rect 4030 11915 4400 12000
rect 4030 11855 4034 11915
rect 4086 11855 4344 11915
rect 4396 11855 4400 11915
rect 4030 11845 4400 11855
rect 4430 11915 4800 12000
rect 4430 11855 4434 11915
rect 4486 11855 4744 11915
rect 4796 11855 4800 11915
rect 4430 11845 4800 11855
rect 4830 11915 5200 12000
rect 4830 11855 4834 11915
rect 4886 11855 5144 11915
rect 5196 11855 5200 11915
rect 4830 11845 5200 11855
rect 5230 11915 5600 12000
rect 5230 11855 5234 11915
rect 5286 11855 5544 11915
rect 5596 11855 5600 11915
rect 5230 11845 5600 11855
rect 5630 12175 6000 12185
rect 5630 12115 5634 12175
rect 5686 12115 5944 12175
rect 5996 12115 6000 12175
rect 5630 12040 6000 12115
rect 6030 12175 6400 12185
rect 6030 12115 6034 12175
rect 6086 12115 6344 12175
rect 6396 12115 6400 12175
rect 6030 12040 6400 12115
rect 6430 12175 6800 12185
rect 6430 12115 6434 12175
rect 6486 12115 6744 12175
rect 6796 12115 6800 12175
rect 6430 12040 6800 12115
rect 6830 12175 7200 12185
rect 6830 12115 6834 12175
rect 6886 12115 7144 12175
rect 7196 12115 7200 12175
rect 6830 12040 7200 12115
rect 7230 12175 7600 12185
rect 7230 12115 7234 12175
rect 7286 12115 7544 12175
rect 7596 12115 7600 12175
rect 7230 12040 7600 12115
rect 5630 12000 7600 12040
rect 5630 11915 6000 12000
rect 5630 11855 5634 11915
rect 5686 11855 5944 11915
rect 5996 11855 6000 11915
rect 5630 11845 6000 11855
rect 6030 11915 6400 12000
rect 6030 11855 6034 11915
rect 6086 11855 6344 11915
rect 6396 11855 6400 11915
rect 6030 11845 6400 11855
rect 6430 11915 6800 12000
rect 6430 11855 6434 11915
rect 6486 11855 6744 11915
rect 6796 11855 6800 11915
rect 6430 11845 6800 11855
rect 6830 11915 7200 12000
rect 6830 11855 6834 11915
rect 6886 11855 7144 11915
rect 7196 11855 7200 11915
rect 6830 11845 7200 11855
rect 7230 11915 7600 12000
rect 7230 11855 7234 11915
rect 7286 11855 7544 11915
rect 7596 11855 7600 11915
rect 7230 11845 7600 11855
rect 7630 12175 8000 12185
rect 7630 12115 7634 12175
rect 7686 12115 7944 12175
rect 7996 12115 8000 12175
rect 7630 12040 8000 12115
rect 8030 12175 8400 12185
rect 8030 12115 8034 12175
rect 8086 12115 8344 12175
rect 8396 12115 8400 12175
rect 8030 12040 8400 12115
rect 7630 12000 8400 12040
rect 7630 11915 8000 12000
rect 7630 11855 7634 11915
rect 7686 11855 7944 11915
rect 7996 11855 8000 11915
rect 7630 11845 8000 11855
rect 8030 11915 8400 12000
rect 8030 11855 8034 11915
rect 8086 11855 8344 11915
rect 8396 11855 8400 11915
rect 8030 11845 8400 11855
rect 8430 12175 8800 12185
rect 8430 12115 8434 12175
rect 8486 12115 8744 12175
rect 8796 12115 8800 12175
rect 8430 11915 8800 12115
rect 8430 11855 8434 11915
rect 8486 11855 8744 11915
rect 8796 11855 8800 11915
rect 8430 11845 8800 11855
rect 8830 12175 9200 12185
rect 8830 12115 8834 12175
rect 8886 12115 9144 12175
rect 9196 12115 9200 12175
rect 8830 12040 9200 12115
rect 9230 12175 9600 12185
rect 9230 12115 9234 12175
rect 9286 12115 9544 12175
rect 9596 12115 9600 12175
rect 9230 12040 9600 12115
rect 9630 12175 10000 12185
rect 9630 12115 9634 12175
rect 9686 12115 9944 12175
rect 9996 12115 10000 12175
rect 9630 12040 10000 12115
rect 8830 12000 10000 12040
rect 8830 11915 9200 12000
rect 8830 11855 8834 11915
rect 8886 11855 9144 11915
rect 9196 11855 9200 11915
rect 8830 11845 9200 11855
rect 9230 11915 9600 12000
rect 9230 11855 9234 11915
rect 9286 11855 9544 11915
rect 9596 11855 9600 11915
rect 9230 11845 9600 11855
rect 9630 11915 10000 12000
rect 9630 11855 9634 11915
rect 9686 11855 9944 11915
rect 9996 11855 10000 11915
rect 9630 11845 10000 11855
rect 10030 12175 10400 12185
rect 10030 12115 10034 12175
rect 10086 12115 10344 12175
rect 10396 12115 10400 12175
rect 10030 12040 10400 12115
rect 10430 12175 10800 12185
rect 10430 12115 10434 12175
rect 10486 12115 10744 12175
rect 10796 12115 10800 12175
rect 10430 12040 10800 12115
rect 10830 12175 11200 12185
rect 10830 12115 10834 12175
rect 10886 12115 11144 12175
rect 11196 12115 11200 12175
rect 10830 12040 11200 12115
rect 10030 12000 11200 12040
rect 10030 11915 10400 12000
rect 10030 11855 10034 11915
rect 10086 11855 10344 11915
rect 10396 11855 10400 11915
rect 10030 11845 10400 11855
rect 10430 11915 10800 12000
rect 10430 11855 10434 11915
rect 10486 11855 10744 11915
rect 10796 11855 10800 11915
rect 10430 11845 10800 11855
rect 10830 11915 11200 12000
rect 10830 11855 10834 11915
rect 10886 11855 11144 11915
rect 11196 11855 11200 11915
rect 10830 11845 11200 11855
rect 11230 12175 11600 12185
rect 11230 12115 11234 12175
rect 11286 12115 11544 12175
rect 11596 12115 11600 12175
rect 11230 11915 11600 12115
rect 11230 11855 11234 11915
rect 11286 11855 11544 11915
rect 11596 11855 11600 11915
rect 11230 11845 11600 11855
rect 11630 12175 12000 12185
rect 11630 12115 11634 12175
rect 11686 12115 11944 12175
rect 11996 12115 12000 12175
rect 11630 11915 12000 12115
rect 11630 11855 11634 11915
rect 11686 11855 11944 11915
rect 11996 11855 12000 11915
rect 11630 11845 12000 11855
rect 12030 12175 12400 12185
rect 12030 12115 12034 12175
rect 12086 12115 12344 12175
rect 12396 12115 12400 12175
rect 12030 11915 12400 12115
rect 12030 11855 12034 11915
rect 12086 11855 12344 11915
rect 12396 11855 12400 11915
rect 12030 11845 12400 11855
rect 12430 12175 12800 12185
rect 12430 12115 12434 12175
rect 12486 12115 12744 12175
rect 12796 12115 12800 12175
rect 12430 12040 12800 12115
rect 12830 12175 13200 12185
rect 12830 12115 12834 12175
rect 12886 12115 13144 12175
rect 13196 12115 13200 12175
rect 12830 12040 13200 12115
rect 12430 12000 13390 12040
rect 12430 11915 12800 12000
rect 12430 11855 12434 11915
rect 12486 11855 12744 11915
rect 12796 11855 12800 11915
rect 12430 11845 12800 11855
rect 12830 11915 13200 12000
rect 12830 11855 12834 11915
rect 12886 11855 13144 11915
rect 13196 11855 13200 11915
rect 12830 11845 13200 11855
rect -330 11815 -324 11845
rect 30 11815 70 11845
rect 430 11815 470 11845
rect 830 11815 870 11845
rect 1230 11815 1270 11845
rect 1630 11815 1670 11845
rect 2030 11815 2070 11845
rect 2430 11815 2470 11845
rect 2830 11815 2870 11845
rect 3230 11815 3270 11845
rect 3630 11815 3670 11845
rect 4030 11815 4070 11845
rect 4430 11815 4470 11845
rect 4830 11815 4870 11845
rect 5230 11815 5270 11845
rect 5630 11815 5670 11845
rect 6030 11815 6070 11845
rect 6430 11815 6470 11845
rect 6830 11815 6870 11845
rect 7230 11815 7270 11845
rect 7630 11815 7670 11845
rect 8030 11815 8070 11845
rect 8430 11815 8470 11845
rect 8830 11815 8870 11845
rect 9230 11815 9270 11845
rect 9630 11815 9670 11845
rect 10030 11815 10070 11845
rect 10430 11815 10470 11845
rect 10830 11815 10870 11845
rect 11230 11815 11270 11845
rect 11630 11815 11670 11845
rect 12030 11815 12070 11845
rect -330 11805 0 11815
rect -314 11745 -56 11805
rect -4 11745 0 11805
rect -330 11545 0 11745
rect -314 11485 -56 11545
rect -4 11485 0 11545
rect -330 11475 0 11485
rect 30 11805 400 11815
rect 30 11745 34 11805
rect 86 11745 344 11805
rect 396 11745 400 11805
rect 30 11670 400 11745
rect 430 11805 800 11815
rect 430 11745 434 11805
rect 486 11745 744 11805
rect 796 11745 800 11805
rect 430 11670 800 11745
rect 830 11805 1200 11815
rect 830 11745 834 11805
rect 886 11745 1144 11805
rect 1196 11745 1200 11805
rect 830 11670 1200 11745
rect 1230 11805 1600 11815
rect 1230 11745 1234 11805
rect 1286 11745 1544 11805
rect 1596 11745 1600 11805
rect 1230 11670 1600 11745
rect 1630 11805 2000 11815
rect 1630 11745 1634 11805
rect 1686 11745 1944 11805
rect 1996 11745 2000 11805
rect 1630 11670 2000 11745
rect 2030 11805 2400 11815
rect 2030 11745 2034 11805
rect 2086 11745 2344 11805
rect 2396 11745 2400 11805
rect 2030 11670 2400 11745
rect 2430 11805 2800 11815
rect 2430 11745 2434 11805
rect 2486 11745 2744 11805
rect 2796 11745 2800 11805
rect 2430 11670 2800 11745
rect 30 11630 2800 11670
rect 30 11545 400 11630
rect 30 11485 34 11545
rect 86 11485 344 11545
rect 396 11485 400 11545
rect 30 11475 400 11485
rect 430 11545 800 11630
rect 430 11485 434 11545
rect 486 11485 744 11545
rect 796 11485 800 11545
rect 430 11475 800 11485
rect 830 11545 1200 11630
rect 830 11485 834 11545
rect 886 11485 1144 11545
rect 1196 11485 1200 11545
rect 830 11475 1200 11485
rect 1230 11545 1600 11630
rect 1230 11485 1234 11545
rect 1286 11485 1544 11545
rect 1596 11485 1600 11545
rect 1230 11475 1600 11485
rect 1630 11545 2000 11630
rect 1630 11485 1634 11545
rect 1686 11485 1944 11545
rect 1996 11485 2000 11545
rect 1630 11475 2000 11485
rect 2030 11545 2400 11630
rect 2030 11485 2034 11545
rect 2086 11485 2344 11545
rect 2396 11485 2400 11545
rect 2030 11475 2400 11485
rect 2430 11545 2800 11630
rect 2430 11485 2434 11545
rect 2486 11485 2744 11545
rect 2796 11485 2800 11545
rect 2430 11475 2800 11485
rect 2830 11805 3200 11815
rect 2830 11745 2834 11805
rect 2886 11745 3144 11805
rect 3196 11745 3200 11805
rect 2830 11670 3200 11745
rect 3230 11805 3600 11815
rect 3230 11745 3234 11805
rect 3286 11745 3544 11805
rect 3596 11745 3600 11805
rect 3230 11670 3600 11745
rect 3630 11805 4000 11815
rect 3630 11745 3634 11805
rect 3686 11745 3944 11805
rect 3996 11745 4000 11805
rect 3630 11670 4000 11745
rect 4030 11805 4400 11815
rect 4030 11745 4034 11805
rect 4086 11745 4344 11805
rect 4396 11745 4400 11805
rect 4030 11670 4400 11745
rect 4430 11805 4800 11815
rect 4430 11745 4434 11805
rect 4486 11745 4744 11805
rect 4796 11745 4800 11805
rect 4430 11670 4800 11745
rect 4830 11805 5200 11815
rect 4830 11745 4834 11805
rect 4886 11745 5144 11805
rect 5196 11745 5200 11805
rect 4830 11670 5200 11745
rect 5230 11805 5600 11815
rect 5230 11745 5234 11805
rect 5286 11745 5544 11805
rect 5596 11745 5600 11805
rect 5230 11670 5600 11745
rect 2830 11630 5600 11670
rect 2830 11545 3200 11630
rect 2830 11485 2834 11545
rect 2886 11485 3144 11545
rect 3196 11485 3200 11545
rect 2830 11475 3200 11485
rect 3230 11545 3600 11630
rect 3230 11485 3234 11545
rect 3286 11485 3544 11545
rect 3596 11485 3600 11545
rect 3230 11475 3600 11485
rect 3630 11545 4000 11630
rect 3630 11485 3634 11545
rect 3686 11485 3944 11545
rect 3996 11485 4000 11545
rect 3630 11475 4000 11485
rect 4030 11545 4400 11630
rect 4030 11485 4034 11545
rect 4086 11485 4344 11545
rect 4396 11485 4400 11545
rect 4030 11475 4400 11485
rect 4430 11545 4800 11630
rect 4430 11485 4434 11545
rect 4486 11485 4744 11545
rect 4796 11485 4800 11545
rect 4430 11475 4800 11485
rect 4830 11545 5200 11630
rect 4830 11485 4834 11545
rect 4886 11485 5144 11545
rect 5196 11485 5200 11545
rect 4830 11475 5200 11485
rect 5230 11545 5600 11630
rect 5230 11485 5234 11545
rect 5286 11485 5544 11545
rect 5596 11485 5600 11545
rect 5230 11475 5600 11485
rect 5630 11805 6000 11815
rect 5630 11745 5634 11805
rect 5686 11745 5944 11805
rect 5996 11745 6000 11805
rect 5630 11670 6000 11745
rect 6030 11805 6400 11815
rect 6030 11745 6034 11805
rect 6086 11745 6344 11805
rect 6396 11745 6400 11805
rect 6030 11670 6400 11745
rect 6430 11805 6800 11815
rect 6430 11745 6434 11805
rect 6486 11745 6744 11805
rect 6796 11745 6800 11805
rect 6430 11670 6800 11745
rect 6830 11805 7200 11815
rect 6830 11745 6834 11805
rect 6886 11745 7144 11805
rect 7196 11745 7200 11805
rect 6830 11670 7200 11745
rect 7230 11805 7600 11815
rect 7230 11745 7234 11805
rect 7286 11745 7544 11805
rect 7596 11745 7600 11805
rect 7230 11670 7600 11745
rect 5630 11630 7600 11670
rect 5630 11545 6000 11630
rect 5630 11485 5634 11545
rect 5686 11485 5944 11545
rect 5996 11485 6000 11545
rect 5630 11475 6000 11485
rect 6030 11545 6400 11630
rect 6030 11485 6034 11545
rect 6086 11485 6344 11545
rect 6396 11485 6400 11545
rect 6030 11475 6400 11485
rect 6430 11545 6800 11630
rect 6430 11485 6434 11545
rect 6486 11485 6744 11545
rect 6796 11485 6800 11545
rect 6430 11475 6800 11485
rect 6830 11545 7200 11630
rect 6830 11485 6834 11545
rect 6886 11485 7144 11545
rect 7196 11485 7200 11545
rect 6830 11475 7200 11485
rect 7230 11545 7600 11630
rect 7230 11485 7234 11545
rect 7286 11485 7544 11545
rect 7596 11485 7600 11545
rect 7230 11475 7600 11485
rect 7630 11805 8000 11815
rect 7630 11745 7634 11805
rect 7686 11745 7944 11805
rect 7996 11745 8000 11805
rect 7630 11670 8000 11745
rect 8030 11805 8400 11815
rect 8030 11745 8034 11805
rect 8086 11745 8344 11805
rect 8396 11745 8400 11805
rect 8030 11670 8400 11745
rect 7630 11630 8400 11670
rect 7630 11545 8000 11630
rect 7630 11485 7634 11545
rect 7686 11485 7944 11545
rect 7996 11485 8000 11545
rect 7630 11475 8000 11485
rect 8030 11545 8400 11630
rect 8030 11485 8034 11545
rect 8086 11485 8344 11545
rect 8396 11485 8400 11545
rect 8030 11475 8400 11485
rect 8430 11805 8800 11815
rect 8430 11745 8434 11805
rect 8486 11745 8744 11805
rect 8796 11745 8800 11805
rect 8430 11545 8800 11745
rect 8430 11485 8434 11545
rect 8486 11485 8744 11545
rect 8796 11485 8800 11545
rect 8430 11475 8800 11485
rect 8830 11805 9200 11815
rect 8830 11745 8834 11805
rect 8886 11745 9144 11805
rect 9196 11745 9200 11805
rect 8830 11670 9200 11745
rect 9230 11805 9600 11815
rect 9230 11745 9234 11805
rect 9286 11745 9544 11805
rect 9596 11745 9600 11805
rect 9230 11670 9600 11745
rect 9630 11805 10000 11815
rect 9630 11745 9634 11805
rect 9686 11745 9944 11805
rect 9996 11745 10000 11805
rect 9630 11670 10000 11745
rect 8830 11630 10000 11670
rect 8830 11545 9200 11630
rect 8830 11485 8834 11545
rect 8886 11485 9144 11545
rect 9196 11485 9200 11545
rect 8830 11475 9200 11485
rect 9230 11545 9600 11630
rect 9230 11485 9234 11545
rect 9286 11485 9544 11545
rect 9596 11485 9600 11545
rect 9230 11475 9600 11485
rect 9630 11545 10000 11630
rect 9630 11485 9634 11545
rect 9686 11485 9944 11545
rect 9996 11485 10000 11545
rect 9630 11475 10000 11485
rect 10030 11805 10400 11815
rect 10030 11745 10034 11805
rect 10086 11745 10344 11805
rect 10396 11745 10400 11805
rect 10030 11670 10400 11745
rect 10430 11805 10800 11815
rect 10430 11745 10434 11805
rect 10486 11745 10744 11805
rect 10796 11745 10800 11805
rect 10430 11670 10800 11745
rect 10830 11805 11200 11815
rect 10830 11745 10834 11805
rect 10886 11745 11144 11805
rect 11196 11745 11200 11805
rect 10830 11670 11200 11745
rect 10030 11630 11200 11670
rect 10030 11545 10400 11630
rect 10030 11485 10034 11545
rect 10086 11485 10344 11545
rect 10396 11485 10400 11545
rect 10030 11475 10400 11485
rect 10430 11545 10800 11630
rect 10430 11485 10434 11545
rect 10486 11485 10744 11545
rect 10796 11485 10800 11545
rect 10430 11475 10800 11485
rect 10830 11545 11200 11630
rect 10830 11485 10834 11545
rect 10886 11485 11144 11545
rect 11196 11485 11200 11545
rect 10830 11475 11200 11485
rect 11230 11805 11600 11815
rect 11230 11745 11234 11805
rect 11286 11745 11544 11805
rect 11596 11745 11600 11805
rect 11230 11545 11600 11745
rect 11230 11485 11234 11545
rect 11286 11485 11544 11545
rect 11596 11485 11600 11545
rect 11230 11475 11600 11485
rect 11630 11805 12000 11815
rect 11630 11745 11634 11805
rect 11686 11745 11944 11805
rect 11996 11745 12000 11805
rect 11630 11545 12000 11745
rect 11630 11485 11634 11545
rect 11686 11485 11944 11545
rect 11996 11485 12000 11545
rect 11630 11475 12000 11485
rect 12030 11805 12400 11815
rect 12030 11745 12034 11805
rect 12086 11745 12344 11805
rect 12396 11745 12400 11805
rect 12030 11545 12400 11745
rect 12030 11485 12034 11545
rect 12086 11485 12344 11545
rect 12396 11485 12400 11545
rect 12030 11475 12400 11485
rect 12430 11805 12800 11815
rect 12430 11745 12434 11805
rect 12486 11745 12744 11805
rect 12796 11745 12800 11805
rect 12430 11670 12800 11745
rect 12830 11805 13200 11815
rect 12830 11745 12834 11805
rect 12886 11745 13144 11805
rect 13196 11745 13200 11805
rect 12830 11670 13200 11745
rect 12430 11630 13390 11670
rect 12430 11545 12800 11630
rect 12430 11485 12434 11545
rect 12486 11485 12744 11545
rect 12796 11485 12800 11545
rect 12430 11475 12800 11485
rect 12830 11545 13200 11630
rect 12830 11485 12834 11545
rect 12886 11485 13144 11545
rect 13196 11485 13200 11545
rect 12830 11475 13200 11485
rect -330 11445 -324 11475
rect 30 11445 70 11475
rect 430 11445 470 11475
rect 830 11445 870 11475
rect 1230 11445 1270 11475
rect 1630 11445 1670 11475
rect 2030 11445 2070 11475
rect 2430 11445 2470 11475
rect 2830 11445 2870 11475
rect 3230 11445 3270 11475
rect 3630 11445 3670 11475
rect 4030 11445 4070 11475
rect 4430 11445 4470 11475
rect 4830 11445 4870 11475
rect 5230 11445 5270 11475
rect 6030 11445 6070 11475
rect 6430 11445 6470 11475
rect 6830 11445 6870 11475
rect 7230 11445 7270 11475
rect 7630 11445 7670 11475
rect 8030 11445 8070 11475
rect 8430 11445 8470 11475
rect 9230 11445 9270 11475
rect 9630 11445 9670 11475
rect 10030 11445 10070 11475
rect 10430 11445 10470 11475
rect 10830 11445 10870 11475
rect 11230 11445 11270 11475
rect 11630 11445 11670 11475
rect 12030 11445 12070 11475
rect -330 11435 0 11445
rect -314 11375 -56 11435
rect -4 11375 0 11435
rect -330 11175 0 11375
rect -314 11115 -56 11175
rect -4 11115 0 11175
rect -330 11105 0 11115
rect 30 11435 400 11445
rect 30 11375 34 11435
rect 86 11375 344 11435
rect 396 11375 400 11435
rect 30 11300 400 11375
rect 430 11435 800 11445
rect 430 11375 434 11435
rect 486 11375 744 11435
rect 796 11375 800 11435
rect 430 11300 800 11375
rect 830 11435 1200 11445
rect 830 11375 834 11435
rect 886 11375 1144 11435
rect 1196 11375 1200 11435
rect 830 11300 1200 11375
rect 1230 11435 1600 11445
rect 1230 11375 1234 11435
rect 1286 11375 1544 11435
rect 1596 11375 1600 11435
rect 1230 11300 1600 11375
rect 1630 11435 2000 11445
rect 1630 11375 1634 11435
rect 1686 11375 1944 11435
rect 1996 11375 2000 11435
rect 1630 11300 2000 11375
rect 2030 11435 2400 11445
rect 2030 11375 2034 11435
rect 2086 11375 2344 11435
rect 2396 11375 2400 11435
rect 2030 11300 2400 11375
rect 2430 11435 2800 11445
rect 2430 11375 2434 11435
rect 2486 11375 2744 11435
rect 2796 11375 2800 11435
rect 2430 11300 2800 11375
rect 30 11260 2800 11300
rect 30 11175 400 11260
rect 30 11115 34 11175
rect 86 11115 344 11175
rect 396 11115 400 11175
rect 30 11105 400 11115
rect 430 11175 800 11260
rect 430 11115 434 11175
rect 486 11115 744 11175
rect 796 11115 800 11175
rect 430 11105 800 11115
rect 830 11175 1200 11260
rect 830 11115 834 11175
rect 886 11115 1144 11175
rect 1196 11115 1200 11175
rect 830 11105 1200 11115
rect 1230 11175 1600 11260
rect 1230 11115 1234 11175
rect 1286 11115 1544 11175
rect 1596 11115 1600 11175
rect 1230 11105 1600 11115
rect 1630 11175 2000 11260
rect 1630 11115 1634 11175
rect 1686 11115 1944 11175
rect 1996 11115 2000 11175
rect 1630 11105 2000 11115
rect 2030 11175 2400 11260
rect 2030 11115 2034 11175
rect 2086 11115 2344 11175
rect 2396 11115 2400 11175
rect 2030 11105 2400 11115
rect 2430 11175 2800 11260
rect 2430 11115 2434 11175
rect 2486 11115 2744 11175
rect 2796 11115 2800 11175
rect 2430 11105 2800 11115
rect 2830 11435 3200 11445
rect 2830 11375 2834 11435
rect 2886 11375 3144 11435
rect 3196 11375 3200 11435
rect 2830 11300 3200 11375
rect 3230 11435 3600 11445
rect 3230 11375 3234 11435
rect 3286 11375 3544 11435
rect 3596 11375 3600 11435
rect 3230 11300 3600 11375
rect 3630 11435 4000 11445
rect 3630 11375 3634 11435
rect 3686 11375 3944 11435
rect 3996 11375 4000 11435
rect 3630 11300 4000 11375
rect 4030 11435 4400 11445
rect 4030 11375 4034 11435
rect 4086 11375 4344 11435
rect 4396 11375 4400 11435
rect 4030 11300 4400 11375
rect 4430 11435 4800 11445
rect 4430 11375 4434 11435
rect 4486 11375 4744 11435
rect 4796 11375 4800 11435
rect 4430 11300 4800 11375
rect 4830 11435 5200 11445
rect 4830 11375 4834 11435
rect 4886 11375 5144 11435
rect 5196 11375 5200 11435
rect 4830 11300 5200 11375
rect 5230 11435 5600 11445
rect 5230 11375 5234 11435
rect 5286 11375 5544 11435
rect 5596 11375 5600 11435
rect 5230 11300 5600 11375
rect 5630 11435 6000 11445
rect 5630 11375 5634 11435
rect 5686 11375 5944 11435
rect 5996 11375 6000 11435
rect 5630 11300 6000 11375
rect 2830 11260 6000 11300
rect 2830 11175 3200 11260
rect 2830 11115 2834 11175
rect 2886 11115 3144 11175
rect 3196 11115 3200 11175
rect 2830 11105 3200 11115
rect 3230 11175 3600 11260
rect 3230 11115 3234 11175
rect 3286 11115 3544 11175
rect 3596 11115 3600 11175
rect 3230 11105 3600 11115
rect 3630 11175 4000 11260
rect 3630 11115 3634 11175
rect 3686 11115 3944 11175
rect 3996 11115 4000 11175
rect 3630 11105 4000 11115
rect 4030 11175 4400 11260
rect 4030 11115 4034 11175
rect 4086 11115 4344 11175
rect 4396 11115 4400 11175
rect 4030 11105 4400 11115
rect 4430 11175 4800 11260
rect 4430 11115 4434 11175
rect 4486 11115 4744 11175
rect 4796 11115 4800 11175
rect 4430 11105 4800 11115
rect 4830 11175 5200 11260
rect 4830 11115 4834 11175
rect 4886 11115 5144 11175
rect 5196 11115 5200 11175
rect 4830 11105 5200 11115
rect 5230 11175 5600 11260
rect 5230 11115 5234 11175
rect 5286 11115 5544 11175
rect 5596 11115 5600 11175
rect 5230 11105 5600 11115
rect 5630 11175 6000 11260
rect 5630 11115 5634 11175
rect 5686 11115 5944 11175
rect 5996 11115 6000 11175
rect 5630 11105 6000 11115
rect 6030 11435 6400 11445
rect 6030 11375 6034 11435
rect 6086 11375 6344 11435
rect 6396 11375 6400 11435
rect 6030 11300 6400 11375
rect 6430 11435 6800 11445
rect 6430 11375 6434 11435
rect 6486 11375 6744 11435
rect 6796 11375 6800 11435
rect 6430 11300 6800 11375
rect 6830 11435 7200 11445
rect 6830 11375 6834 11435
rect 6886 11375 7144 11435
rect 7196 11375 7200 11435
rect 6830 11300 7200 11375
rect 7230 11435 7600 11445
rect 7230 11375 7234 11435
rect 7286 11375 7544 11435
rect 7596 11375 7600 11435
rect 7230 11300 7600 11375
rect 6030 11260 7600 11300
rect 6030 11175 6400 11260
rect 6030 11115 6034 11175
rect 6086 11115 6344 11175
rect 6396 11115 6400 11175
rect 6030 11105 6400 11115
rect 6430 11175 6800 11260
rect 6430 11115 6434 11175
rect 6486 11115 6744 11175
rect 6796 11115 6800 11175
rect 6430 11105 6800 11115
rect 6830 11175 7200 11260
rect 6830 11115 6834 11175
rect 6886 11115 7144 11175
rect 7196 11115 7200 11175
rect 6830 11105 7200 11115
rect 7230 11175 7600 11260
rect 7230 11115 7234 11175
rect 7286 11115 7544 11175
rect 7596 11115 7600 11175
rect 7230 11105 7600 11115
rect 7630 11435 8000 11445
rect 7630 11375 7634 11435
rect 7686 11375 7944 11435
rect 7996 11375 8000 11435
rect 7630 11300 8000 11375
rect 8030 11435 8400 11445
rect 8030 11375 8034 11435
rect 8086 11375 8344 11435
rect 8396 11375 8400 11435
rect 8030 11300 8400 11375
rect 7630 11260 8400 11300
rect 7630 11175 8000 11260
rect 7630 11115 7634 11175
rect 7686 11115 7944 11175
rect 7996 11115 8000 11175
rect 7630 11105 8000 11115
rect 8030 11175 8400 11260
rect 8030 11115 8034 11175
rect 8086 11115 8344 11175
rect 8396 11115 8400 11175
rect 8030 11105 8400 11115
rect 8430 11435 8800 11445
rect 8430 11375 8434 11435
rect 8486 11375 8744 11435
rect 8796 11375 8800 11435
rect 8430 11175 8800 11375
rect 8430 11115 8434 11175
rect 8486 11115 8744 11175
rect 8796 11115 8800 11175
rect 8430 11105 8800 11115
rect 8830 11435 9200 11445
rect 8830 11375 8834 11435
rect 8886 11375 9144 11435
rect 9196 11375 9200 11435
rect 8830 11175 9200 11375
rect 8830 11115 8834 11175
rect 8886 11115 9144 11175
rect 9196 11115 9200 11175
rect 8830 11105 9200 11115
rect 9230 11435 9600 11445
rect 9230 11375 9234 11435
rect 9286 11375 9544 11435
rect 9596 11375 9600 11435
rect 9230 11300 9600 11375
rect 9630 11435 10000 11445
rect 9630 11375 9634 11435
rect 9686 11375 9944 11435
rect 9996 11375 10000 11435
rect 9630 11300 10000 11375
rect 9230 11260 10000 11300
rect 9230 11175 9600 11260
rect 9230 11115 9234 11175
rect 9286 11115 9544 11175
rect 9596 11115 9600 11175
rect 9230 11105 9600 11115
rect 9630 11175 10000 11260
rect 9630 11115 9634 11175
rect 9686 11115 9944 11175
rect 9996 11115 10000 11175
rect 9630 11105 10000 11115
rect 10030 11435 10400 11445
rect 10030 11375 10034 11435
rect 10086 11375 10344 11435
rect 10396 11375 10400 11435
rect 10030 11300 10400 11375
rect 10430 11435 10800 11445
rect 10430 11375 10434 11435
rect 10486 11375 10744 11435
rect 10796 11375 10800 11435
rect 10430 11300 10800 11375
rect 10830 11435 11200 11445
rect 10830 11375 10834 11435
rect 10886 11375 11144 11435
rect 11196 11375 11200 11435
rect 10830 11300 11200 11375
rect 10030 11260 11200 11300
rect 10030 11175 10400 11260
rect 10030 11115 10034 11175
rect 10086 11115 10344 11175
rect 10396 11115 10400 11175
rect 10030 11105 10400 11115
rect 10430 11175 10800 11260
rect 10430 11115 10434 11175
rect 10486 11115 10744 11175
rect 10796 11115 10800 11175
rect 10430 11105 10800 11115
rect 10830 11175 11200 11260
rect 10830 11115 10834 11175
rect 10886 11115 11144 11175
rect 11196 11115 11200 11175
rect 10830 11105 11200 11115
rect 11230 11435 11600 11445
rect 11230 11375 11234 11435
rect 11286 11375 11544 11435
rect 11596 11375 11600 11435
rect 11230 11175 11600 11375
rect 11230 11115 11234 11175
rect 11286 11115 11544 11175
rect 11596 11115 11600 11175
rect 11230 11105 11600 11115
rect 11630 11435 12000 11445
rect 11630 11375 11634 11435
rect 11686 11375 11944 11435
rect 11996 11375 12000 11435
rect 11630 11175 12000 11375
rect 11630 11115 11634 11175
rect 11686 11115 11944 11175
rect 11996 11115 12000 11175
rect 11630 11105 12000 11115
rect 12030 11435 12400 11445
rect 12030 11375 12034 11435
rect 12086 11375 12344 11435
rect 12396 11375 12400 11435
rect 12030 11300 12400 11375
rect 12430 11435 12800 11445
rect 12430 11375 12434 11435
rect 12486 11375 12744 11435
rect 12796 11375 12800 11435
rect 12430 11300 12800 11375
rect 12830 11435 13200 11445
rect 12830 11375 12834 11435
rect 12886 11375 13144 11435
rect 13196 11375 13200 11435
rect 12830 11300 13200 11375
rect 12030 11260 13390 11300
rect 12030 11175 12400 11260
rect 12030 11115 12034 11175
rect 12086 11115 12344 11175
rect 12396 11115 12400 11175
rect 12030 11105 12400 11115
rect 12430 11175 12800 11260
rect 12430 11115 12434 11175
rect 12486 11115 12744 11175
rect 12796 11115 12800 11175
rect 12430 11105 12800 11115
rect 12830 11175 13200 11260
rect 12830 11115 12834 11175
rect 12886 11115 13144 11175
rect 13196 11115 13200 11175
rect 12830 11105 13200 11115
rect -330 11075 -324 11105
rect 30 11075 70 11105
rect 430 11075 470 11105
rect 830 11075 870 11105
rect 1230 11075 1270 11105
rect 1630 11075 1670 11105
rect 2030 11075 2070 11105
rect 2430 11075 2470 11105
rect 2830 11075 2870 11105
rect 3230 11075 3270 11105
rect 3630 11075 3670 11105
rect 4030 11075 4070 11105
rect 4430 11075 4470 11105
rect 4830 11075 4870 11105
rect 5230 11075 5270 11105
rect 5630 11075 5670 11105
rect 6030 11075 6070 11105
rect 6430 11075 6470 11105
rect 6830 11075 6870 11105
rect 7230 11075 7270 11105
rect 7630 11075 7670 11105
rect 8030 11075 8070 11105
rect 8430 11075 8470 11105
rect 8830 11075 8870 11105
rect 9230 11075 9270 11105
rect 9630 11075 9670 11105
rect 10430 11075 10470 11105
rect 10830 11075 10870 11105
rect 11230 11075 11270 11105
rect 11630 11075 11670 11105
rect -330 11065 0 11075
rect -314 11005 -56 11065
rect -4 11005 0 11065
rect -330 10805 0 11005
rect -314 10745 -56 10805
rect -4 10745 0 10805
rect -330 10735 0 10745
rect 30 11065 400 11075
rect 30 11005 34 11065
rect 86 11005 344 11065
rect 396 11005 400 11065
rect 30 10930 400 11005
rect 430 11065 800 11075
rect 430 11005 434 11065
rect 486 11005 744 11065
rect 796 11005 800 11065
rect 430 10930 800 11005
rect 830 11065 1200 11075
rect 830 11005 834 11065
rect 886 11005 1144 11065
rect 1196 11005 1200 11065
rect 830 10930 1200 11005
rect 1230 11065 1600 11075
rect 1230 11005 1234 11065
rect 1286 11005 1544 11065
rect 1596 11005 1600 11065
rect 1230 10930 1600 11005
rect 1630 11065 2000 11075
rect 1630 11005 1634 11065
rect 1686 11005 1944 11065
rect 1996 11005 2000 11065
rect 1630 10930 2000 11005
rect 2030 11065 2400 11075
rect 2030 11005 2034 11065
rect 2086 11005 2344 11065
rect 2396 11005 2400 11065
rect 2030 10930 2400 11005
rect 2430 11065 2800 11075
rect 2430 11005 2434 11065
rect 2486 11005 2744 11065
rect 2796 11005 2800 11065
rect 2430 10930 2800 11005
rect 30 10890 2800 10930
rect 30 10805 400 10890
rect 30 10745 34 10805
rect 86 10745 344 10805
rect 396 10745 400 10805
rect 30 10735 400 10745
rect 430 10805 800 10890
rect 430 10745 434 10805
rect 486 10745 744 10805
rect 796 10745 800 10805
rect 430 10735 800 10745
rect 830 10805 1200 10890
rect 830 10745 834 10805
rect 886 10745 1144 10805
rect 1196 10745 1200 10805
rect 830 10735 1200 10745
rect 1230 10805 1600 10890
rect 1230 10745 1234 10805
rect 1286 10745 1544 10805
rect 1596 10745 1600 10805
rect 1230 10735 1600 10745
rect 1630 10805 2000 10890
rect 1630 10745 1634 10805
rect 1686 10745 1944 10805
rect 1996 10745 2000 10805
rect 1630 10735 2000 10745
rect 2030 10805 2400 10890
rect 2030 10745 2034 10805
rect 2086 10745 2344 10805
rect 2396 10745 2400 10805
rect 2030 10735 2400 10745
rect 2430 10805 2800 10890
rect 2430 10745 2434 10805
rect 2486 10745 2744 10805
rect 2796 10745 2800 10805
rect 2430 10735 2800 10745
rect 2830 11065 3200 11075
rect 2830 11005 2834 11065
rect 2886 11005 3144 11065
rect 3196 11005 3200 11065
rect 2830 10930 3200 11005
rect 3230 11065 3600 11075
rect 3230 11005 3234 11065
rect 3286 11005 3544 11065
rect 3596 11005 3600 11065
rect 3230 10930 3600 11005
rect 3630 11065 4000 11075
rect 3630 11005 3634 11065
rect 3686 11005 3944 11065
rect 3996 11005 4000 11065
rect 3630 10930 4000 11005
rect 4030 11065 4400 11075
rect 4030 11005 4034 11065
rect 4086 11005 4344 11065
rect 4396 11005 4400 11065
rect 4030 10930 4400 11005
rect 4430 11065 4800 11075
rect 4430 11005 4434 11065
rect 4486 11005 4744 11065
rect 4796 11005 4800 11065
rect 4430 10930 4800 11005
rect 4830 11065 5200 11075
rect 4830 11005 4834 11065
rect 4886 11005 5144 11065
rect 5196 11005 5200 11065
rect 4830 10930 5200 11005
rect 5230 11065 5600 11075
rect 5230 11005 5234 11065
rect 5286 11005 5544 11065
rect 5596 11005 5600 11065
rect 5230 10930 5600 11005
rect 5630 11065 6000 11075
rect 5630 11005 5634 11065
rect 5686 11005 5944 11065
rect 5996 11005 6000 11065
rect 5630 10930 6000 11005
rect 2830 10890 6000 10930
rect 2830 10805 3200 10890
rect 2830 10745 2834 10805
rect 2886 10745 3144 10805
rect 3196 10745 3200 10805
rect 2830 10735 3200 10745
rect 3230 10805 3600 10890
rect 3230 10745 3234 10805
rect 3286 10745 3544 10805
rect 3596 10745 3600 10805
rect 3230 10735 3600 10745
rect 3630 10805 4000 10890
rect 3630 10745 3634 10805
rect 3686 10745 3944 10805
rect 3996 10745 4000 10805
rect 3630 10735 4000 10745
rect 4030 10805 4400 10890
rect 4030 10745 4034 10805
rect 4086 10745 4344 10805
rect 4396 10745 4400 10805
rect 4030 10735 4400 10745
rect 4430 10805 4800 10890
rect 4430 10745 4434 10805
rect 4486 10745 4744 10805
rect 4796 10745 4800 10805
rect 4430 10735 4800 10745
rect 4830 10805 5200 10890
rect 4830 10745 4834 10805
rect 4886 10745 5144 10805
rect 5196 10745 5200 10805
rect 4830 10735 5200 10745
rect 5230 10805 5600 10890
rect 5230 10745 5234 10805
rect 5286 10745 5544 10805
rect 5596 10745 5600 10805
rect 5230 10735 5600 10745
rect 5630 10805 6000 10890
rect 5630 10745 5634 10805
rect 5686 10745 5944 10805
rect 5996 10745 6000 10805
rect 5630 10735 6000 10745
rect 6030 11065 6400 11075
rect 6030 11005 6034 11065
rect 6086 11005 6344 11065
rect 6396 11005 6400 11065
rect 6030 10930 6400 11005
rect 6430 11065 6800 11075
rect 6430 11005 6434 11065
rect 6486 11005 6744 11065
rect 6796 11005 6800 11065
rect 6430 10930 6800 11005
rect 6830 11065 7200 11075
rect 6830 11005 6834 11065
rect 6886 11005 7144 11065
rect 7196 11005 7200 11065
rect 6830 10930 7200 11005
rect 7230 11065 7600 11075
rect 7230 11005 7234 11065
rect 7286 11005 7544 11065
rect 7596 11005 7600 11065
rect 7230 10930 7600 11005
rect 6030 10890 7600 10930
rect 6030 10805 6400 10890
rect 6030 10745 6034 10805
rect 6086 10745 6344 10805
rect 6396 10745 6400 10805
rect 6030 10735 6400 10745
rect 6430 10805 6800 10890
rect 6430 10745 6434 10805
rect 6486 10745 6744 10805
rect 6796 10745 6800 10805
rect 6430 10735 6800 10745
rect 6830 10805 7200 10890
rect 6830 10745 6834 10805
rect 6886 10745 7144 10805
rect 7196 10745 7200 10805
rect 6830 10735 7200 10745
rect 7230 10805 7600 10890
rect 7230 10745 7234 10805
rect 7286 10745 7544 10805
rect 7596 10745 7600 10805
rect 7230 10735 7600 10745
rect 7630 11065 8000 11075
rect 7630 11005 7634 11065
rect 7686 11005 7944 11065
rect 7996 11005 8000 11065
rect 7630 10930 8000 11005
rect 8030 11065 8400 11075
rect 8030 11005 8034 11065
rect 8086 11005 8344 11065
rect 8396 11005 8400 11065
rect 8030 10930 8400 11005
rect 7630 10890 8400 10930
rect 7630 10805 8000 10890
rect 7630 10745 7634 10805
rect 7686 10745 7944 10805
rect 7996 10745 8000 10805
rect 7630 10735 8000 10745
rect 8030 10805 8400 10890
rect 8030 10745 8034 10805
rect 8086 10745 8344 10805
rect 8396 10745 8400 10805
rect 8030 10735 8400 10745
rect 8430 11065 8800 11075
rect 8430 11005 8434 11065
rect 8486 11005 8744 11065
rect 8796 11005 8800 11065
rect 8430 10805 8800 11005
rect 8430 10745 8434 10805
rect 8486 10745 8744 10805
rect 8796 10745 8800 10805
rect 8430 10735 8800 10745
rect 8830 11065 9200 11075
rect 8830 11005 8834 11065
rect 8886 11005 9144 11065
rect 9196 11005 9200 11065
rect 8830 10805 9200 11005
rect 8830 10745 8834 10805
rect 8886 10745 9144 10805
rect 9196 10745 9200 10805
rect 8830 10735 9200 10745
rect 9230 11065 9600 11075
rect 9230 11005 9234 11065
rect 9286 11005 9544 11065
rect 9596 11005 9600 11065
rect 9230 10930 9600 11005
rect 9630 11065 10000 11075
rect 9630 11005 9634 11065
rect 9686 11005 9944 11065
rect 9996 11005 10000 11065
rect 9630 10930 10000 11005
rect 10030 11065 10400 11075
rect 10030 11005 10034 11065
rect 10086 11005 10344 11065
rect 10396 11005 10400 11065
rect 10030 10930 10400 11005
rect 9230 10890 10400 10930
rect 9230 10805 9600 10890
rect 9230 10745 9234 10805
rect 9286 10745 9544 10805
rect 9596 10745 9600 10805
rect 9230 10735 9600 10745
rect 9630 10805 10000 10890
rect 9630 10745 9634 10805
rect 9686 10745 9944 10805
rect 9996 10745 10000 10805
rect 9630 10735 10000 10745
rect 10030 10805 10400 10890
rect 10030 10745 10034 10805
rect 10086 10745 10344 10805
rect 10396 10745 10400 10805
rect 10030 10735 10400 10745
rect 10430 11065 10800 11075
rect 10430 11005 10434 11065
rect 10486 11005 10744 11065
rect 10796 11005 10800 11065
rect 10430 10930 10800 11005
rect 10830 11065 11200 11075
rect 10830 11005 10834 11065
rect 10886 11005 11144 11065
rect 11196 11005 11200 11065
rect 10830 10930 11200 11005
rect 10430 10890 11200 10930
rect 10430 10805 10800 10890
rect 10430 10745 10434 10805
rect 10486 10745 10744 10805
rect 10796 10745 10800 10805
rect 10430 10735 10800 10745
rect 10830 10805 11200 10890
rect 10830 10745 10834 10805
rect 10886 10745 11144 10805
rect 11196 10745 11200 10805
rect 10830 10735 11200 10745
rect 11230 11065 11600 11075
rect 11230 11005 11234 11065
rect 11286 11005 11544 11065
rect 11596 11005 11600 11065
rect 11230 10805 11600 11005
rect 11230 10745 11234 10805
rect 11286 10745 11544 10805
rect 11596 10745 11600 10805
rect 11230 10735 11600 10745
rect 11630 11065 12000 11075
rect 11630 11005 11634 11065
rect 11686 11005 11944 11065
rect 11996 11005 12000 11065
rect 11630 10805 12000 11005
rect 11630 10745 11634 10805
rect 11686 10745 11944 10805
rect 11996 10745 12000 10805
rect 11630 10735 12000 10745
rect 12030 11065 12400 11075
rect 12030 11005 12034 11065
rect 12086 11005 12344 11065
rect 12396 11005 12400 11065
rect 12030 10930 12400 11005
rect 12430 11065 12800 11075
rect 12430 11005 12434 11065
rect 12486 11005 12744 11065
rect 12796 11005 12800 11065
rect 12430 10930 12800 11005
rect 12830 11065 13200 11075
rect 12830 11005 12834 11065
rect 12886 11005 13144 11065
rect 13196 11005 13200 11065
rect 12830 10930 13200 11005
rect 12030 10890 13390 10930
rect 12030 10805 12400 10890
rect 12030 10745 12034 10805
rect 12086 10745 12344 10805
rect 12396 10745 12400 10805
rect 12030 10735 12400 10745
rect 12430 10805 12800 10890
rect 12430 10745 12434 10805
rect 12486 10745 12744 10805
rect 12796 10745 12800 10805
rect 12430 10735 12800 10745
rect 12830 10805 13200 10890
rect 12830 10745 12834 10805
rect 12886 10745 13144 10805
rect 13196 10745 13200 10805
rect 12830 10735 13200 10745
rect -330 10705 -324 10735
rect 30 10705 70 10735
rect 430 10705 470 10735
rect 830 10705 870 10735
rect 1230 10705 1270 10735
rect 1630 10705 1670 10735
rect 2030 10705 2070 10735
rect 2430 10705 2470 10735
rect 2830 10705 2870 10735
rect 3230 10705 3270 10735
rect 3630 10705 3670 10735
rect 4030 10705 4070 10735
rect 4430 10705 4470 10735
rect 4830 10705 4870 10735
rect 5230 10705 5270 10735
rect 5630 10705 5670 10735
rect 6030 10705 6070 10735
rect 6430 10705 6470 10735
rect 6830 10705 6870 10735
rect 7230 10705 7270 10735
rect 7630 10705 7670 10735
rect 8030 10705 8070 10735
rect 8430 10705 8470 10735
rect 8830 10705 8870 10735
rect 9230 10705 9270 10735
rect 9630 10705 9670 10735
rect 10030 10705 10070 10735
rect 10430 10705 10470 10735
rect 10830 10705 10870 10735
rect 11230 10705 11270 10735
rect 12030 10705 12070 10735
rect 12430 10705 12470 10735
rect -330 10695 0 10705
rect -314 10635 -56 10695
rect -4 10635 0 10695
rect -330 10435 0 10635
rect -314 10375 -56 10435
rect -4 10375 0 10435
rect -330 10365 0 10375
rect 30 10695 400 10705
rect 30 10635 34 10695
rect 86 10635 344 10695
rect 396 10635 400 10695
rect 30 10560 400 10635
rect 430 10695 800 10705
rect 430 10635 434 10695
rect 486 10635 744 10695
rect 796 10635 800 10695
rect 430 10560 800 10635
rect 830 10695 1200 10705
rect 830 10635 834 10695
rect 886 10635 1144 10695
rect 1196 10635 1200 10695
rect 830 10560 1200 10635
rect 1230 10695 1600 10705
rect 1230 10635 1234 10695
rect 1286 10635 1544 10695
rect 1596 10635 1600 10695
rect 1230 10560 1600 10635
rect 1630 10695 2000 10705
rect 1630 10635 1634 10695
rect 1686 10635 1944 10695
rect 1996 10635 2000 10695
rect 1630 10560 2000 10635
rect 2030 10695 2400 10705
rect 2030 10635 2034 10695
rect 2086 10635 2344 10695
rect 2396 10635 2400 10695
rect 2030 10560 2400 10635
rect 2430 10695 2800 10705
rect 2430 10635 2434 10695
rect 2486 10635 2744 10695
rect 2796 10635 2800 10695
rect 2430 10560 2800 10635
rect 30 10520 2800 10560
rect 30 10435 400 10520
rect 30 10375 34 10435
rect 86 10375 344 10435
rect 396 10375 400 10435
rect 30 10365 400 10375
rect 430 10435 800 10520
rect 430 10375 434 10435
rect 486 10375 744 10435
rect 796 10375 800 10435
rect 430 10365 800 10375
rect 830 10435 1200 10520
rect 830 10375 834 10435
rect 886 10375 1144 10435
rect 1196 10375 1200 10435
rect 830 10365 1200 10375
rect 1230 10435 1600 10520
rect 1230 10375 1234 10435
rect 1286 10375 1544 10435
rect 1596 10375 1600 10435
rect 1230 10365 1600 10375
rect 1630 10435 2000 10520
rect 1630 10375 1634 10435
rect 1686 10375 1944 10435
rect 1996 10375 2000 10435
rect 1630 10365 2000 10375
rect 2030 10435 2400 10520
rect 2030 10375 2034 10435
rect 2086 10375 2344 10435
rect 2396 10375 2400 10435
rect 2030 10365 2400 10375
rect 2430 10435 2800 10520
rect 2430 10375 2434 10435
rect 2486 10375 2744 10435
rect 2796 10375 2800 10435
rect 2430 10365 2800 10375
rect 2830 10695 3200 10705
rect 2830 10635 2834 10695
rect 2886 10635 3144 10695
rect 3196 10635 3200 10695
rect 2830 10560 3200 10635
rect 3230 10695 3600 10705
rect 3230 10635 3234 10695
rect 3286 10635 3544 10695
rect 3596 10635 3600 10695
rect 3230 10560 3600 10635
rect 3630 10695 4000 10705
rect 3630 10635 3634 10695
rect 3686 10635 3944 10695
rect 3996 10635 4000 10695
rect 3630 10560 4000 10635
rect 4030 10695 4400 10705
rect 4030 10635 4034 10695
rect 4086 10635 4344 10695
rect 4396 10635 4400 10695
rect 4030 10560 4400 10635
rect 4430 10695 4800 10705
rect 4430 10635 4434 10695
rect 4486 10635 4744 10695
rect 4796 10635 4800 10695
rect 4430 10560 4800 10635
rect 4830 10695 5200 10705
rect 4830 10635 4834 10695
rect 4886 10635 5144 10695
rect 5196 10635 5200 10695
rect 4830 10560 5200 10635
rect 5230 10695 5600 10705
rect 5230 10635 5234 10695
rect 5286 10635 5544 10695
rect 5596 10635 5600 10695
rect 5230 10560 5600 10635
rect 5630 10695 6000 10705
rect 5630 10635 5634 10695
rect 5686 10635 5944 10695
rect 5996 10635 6000 10695
rect 5630 10560 6000 10635
rect 2830 10520 6000 10560
rect 2830 10435 3200 10520
rect 2830 10375 2834 10435
rect 2886 10375 3144 10435
rect 3196 10375 3200 10435
rect 2830 10365 3200 10375
rect 3230 10435 3600 10520
rect 3230 10375 3234 10435
rect 3286 10375 3544 10435
rect 3596 10375 3600 10435
rect 3230 10365 3600 10375
rect 3630 10435 4000 10520
rect 3630 10375 3634 10435
rect 3686 10375 3944 10435
rect 3996 10375 4000 10435
rect 3630 10365 4000 10375
rect 4030 10435 4400 10520
rect 4030 10375 4034 10435
rect 4086 10375 4344 10435
rect 4396 10375 4400 10435
rect 4030 10365 4400 10375
rect 4430 10435 4800 10520
rect 4430 10375 4434 10435
rect 4486 10375 4744 10435
rect 4796 10375 4800 10435
rect 4430 10365 4800 10375
rect 4830 10435 5200 10520
rect 4830 10375 4834 10435
rect 4886 10375 5144 10435
rect 5196 10375 5200 10435
rect 4830 10365 5200 10375
rect 5230 10435 5600 10520
rect 5230 10375 5234 10435
rect 5286 10375 5544 10435
rect 5596 10375 5600 10435
rect 5230 10365 5600 10375
rect 5630 10435 6000 10520
rect 5630 10375 5634 10435
rect 5686 10375 5944 10435
rect 5996 10375 6000 10435
rect 5630 10365 6000 10375
rect 6030 10695 6400 10705
rect 6030 10635 6034 10695
rect 6086 10635 6344 10695
rect 6396 10635 6400 10695
rect 6030 10560 6400 10635
rect 6430 10695 6800 10705
rect 6430 10635 6434 10695
rect 6486 10635 6744 10695
rect 6796 10635 6800 10695
rect 6430 10560 6800 10635
rect 6830 10695 7200 10705
rect 6830 10635 6834 10695
rect 6886 10635 7144 10695
rect 7196 10635 7200 10695
rect 6830 10560 7200 10635
rect 7230 10695 7600 10705
rect 7230 10635 7234 10695
rect 7286 10635 7544 10695
rect 7596 10635 7600 10695
rect 7230 10560 7600 10635
rect 6030 10520 7600 10560
rect 6030 10435 6400 10520
rect 6030 10375 6034 10435
rect 6086 10375 6344 10435
rect 6396 10375 6400 10435
rect 6030 10365 6400 10375
rect 6430 10435 6800 10520
rect 6430 10375 6434 10435
rect 6486 10375 6744 10435
rect 6796 10375 6800 10435
rect 6430 10365 6800 10375
rect 6830 10435 7200 10520
rect 6830 10375 6834 10435
rect 6886 10375 7144 10435
rect 7196 10375 7200 10435
rect 6830 10365 7200 10375
rect 7230 10435 7600 10520
rect 7230 10375 7234 10435
rect 7286 10375 7544 10435
rect 7596 10375 7600 10435
rect 7230 10365 7600 10375
rect 7630 10695 8000 10705
rect 7630 10635 7634 10695
rect 7686 10635 7944 10695
rect 7996 10635 8000 10695
rect 7630 10560 8000 10635
rect 8030 10695 8400 10705
rect 8030 10635 8034 10695
rect 8086 10635 8344 10695
rect 8396 10635 8400 10695
rect 8030 10560 8400 10635
rect 7630 10520 8400 10560
rect 7630 10435 8000 10520
rect 7630 10375 7634 10435
rect 7686 10375 7944 10435
rect 7996 10375 8000 10435
rect 7630 10365 8000 10375
rect 8030 10435 8400 10520
rect 8030 10375 8034 10435
rect 8086 10375 8344 10435
rect 8396 10375 8400 10435
rect 8030 10365 8400 10375
rect 8430 10695 8800 10705
rect 8430 10635 8434 10695
rect 8486 10635 8744 10695
rect 8796 10635 8800 10695
rect 8430 10435 8800 10635
rect 8430 10375 8434 10435
rect 8486 10375 8744 10435
rect 8796 10375 8800 10435
rect 8430 10365 8800 10375
rect 8830 10695 9200 10705
rect 8830 10635 8834 10695
rect 8886 10635 9144 10695
rect 9196 10635 9200 10695
rect 8830 10435 9200 10635
rect 8830 10375 8834 10435
rect 8886 10375 9144 10435
rect 9196 10375 9200 10435
rect 8830 10365 9200 10375
rect 9230 10695 9600 10705
rect 9230 10635 9234 10695
rect 9286 10635 9544 10695
rect 9596 10635 9600 10695
rect 9230 10560 9600 10635
rect 9630 10695 10000 10705
rect 9630 10635 9634 10695
rect 9686 10635 9944 10695
rect 9996 10635 10000 10695
rect 9630 10560 10000 10635
rect 10030 10695 10400 10705
rect 10030 10635 10034 10695
rect 10086 10635 10344 10695
rect 10396 10635 10400 10695
rect 10030 10560 10400 10635
rect 9230 10520 10400 10560
rect 9230 10435 9600 10520
rect 9230 10375 9234 10435
rect 9286 10375 9544 10435
rect 9596 10375 9600 10435
rect 9230 10365 9600 10375
rect 9630 10435 10000 10520
rect 9630 10375 9634 10435
rect 9686 10375 9944 10435
rect 9996 10375 10000 10435
rect 9630 10365 10000 10375
rect 10030 10435 10400 10520
rect 10030 10375 10034 10435
rect 10086 10375 10344 10435
rect 10396 10375 10400 10435
rect 10030 10365 10400 10375
rect 10430 10695 10800 10705
rect 10430 10635 10434 10695
rect 10486 10635 10744 10695
rect 10796 10635 10800 10695
rect 10430 10560 10800 10635
rect 10830 10695 11200 10705
rect 10830 10635 10834 10695
rect 10886 10635 11144 10695
rect 11196 10635 11200 10695
rect 10830 10560 11200 10635
rect 10430 10520 11200 10560
rect 10430 10435 10800 10520
rect 10430 10375 10434 10435
rect 10486 10375 10744 10435
rect 10796 10375 10800 10435
rect 10430 10365 10800 10375
rect 10830 10435 11200 10520
rect 10830 10375 10834 10435
rect 10886 10375 11144 10435
rect 11196 10375 11200 10435
rect 10830 10365 11200 10375
rect 11230 10695 11600 10705
rect 11230 10635 11234 10695
rect 11286 10635 11544 10695
rect 11596 10635 11600 10695
rect 11230 10560 11600 10635
rect 11630 10695 12000 10705
rect 11630 10635 11634 10695
rect 11686 10635 11944 10695
rect 11996 10635 12000 10695
rect 11630 10560 12000 10635
rect 12030 10695 12400 10705
rect 12030 10635 12034 10695
rect 12086 10635 12344 10695
rect 12396 10635 12400 10695
rect 12030 10560 12400 10635
rect 12430 10695 12800 10705
rect 12430 10635 12434 10695
rect 12486 10635 12744 10695
rect 12796 10635 12800 10695
rect 12430 10560 12800 10635
rect 12830 10695 13200 10705
rect 12830 10635 12834 10695
rect 12886 10635 13144 10695
rect 13196 10635 13200 10695
rect 12830 10560 13200 10635
rect 11230 10520 13200 10560
rect 11230 10435 11600 10520
rect 11230 10375 11234 10435
rect 11286 10375 11544 10435
rect 11596 10375 11600 10435
rect 11230 10365 11600 10375
rect 11630 10435 12000 10520
rect 11630 10375 11634 10435
rect 11686 10375 11944 10435
rect 11996 10375 12000 10435
rect 11630 10365 12000 10375
rect 12030 10435 12400 10520
rect 12030 10375 12034 10435
rect 12086 10375 12344 10435
rect 12396 10375 12400 10435
rect 12030 10365 12400 10375
rect 12430 10435 12800 10520
rect 12430 10375 12434 10435
rect 12486 10375 12744 10435
rect 12796 10375 12800 10435
rect 12430 10365 12800 10375
rect 12830 10435 13200 10520
rect 12830 10375 12834 10435
rect 12886 10375 13144 10435
rect 13196 10375 13200 10435
rect 12830 10365 13200 10375
rect -330 10335 -324 10365
rect 30 10335 70 10365
rect 430 10335 470 10365
rect 830 10335 870 10365
rect 1230 10335 1270 10365
rect 1630 10335 1670 10365
rect 2030 10335 2070 10365
rect 2430 10335 2470 10365
rect 2830 10335 2870 10365
rect 3230 10335 3270 10365
rect 3630 10335 3670 10365
rect 4030 10335 4070 10365
rect 4430 10335 4470 10365
rect 4830 10335 4870 10365
rect 5230 10335 5270 10365
rect 5630 10335 5670 10365
rect 6030 10335 6070 10365
rect 6430 10335 6470 10365
rect 6830 10335 6870 10365
rect 7230 10335 7270 10365
rect 7630 10335 7670 10365
rect 8030 10335 8070 10365
rect 8430 10335 8470 10365
rect 8830 10335 8870 10365
rect 9230 10335 9270 10365
rect 9630 10335 9670 10365
rect 10030 10335 10070 10365
rect 10430 10335 10470 10365
rect 10830 10335 10870 10365
rect -330 10325 0 10335
rect -314 10265 -56 10325
rect -4 10265 0 10325
rect -330 10065 0 10265
rect -314 10005 -56 10065
rect -4 10005 0 10065
rect -330 9995 0 10005
rect 30 10325 400 10335
rect 30 10265 34 10325
rect 86 10265 344 10325
rect 396 10265 400 10325
rect 30 10190 400 10265
rect 430 10325 800 10335
rect 430 10265 434 10325
rect 486 10265 744 10325
rect 796 10265 800 10325
rect 430 10190 800 10265
rect 830 10325 1200 10335
rect 830 10265 834 10325
rect 886 10265 1144 10325
rect 1196 10265 1200 10325
rect 830 10190 1200 10265
rect 1230 10325 1600 10335
rect 1230 10265 1234 10325
rect 1286 10265 1544 10325
rect 1596 10265 1600 10325
rect 1230 10190 1600 10265
rect 1630 10325 2000 10335
rect 1630 10265 1634 10325
rect 1686 10265 1944 10325
rect 1996 10265 2000 10325
rect 1630 10190 2000 10265
rect 2030 10325 2400 10335
rect 2030 10265 2034 10325
rect 2086 10265 2344 10325
rect 2396 10265 2400 10325
rect 2030 10190 2400 10265
rect 2430 10325 2800 10335
rect 2430 10265 2434 10325
rect 2486 10265 2744 10325
rect 2796 10265 2800 10325
rect 2430 10190 2800 10265
rect 30 10150 2800 10190
rect 30 10065 400 10150
rect 30 10005 34 10065
rect 86 10005 344 10065
rect 396 10005 400 10065
rect 30 9995 400 10005
rect 430 10065 800 10150
rect 430 10005 434 10065
rect 486 10005 744 10065
rect 796 10005 800 10065
rect 430 9995 800 10005
rect 830 10065 1200 10150
rect 830 10005 834 10065
rect 886 10005 1144 10065
rect 1196 10005 1200 10065
rect 830 9995 1200 10005
rect 1230 10065 1600 10150
rect 1230 10005 1234 10065
rect 1286 10005 1544 10065
rect 1596 10005 1600 10065
rect 1230 9995 1600 10005
rect 1630 10065 2000 10150
rect 1630 10005 1634 10065
rect 1686 10005 1944 10065
rect 1996 10005 2000 10065
rect 1630 9995 2000 10005
rect 2030 10065 2400 10150
rect 2030 10005 2034 10065
rect 2086 10005 2344 10065
rect 2396 10005 2400 10065
rect 2030 9995 2400 10005
rect 2430 10065 2800 10150
rect 2430 10005 2434 10065
rect 2486 10005 2744 10065
rect 2796 10005 2800 10065
rect 2430 9995 2800 10005
rect 2830 10325 3200 10335
rect 2830 10265 2834 10325
rect 2886 10265 3144 10325
rect 3196 10265 3200 10325
rect 2830 10190 3200 10265
rect 3230 10325 3600 10335
rect 3230 10265 3234 10325
rect 3286 10265 3544 10325
rect 3596 10265 3600 10325
rect 3230 10190 3600 10265
rect 3630 10325 4000 10335
rect 3630 10265 3634 10325
rect 3686 10265 3944 10325
rect 3996 10265 4000 10325
rect 3630 10190 4000 10265
rect 4030 10325 4400 10335
rect 4030 10265 4034 10325
rect 4086 10265 4344 10325
rect 4396 10265 4400 10325
rect 4030 10190 4400 10265
rect 4430 10325 4800 10335
rect 4430 10265 4434 10325
rect 4486 10265 4744 10325
rect 4796 10265 4800 10325
rect 4430 10190 4800 10265
rect 4830 10325 5200 10335
rect 4830 10265 4834 10325
rect 4886 10265 5144 10325
rect 5196 10265 5200 10325
rect 4830 10190 5200 10265
rect 5230 10325 5600 10335
rect 5230 10265 5234 10325
rect 5286 10265 5544 10325
rect 5596 10265 5600 10325
rect 5230 10190 5600 10265
rect 5630 10325 6000 10335
rect 5630 10265 5634 10325
rect 5686 10265 5944 10325
rect 5996 10265 6000 10325
rect 5630 10190 6000 10265
rect 2830 10150 6000 10190
rect 2830 10065 3200 10150
rect 2830 10005 2834 10065
rect 2886 10005 3144 10065
rect 3196 10005 3200 10065
rect 2830 9995 3200 10005
rect 3230 10065 3600 10150
rect 3230 10005 3234 10065
rect 3286 10005 3544 10065
rect 3596 10005 3600 10065
rect 3230 9995 3600 10005
rect 3630 10065 4000 10150
rect 3630 10005 3634 10065
rect 3686 10005 3944 10065
rect 3996 10005 4000 10065
rect 3630 9995 4000 10005
rect 4030 10065 4400 10150
rect 4030 10005 4034 10065
rect 4086 10005 4344 10065
rect 4396 10005 4400 10065
rect 4030 9995 4400 10005
rect 4430 10065 4800 10150
rect 4430 10005 4434 10065
rect 4486 10005 4744 10065
rect 4796 10005 4800 10065
rect 4430 9995 4800 10005
rect 4830 10065 5200 10150
rect 4830 10005 4834 10065
rect 4886 10005 5144 10065
rect 5196 10005 5200 10065
rect 4830 9995 5200 10005
rect 5230 10065 5600 10150
rect 5230 10005 5234 10065
rect 5286 10005 5544 10065
rect 5596 10005 5600 10065
rect 5230 9995 5600 10005
rect 5630 10065 6000 10150
rect 5630 10005 5634 10065
rect 5686 10005 5944 10065
rect 5996 10005 6000 10065
rect 5630 9995 6000 10005
rect 6030 10325 6400 10335
rect 6030 10265 6034 10325
rect 6086 10265 6344 10325
rect 6396 10265 6400 10325
rect 6030 10190 6400 10265
rect 6430 10325 6800 10335
rect 6430 10265 6434 10325
rect 6486 10265 6744 10325
rect 6796 10265 6800 10325
rect 6430 10190 6800 10265
rect 6830 10325 7200 10335
rect 6830 10265 6834 10325
rect 6886 10265 7144 10325
rect 7196 10265 7200 10325
rect 6830 10190 7200 10265
rect 7230 10325 7600 10335
rect 7230 10265 7234 10325
rect 7286 10265 7544 10325
rect 7596 10265 7600 10325
rect 7230 10190 7600 10265
rect 6030 10150 7600 10190
rect 6030 10065 6400 10150
rect 6030 10005 6034 10065
rect 6086 10005 6344 10065
rect 6396 10005 6400 10065
rect 6030 9995 6400 10005
rect 6430 10065 6800 10150
rect 6430 10005 6434 10065
rect 6486 10005 6744 10065
rect 6796 10005 6800 10065
rect 6430 9995 6800 10005
rect 6830 10065 7200 10150
rect 6830 10005 6834 10065
rect 6886 10005 7144 10065
rect 7196 10005 7200 10065
rect 6830 9995 7200 10005
rect 7230 10065 7600 10150
rect 7230 10005 7234 10065
rect 7286 10005 7544 10065
rect 7596 10005 7600 10065
rect 7230 9995 7600 10005
rect 7630 10325 8000 10335
rect 7630 10265 7634 10325
rect 7686 10265 7944 10325
rect 7996 10265 8000 10325
rect 7630 10190 8000 10265
rect 8030 10325 8400 10335
rect 8030 10265 8034 10325
rect 8086 10265 8344 10325
rect 8396 10265 8400 10325
rect 8030 10190 8400 10265
rect 7630 10150 8400 10190
rect 7630 10065 8000 10150
rect 7630 10005 7634 10065
rect 7686 10005 7944 10065
rect 7996 10005 8000 10065
rect 7630 9995 8000 10005
rect 8030 10065 8400 10150
rect 8030 10005 8034 10065
rect 8086 10005 8344 10065
rect 8396 10005 8400 10065
rect 8030 9995 8400 10005
rect 8430 10325 8800 10335
rect 8430 10265 8434 10325
rect 8486 10265 8744 10325
rect 8796 10265 8800 10325
rect 8430 10065 8800 10265
rect 8430 10005 8434 10065
rect 8486 10005 8744 10065
rect 8796 10005 8800 10065
rect 8430 9995 8800 10005
rect 8830 10325 9200 10335
rect 8830 10265 8834 10325
rect 8886 10265 9144 10325
rect 9196 10265 9200 10325
rect 8830 10065 9200 10265
rect 8830 10005 8834 10065
rect 8886 10005 9144 10065
rect 9196 10005 9200 10065
rect 8830 9995 9200 10005
rect 9230 10325 9600 10335
rect 9230 10265 9234 10325
rect 9286 10265 9544 10325
rect 9596 10265 9600 10325
rect 9230 10190 9600 10265
rect 9630 10325 10000 10335
rect 9630 10265 9634 10325
rect 9686 10265 9944 10325
rect 9996 10265 10000 10325
rect 9630 10190 10000 10265
rect 10030 10325 10400 10335
rect 10030 10265 10034 10325
rect 10086 10265 10344 10325
rect 10396 10265 10400 10325
rect 10030 10190 10400 10265
rect 9230 10150 10400 10190
rect 9230 10065 9600 10150
rect 9230 10005 9234 10065
rect 9286 10005 9544 10065
rect 9596 10005 9600 10065
rect 9230 9995 9600 10005
rect 9630 10065 10000 10150
rect 9630 10005 9634 10065
rect 9686 10005 9944 10065
rect 9996 10005 10000 10065
rect 9630 9995 10000 10005
rect 10030 10065 10400 10150
rect 10030 10005 10034 10065
rect 10086 10005 10344 10065
rect 10396 10005 10400 10065
rect 10030 9995 10400 10005
rect 10430 10325 10800 10335
rect 10430 10265 10434 10325
rect 10486 10265 10744 10325
rect 10796 10265 10800 10325
rect 10430 10190 10800 10265
rect 10830 10325 11200 10335
rect 10830 10265 10834 10325
rect 10886 10265 11144 10325
rect 11196 10265 11200 10325
rect 10830 10190 11200 10265
rect 11230 10325 11600 10335
rect 11230 10265 11234 10325
rect 11286 10265 11544 10325
rect 11596 10265 11600 10325
rect 11230 10190 11600 10265
rect 11630 10325 12000 10335
rect 11630 10265 11634 10325
rect 11686 10265 11944 10325
rect 11996 10265 12000 10325
rect 11630 10190 12000 10265
rect 12030 10325 12400 10335
rect 12030 10265 12034 10325
rect 12086 10265 12344 10325
rect 12396 10265 12400 10325
rect 12030 10190 12400 10265
rect 12430 10325 12800 10335
rect 12430 10265 12434 10325
rect 12486 10265 12744 10325
rect 12796 10265 12800 10325
rect 12430 10190 12800 10265
rect 12830 10325 13200 10335
rect 12830 10265 12834 10325
rect 12886 10265 13144 10325
rect 13196 10265 13200 10325
rect 12830 10190 13200 10265
rect 10430 10150 13390 10190
rect 10430 10065 10800 10150
rect 10430 10005 10434 10065
rect 10486 10005 10744 10065
rect 10796 10005 10800 10065
rect 10430 9995 10800 10005
rect 10830 10065 11200 10150
rect 10830 10005 10834 10065
rect 10886 10005 11144 10065
rect 11196 10005 11200 10065
rect 10830 9995 11200 10005
rect 11230 10065 11600 10150
rect 11230 10005 11234 10065
rect 11286 10005 11544 10065
rect 11596 10005 11600 10065
rect 11230 9995 11600 10005
rect 11630 10065 12000 10150
rect 11630 10005 11634 10065
rect 11686 10005 11944 10065
rect 11996 10005 12000 10065
rect 11630 9995 12000 10005
rect 12030 10065 12400 10150
rect 12030 10005 12034 10065
rect 12086 10005 12344 10065
rect 12396 10005 12400 10065
rect 12030 9995 12400 10005
rect 12430 10065 12800 10150
rect 12430 10005 12434 10065
rect 12486 10005 12744 10065
rect 12796 10005 12800 10065
rect 12430 9995 12800 10005
rect 12830 10065 13200 10150
rect 12830 10005 12834 10065
rect 12886 10005 13144 10065
rect 13196 10005 13200 10065
rect 12830 9995 13200 10005
rect -330 9965 -324 9995
rect 30 9965 70 9995
rect 430 9965 470 9995
rect 830 9965 870 9995
rect 1230 9965 1270 9995
rect 1630 9965 1670 9995
rect 2030 9965 2070 9995
rect 2430 9965 2470 9995
rect 2830 9965 2870 9995
rect 3230 9965 3270 9995
rect 3630 9965 3670 9995
rect 4030 9965 4070 9995
rect 4430 9965 4470 9995
rect 4830 9965 4870 9995
rect 5230 9965 5270 9995
rect 5630 9965 5670 9995
rect 6030 9965 6070 9995
rect 6430 9965 6470 9995
rect 6830 9965 6870 9995
rect 7230 9965 7270 9995
rect 7630 9965 7670 9995
rect 8030 9965 8070 9995
rect 8430 9965 8470 9995
rect 8830 9965 8870 9995
rect 9230 9965 9270 9995
rect 9630 9965 9670 9995
rect 10030 9965 10070 9995
rect -330 9955 0 9965
rect -314 9895 -56 9955
rect -4 9895 0 9955
rect -330 9695 0 9895
rect -314 9635 -56 9695
rect -4 9635 0 9695
rect -330 9625 0 9635
rect 30 9955 400 9965
rect 30 9895 34 9955
rect 86 9895 344 9955
rect 396 9895 400 9955
rect 30 9820 400 9895
rect 430 9955 800 9965
rect 430 9895 434 9955
rect 486 9895 744 9955
rect 796 9895 800 9955
rect 430 9820 800 9895
rect 830 9955 1200 9965
rect 830 9895 834 9955
rect 886 9895 1144 9955
rect 1196 9895 1200 9955
rect 830 9820 1200 9895
rect 1230 9955 1600 9965
rect 1230 9895 1234 9955
rect 1286 9895 1544 9955
rect 1596 9895 1600 9955
rect 1230 9820 1600 9895
rect 1630 9955 2000 9965
rect 1630 9895 1634 9955
rect 1686 9895 1944 9955
rect 1996 9895 2000 9955
rect 1630 9820 2000 9895
rect 2030 9955 2400 9965
rect 2030 9895 2034 9955
rect 2086 9895 2344 9955
rect 2396 9895 2400 9955
rect 2030 9820 2400 9895
rect 2430 9955 2800 9965
rect 2430 9895 2434 9955
rect 2486 9895 2744 9955
rect 2796 9895 2800 9955
rect 2430 9820 2800 9895
rect 30 9780 2800 9820
rect 30 9695 400 9780
rect 30 9635 34 9695
rect 86 9635 344 9695
rect 396 9635 400 9695
rect 30 9625 400 9635
rect 430 9695 800 9780
rect 430 9635 434 9695
rect 486 9635 744 9695
rect 796 9635 800 9695
rect 430 9625 800 9635
rect 830 9695 1200 9780
rect 830 9635 834 9695
rect 886 9635 1144 9695
rect 1196 9635 1200 9695
rect 830 9625 1200 9635
rect 1230 9695 1600 9780
rect 1230 9635 1234 9695
rect 1286 9635 1544 9695
rect 1596 9635 1600 9695
rect 1230 9625 1600 9635
rect 1630 9695 2000 9780
rect 1630 9635 1634 9695
rect 1686 9635 1944 9695
rect 1996 9635 2000 9695
rect 1630 9625 2000 9635
rect 2030 9695 2400 9780
rect 2030 9635 2034 9695
rect 2086 9635 2344 9695
rect 2396 9635 2400 9695
rect 2030 9625 2400 9635
rect 2430 9695 2800 9780
rect 2430 9635 2434 9695
rect 2486 9635 2744 9695
rect 2796 9635 2800 9695
rect 2430 9625 2800 9635
rect 2830 9955 3200 9965
rect 2830 9895 2834 9955
rect 2886 9895 3144 9955
rect 3196 9895 3200 9955
rect 2830 9820 3200 9895
rect 3230 9955 3600 9965
rect 3230 9895 3234 9955
rect 3286 9895 3544 9955
rect 3596 9895 3600 9955
rect 3230 9820 3600 9895
rect 3630 9955 4000 9965
rect 3630 9895 3634 9955
rect 3686 9895 3944 9955
rect 3996 9895 4000 9955
rect 3630 9820 4000 9895
rect 4030 9955 4400 9965
rect 4030 9895 4034 9955
rect 4086 9895 4344 9955
rect 4396 9895 4400 9955
rect 4030 9820 4400 9895
rect 4430 9955 4800 9965
rect 4430 9895 4434 9955
rect 4486 9895 4744 9955
rect 4796 9895 4800 9955
rect 4430 9820 4800 9895
rect 4830 9955 5200 9965
rect 4830 9895 4834 9955
rect 4886 9895 5144 9955
rect 5196 9895 5200 9955
rect 4830 9820 5200 9895
rect 5230 9955 5600 9965
rect 5230 9895 5234 9955
rect 5286 9895 5544 9955
rect 5596 9895 5600 9955
rect 5230 9820 5600 9895
rect 5630 9955 6000 9965
rect 5630 9895 5634 9955
rect 5686 9895 5944 9955
rect 5996 9895 6000 9955
rect 5630 9820 6000 9895
rect 2830 9780 6000 9820
rect 2830 9695 3200 9780
rect 2830 9635 2834 9695
rect 2886 9635 3144 9695
rect 3196 9635 3200 9695
rect 2830 9625 3200 9635
rect 3230 9695 3600 9780
rect 3230 9635 3234 9695
rect 3286 9635 3544 9695
rect 3596 9635 3600 9695
rect 3230 9625 3600 9635
rect 3630 9695 4000 9780
rect 3630 9635 3634 9695
rect 3686 9635 3944 9695
rect 3996 9635 4000 9695
rect 3630 9625 4000 9635
rect 4030 9695 4400 9780
rect 4030 9635 4034 9695
rect 4086 9635 4344 9695
rect 4396 9635 4400 9695
rect 4030 9625 4400 9635
rect 4430 9695 4800 9780
rect 4430 9635 4434 9695
rect 4486 9635 4744 9695
rect 4796 9635 4800 9695
rect 4430 9625 4800 9635
rect 4830 9695 5200 9780
rect 4830 9635 4834 9695
rect 4886 9635 5144 9695
rect 5196 9635 5200 9695
rect 4830 9625 5200 9635
rect 5230 9695 5600 9780
rect 5230 9635 5234 9695
rect 5286 9635 5544 9695
rect 5596 9635 5600 9695
rect 5230 9625 5600 9635
rect 5630 9695 6000 9780
rect 5630 9635 5634 9695
rect 5686 9635 5944 9695
rect 5996 9635 6000 9695
rect 5630 9625 6000 9635
rect 6030 9955 6400 9965
rect 6030 9895 6034 9955
rect 6086 9895 6344 9955
rect 6396 9895 6400 9955
rect 6030 9820 6400 9895
rect 6430 9955 6800 9965
rect 6430 9895 6434 9955
rect 6486 9895 6744 9955
rect 6796 9895 6800 9955
rect 6430 9820 6800 9895
rect 6830 9955 7200 9965
rect 6830 9895 6834 9955
rect 6886 9895 7144 9955
rect 7196 9895 7200 9955
rect 6830 9820 7200 9895
rect 7230 9955 7600 9965
rect 7230 9895 7234 9955
rect 7286 9895 7544 9955
rect 7596 9895 7600 9955
rect 7230 9820 7600 9895
rect 6030 9780 7600 9820
rect 6030 9695 6400 9780
rect 6030 9635 6034 9695
rect 6086 9635 6344 9695
rect 6396 9635 6400 9695
rect 6030 9625 6400 9635
rect 6430 9695 6800 9780
rect 6430 9635 6434 9695
rect 6486 9635 6744 9695
rect 6796 9635 6800 9695
rect 6430 9625 6800 9635
rect 6830 9695 7200 9780
rect 6830 9635 6834 9695
rect 6886 9635 7144 9695
rect 7196 9635 7200 9695
rect 6830 9625 7200 9635
rect 7230 9695 7600 9780
rect 7230 9635 7234 9695
rect 7286 9635 7544 9695
rect 7596 9635 7600 9695
rect 7230 9625 7600 9635
rect 7630 9955 8000 9965
rect 7630 9895 7634 9955
rect 7686 9895 7944 9955
rect 7996 9895 8000 9955
rect 7630 9820 8000 9895
rect 8030 9955 8400 9965
rect 8030 9895 8034 9955
rect 8086 9895 8344 9955
rect 8396 9895 8400 9955
rect 8030 9820 8400 9895
rect 7630 9780 8400 9820
rect 7630 9695 8000 9780
rect 7630 9635 7634 9695
rect 7686 9635 7944 9695
rect 7996 9635 8000 9695
rect 7630 9625 8000 9635
rect 8030 9695 8400 9780
rect 8030 9635 8034 9695
rect 8086 9635 8344 9695
rect 8396 9635 8400 9695
rect 8030 9625 8400 9635
rect 8430 9955 8800 9965
rect 8430 9895 8434 9955
rect 8486 9895 8744 9955
rect 8796 9895 8800 9955
rect 8430 9695 8800 9895
rect 8430 9635 8434 9695
rect 8486 9635 8744 9695
rect 8796 9635 8800 9695
rect 8430 9625 8800 9635
rect 8830 9955 9200 9965
rect 8830 9895 8834 9955
rect 8886 9895 9144 9955
rect 9196 9895 9200 9955
rect 8830 9695 9200 9895
rect 8830 9635 8834 9695
rect 8886 9635 9144 9695
rect 9196 9635 9200 9695
rect 8830 9625 9200 9635
rect 9230 9955 9600 9965
rect 9230 9895 9234 9955
rect 9286 9895 9544 9955
rect 9596 9895 9600 9955
rect 9230 9820 9600 9895
rect 9630 9955 10000 9965
rect 9630 9895 9634 9955
rect 9686 9895 9944 9955
rect 9996 9895 10000 9955
rect 9630 9820 10000 9895
rect 10030 9955 10400 9965
rect 10030 9895 10034 9955
rect 10086 9895 10344 9955
rect 10396 9895 10400 9955
rect 10030 9820 10400 9895
rect 10430 9955 10800 9965
rect 10430 9895 10434 9955
rect 10486 9895 10744 9955
rect 10796 9895 10800 9955
rect 10430 9820 10800 9895
rect 10830 9955 11200 9965
rect 10830 9895 10834 9955
rect 10886 9895 11144 9955
rect 11196 9895 11200 9955
rect 10830 9820 11200 9895
rect 11230 9955 11600 9965
rect 11230 9895 11234 9955
rect 11286 9895 11544 9955
rect 11596 9895 11600 9955
rect 11230 9820 11600 9895
rect 11630 9955 12000 9965
rect 11630 9895 11634 9955
rect 11686 9895 11944 9955
rect 11996 9895 12000 9955
rect 11630 9820 12000 9895
rect 12030 9955 12400 9965
rect 12030 9895 12034 9955
rect 12086 9895 12344 9955
rect 12396 9895 12400 9955
rect 12030 9820 12400 9895
rect 12430 9955 12800 9965
rect 12430 9895 12434 9955
rect 12486 9895 12744 9955
rect 12796 9895 12800 9955
rect 12430 9820 12800 9895
rect 12830 9955 13200 9965
rect 12830 9895 12834 9955
rect 12886 9895 13144 9955
rect 13196 9895 13200 9955
rect 12830 9820 13200 9895
rect 9230 9780 13390 9820
rect 9230 9695 9600 9780
rect 9230 9635 9234 9695
rect 9286 9635 9544 9695
rect 9596 9635 9600 9695
rect 9230 9625 9600 9635
rect 9630 9695 10000 9780
rect 9630 9635 9634 9695
rect 9686 9635 9944 9695
rect 9996 9635 10000 9695
rect 9630 9625 10000 9635
rect 10030 9695 10400 9780
rect 10030 9635 10034 9695
rect 10086 9635 10344 9695
rect 10396 9635 10400 9695
rect 10030 9625 10400 9635
rect 10430 9695 10800 9780
rect 10430 9635 10434 9695
rect 10486 9635 10744 9695
rect 10796 9635 10800 9695
rect 10430 9625 10800 9635
rect 10830 9695 11200 9780
rect 10830 9635 10834 9695
rect 10886 9635 11144 9695
rect 11196 9635 11200 9695
rect 10830 9625 11200 9635
rect 11230 9695 11600 9780
rect 11230 9635 11234 9695
rect 11286 9635 11544 9695
rect 11596 9635 11600 9695
rect 11230 9625 11600 9635
rect 11630 9695 12000 9780
rect 11630 9635 11634 9695
rect 11686 9635 11944 9695
rect 11996 9635 12000 9695
rect 11630 9625 12000 9635
rect 12030 9695 12400 9780
rect 12030 9635 12034 9695
rect 12086 9635 12344 9695
rect 12396 9635 12400 9695
rect 12030 9625 12400 9635
rect 12430 9695 12800 9780
rect 12430 9635 12434 9695
rect 12486 9635 12744 9695
rect 12796 9635 12800 9695
rect 12430 9625 12800 9635
rect 12830 9695 13200 9780
rect 12830 9635 12834 9695
rect 12886 9635 13144 9695
rect 13196 9635 13200 9695
rect 12830 9625 13200 9635
rect -330 9595 -324 9625
rect 30 9595 70 9625
rect 430 9595 470 9625
rect 830 9595 870 9625
rect 1230 9595 1270 9625
rect 1630 9595 1670 9625
rect 2030 9595 2070 9625
rect 2430 9595 2470 9625
rect 2830 9595 2870 9625
rect 3230 9595 3270 9625
rect 3630 9595 3670 9625
rect 4030 9595 4070 9625
rect 4430 9595 4470 9625
rect 4830 9595 4870 9625
rect 5230 9595 5270 9625
rect 5630 9595 5670 9625
rect 6030 9595 6070 9625
rect 6430 9595 6470 9625
rect 6830 9595 6870 9625
rect 7230 9595 7270 9625
rect 7630 9595 7670 9625
rect 8030 9595 8070 9625
rect 8430 9595 8470 9625
rect 8830 9595 8870 9625
rect 9230 9595 9270 9625
rect 9630 9595 9670 9625
rect 10030 9595 10070 9625
rect 10430 9595 10470 9625
rect 10830 9595 10870 9625
rect 11230 9595 11270 9625
rect 11630 9595 11670 9625
rect 12030 9595 12070 9625
rect 12430 9595 12470 9625
rect -330 9585 0 9595
rect -314 9525 -56 9585
rect -4 9525 0 9585
rect -330 9325 0 9525
rect -314 9265 -56 9325
rect -4 9265 0 9325
rect -330 9255 0 9265
rect 30 9585 400 9595
rect 30 9525 34 9585
rect 86 9525 344 9585
rect 396 9525 400 9585
rect 30 9450 400 9525
rect 430 9585 800 9595
rect 430 9525 434 9585
rect 486 9525 744 9585
rect 796 9525 800 9585
rect 430 9450 800 9525
rect 830 9585 1200 9595
rect 830 9525 834 9585
rect 886 9525 1144 9585
rect 1196 9525 1200 9585
rect 830 9450 1200 9525
rect 1230 9585 1600 9595
rect 1230 9525 1234 9585
rect 1286 9525 1544 9585
rect 1596 9525 1600 9585
rect 1230 9450 1600 9525
rect 1630 9585 2000 9595
rect 1630 9525 1634 9585
rect 1686 9525 1944 9585
rect 1996 9525 2000 9585
rect 1630 9450 2000 9525
rect 2030 9585 2400 9595
rect 2030 9525 2034 9585
rect 2086 9525 2344 9585
rect 2396 9525 2400 9585
rect 2030 9450 2400 9525
rect 2430 9585 2800 9595
rect 2430 9525 2434 9585
rect 2486 9525 2744 9585
rect 2796 9525 2800 9585
rect 2430 9450 2800 9525
rect 30 9410 2800 9450
rect 30 9325 400 9410
rect 30 9265 34 9325
rect 86 9265 344 9325
rect 396 9265 400 9325
rect 30 9255 400 9265
rect 430 9325 800 9410
rect 430 9265 434 9325
rect 486 9265 744 9325
rect 796 9265 800 9325
rect 430 9255 800 9265
rect 830 9325 1200 9410
rect 830 9265 834 9325
rect 886 9265 1144 9325
rect 1196 9265 1200 9325
rect 830 9255 1200 9265
rect 1230 9325 1600 9410
rect 1230 9265 1234 9325
rect 1286 9265 1544 9325
rect 1596 9265 1600 9325
rect 1230 9255 1600 9265
rect 1630 9325 2000 9410
rect 1630 9265 1634 9325
rect 1686 9265 1944 9325
rect 1996 9265 2000 9325
rect 1630 9255 2000 9265
rect 2030 9325 2400 9410
rect 2030 9265 2034 9325
rect 2086 9265 2344 9325
rect 2396 9265 2400 9325
rect 2030 9255 2400 9265
rect 2430 9325 2800 9410
rect 2430 9265 2434 9325
rect 2486 9265 2744 9325
rect 2796 9265 2800 9325
rect 2430 9255 2800 9265
rect 2830 9585 3200 9595
rect 2830 9525 2834 9585
rect 2886 9525 3144 9585
rect 3196 9525 3200 9585
rect 2830 9450 3200 9525
rect 3230 9585 3600 9595
rect 3230 9525 3234 9585
rect 3286 9525 3544 9585
rect 3596 9525 3600 9585
rect 3230 9450 3600 9525
rect 3630 9585 4000 9595
rect 3630 9525 3634 9585
rect 3686 9525 3944 9585
rect 3996 9525 4000 9585
rect 3630 9450 4000 9525
rect 4030 9585 4400 9595
rect 4030 9525 4034 9585
rect 4086 9525 4344 9585
rect 4396 9525 4400 9585
rect 4030 9450 4400 9525
rect 4430 9585 4800 9595
rect 4430 9525 4434 9585
rect 4486 9525 4744 9585
rect 4796 9525 4800 9585
rect 4430 9450 4800 9525
rect 4830 9585 5200 9595
rect 4830 9525 4834 9585
rect 4886 9525 5144 9585
rect 5196 9525 5200 9585
rect 4830 9450 5200 9525
rect 5230 9585 5600 9595
rect 5230 9525 5234 9585
rect 5286 9525 5544 9585
rect 5596 9525 5600 9585
rect 5230 9450 5600 9525
rect 5630 9585 6000 9595
rect 5630 9525 5634 9585
rect 5686 9525 5944 9585
rect 5996 9525 6000 9585
rect 5630 9450 6000 9525
rect 2830 9410 6000 9450
rect 2830 9325 3200 9410
rect 2830 9265 2834 9325
rect 2886 9265 3144 9325
rect 3196 9265 3200 9325
rect 2830 9255 3200 9265
rect 3230 9325 3600 9410
rect 3230 9265 3234 9325
rect 3286 9265 3544 9325
rect 3596 9265 3600 9325
rect 3230 9255 3600 9265
rect 3630 9325 4000 9410
rect 3630 9265 3634 9325
rect 3686 9265 3944 9325
rect 3996 9265 4000 9325
rect 3630 9255 4000 9265
rect 4030 9325 4400 9410
rect 4030 9265 4034 9325
rect 4086 9265 4344 9325
rect 4396 9265 4400 9325
rect 4030 9255 4400 9265
rect 4430 9325 4800 9410
rect 4430 9265 4434 9325
rect 4486 9265 4744 9325
rect 4796 9265 4800 9325
rect 4430 9255 4800 9265
rect 4830 9325 5200 9410
rect 4830 9265 4834 9325
rect 4886 9265 5144 9325
rect 5196 9265 5200 9325
rect 4830 9255 5200 9265
rect 5230 9325 5600 9410
rect 5230 9265 5234 9325
rect 5286 9265 5544 9325
rect 5596 9265 5600 9325
rect 5230 9255 5600 9265
rect 5630 9325 6000 9410
rect 5630 9265 5634 9325
rect 5686 9265 5944 9325
rect 5996 9265 6000 9325
rect 5630 9255 6000 9265
rect 6030 9585 6400 9595
rect 6030 9525 6034 9585
rect 6086 9525 6344 9585
rect 6396 9525 6400 9585
rect 6030 9450 6400 9525
rect 6430 9585 6800 9595
rect 6430 9525 6434 9585
rect 6486 9525 6744 9585
rect 6796 9525 6800 9585
rect 6430 9450 6800 9525
rect 6830 9585 7200 9595
rect 6830 9525 6834 9585
rect 6886 9525 7144 9585
rect 7196 9525 7200 9585
rect 6830 9450 7200 9525
rect 7230 9585 7600 9595
rect 7230 9525 7234 9585
rect 7286 9525 7544 9585
rect 7596 9525 7600 9585
rect 7230 9450 7600 9525
rect 6030 9410 7600 9450
rect 6030 9325 6400 9410
rect 6030 9265 6034 9325
rect 6086 9265 6344 9325
rect 6396 9265 6400 9325
rect 6030 9255 6400 9265
rect 6430 9325 6800 9410
rect 6430 9265 6434 9325
rect 6486 9265 6744 9325
rect 6796 9265 6800 9325
rect 6430 9255 6800 9265
rect 6830 9325 7200 9410
rect 6830 9265 6834 9325
rect 6886 9265 7144 9325
rect 7196 9265 7200 9325
rect 6830 9255 7200 9265
rect 7230 9325 7600 9410
rect 7230 9265 7234 9325
rect 7286 9265 7544 9325
rect 7596 9265 7600 9325
rect 7230 9255 7600 9265
rect 7630 9585 8000 9595
rect 7630 9525 7634 9585
rect 7686 9525 7944 9585
rect 7996 9525 8000 9585
rect 7630 9450 8000 9525
rect 8030 9585 8400 9595
rect 8030 9525 8034 9585
rect 8086 9525 8344 9585
rect 8396 9525 8400 9585
rect 8030 9450 8400 9525
rect 7630 9410 8400 9450
rect 7630 9325 8000 9410
rect 7630 9265 7634 9325
rect 7686 9265 7944 9325
rect 7996 9265 8000 9325
rect 7630 9255 8000 9265
rect 8030 9325 8400 9410
rect 8030 9265 8034 9325
rect 8086 9265 8344 9325
rect 8396 9265 8400 9325
rect 8030 9255 8400 9265
rect 8430 9585 8800 9595
rect 8430 9525 8434 9585
rect 8486 9525 8744 9585
rect 8796 9525 8800 9585
rect 8430 9325 8800 9525
rect 8430 9265 8434 9325
rect 8486 9265 8744 9325
rect 8796 9265 8800 9325
rect 8430 9255 8800 9265
rect 8830 9585 9200 9595
rect 8830 9525 8834 9585
rect 8886 9525 9144 9585
rect 9196 9525 9200 9585
rect 8830 9325 9200 9525
rect 8830 9265 8834 9325
rect 8886 9265 9144 9325
rect 9196 9265 9200 9325
rect 8830 9255 9200 9265
rect 9230 9585 9600 9595
rect 9230 9525 9234 9585
rect 9286 9525 9544 9585
rect 9596 9525 9600 9585
rect 9230 9450 9600 9525
rect 9630 9585 10000 9595
rect 9630 9525 9634 9585
rect 9686 9525 9944 9585
rect 9996 9525 10000 9585
rect 9630 9450 10000 9525
rect 10030 9585 10400 9595
rect 10030 9525 10034 9585
rect 10086 9525 10344 9585
rect 10396 9525 10400 9585
rect 10030 9450 10400 9525
rect 10430 9585 10800 9595
rect 10430 9525 10434 9585
rect 10486 9525 10744 9585
rect 10796 9525 10800 9585
rect 10430 9450 10800 9525
rect 10830 9585 11200 9595
rect 10830 9525 10834 9585
rect 10886 9525 11144 9585
rect 11196 9525 11200 9585
rect 10830 9450 11200 9525
rect 11230 9585 11600 9595
rect 11230 9525 11234 9585
rect 11286 9525 11544 9585
rect 11596 9525 11600 9585
rect 11230 9450 11600 9525
rect 11630 9585 12000 9595
rect 11630 9525 11634 9585
rect 11686 9525 11944 9585
rect 11996 9525 12000 9585
rect 11630 9450 12000 9525
rect 12030 9585 12400 9595
rect 12030 9525 12034 9585
rect 12086 9525 12344 9585
rect 12396 9525 12400 9585
rect 12030 9450 12400 9525
rect 12430 9585 12800 9595
rect 12430 9525 12434 9585
rect 12486 9525 12744 9585
rect 12796 9525 12800 9585
rect 12430 9450 12800 9525
rect 12830 9585 13200 9595
rect 12830 9525 12834 9585
rect 12886 9525 13144 9585
rect 13196 9525 13200 9585
rect 12830 9450 13200 9525
rect 9230 9410 13200 9450
rect 9230 9325 9600 9410
rect 9230 9265 9234 9325
rect 9286 9265 9544 9325
rect 9596 9265 9600 9325
rect 9230 9255 9600 9265
rect 9630 9325 10000 9410
rect 9630 9265 9634 9325
rect 9686 9265 9944 9325
rect 9996 9265 10000 9325
rect 9630 9255 10000 9265
rect 10030 9325 10400 9410
rect 10030 9265 10034 9325
rect 10086 9265 10344 9325
rect 10396 9265 10400 9325
rect 10030 9255 10400 9265
rect 10430 9325 10800 9410
rect 10430 9265 10434 9325
rect 10486 9265 10744 9325
rect 10796 9265 10800 9325
rect 10430 9255 10800 9265
rect 10830 9325 11200 9410
rect 10830 9265 10834 9325
rect 10886 9265 11144 9325
rect 11196 9265 11200 9325
rect 10830 9255 11200 9265
rect 11230 9325 11600 9410
rect 11230 9265 11234 9325
rect 11286 9265 11544 9325
rect 11596 9265 11600 9325
rect 11230 9255 11600 9265
rect 11630 9325 12000 9410
rect 11630 9265 11634 9325
rect 11686 9265 11944 9325
rect 11996 9265 12000 9325
rect 11630 9255 12000 9265
rect 12030 9325 12400 9410
rect 12030 9265 12034 9325
rect 12086 9265 12344 9325
rect 12396 9265 12400 9325
rect 12030 9255 12400 9265
rect 12430 9325 12800 9410
rect 12430 9265 12434 9325
rect 12486 9265 12744 9325
rect 12796 9265 12800 9325
rect 12430 9255 12800 9265
rect 12830 9325 13200 9410
rect 12830 9265 12834 9325
rect 12886 9265 13144 9325
rect 13196 9265 13200 9325
rect 12830 9255 13200 9265
rect -330 9225 -324 9255
rect 30 9225 70 9255
rect 430 9225 470 9255
rect 830 9225 870 9255
rect 1230 9225 1270 9255
rect 1630 9225 1670 9255
rect 2030 9225 2070 9255
rect 2430 9225 2470 9255
rect 2830 9225 2870 9255
rect 3230 9225 3270 9255
rect 3630 9225 3670 9255
rect 4030 9225 4070 9255
rect 4430 9225 4470 9255
rect 4830 9225 4870 9255
rect 5230 9225 5270 9255
rect 5630 9225 5670 9255
rect 6030 9225 6070 9255
rect 6430 9225 6470 9255
rect 6830 9225 6870 9255
rect 7230 9225 7270 9255
rect 7630 9225 7670 9255
rect 8030 9225 8070 9255
rect 8430 9225 8470 9255
rect 8830 9225 8870 9255
rect -330 9215 0 9225
rect -314 9155 -56 9215
rect -4 9155 0 9215
rect -330 8955 0 9155
rect -314 8895 -56 8955
rect -4 8895 0 8955
rect -330 8885 0 8895
rect 30 9215 400 9225
rect 30 9155 34 9215
rect 86 9155 344 9215
rect 396 9155 400 9215
rect 30 9080 400 9155
rect 430 9215 800 9225
rect 430 9155 434 9215
rect 486 9155 744 9215
rect 796 9155 800 9215
rect 430 9080 800 9155
rect 830 9215 1200 9225
rect 830 9155 834 9215
rect 886 9155 1144 9215
rect 1196 9155 1200 9215
rect 830 9080 1200 9155
rect 1230 9215 1600 9225
rect 1230 9155 1234 9215
rect 1286 9155 1544 9215
rect 1596 9155 1600 9215
rect 1230 9080 1600 9155
rect 1630 9215 2000 9225
rect 1630 9155 1634 9215
rect 1686 9155 1944 9215
rect 1996 9155 2000 9215
rect 1630 9080 2000 9155
rect 2030 9215 2400 9225
rect 2030 9155 2034 9215
rect 2086 9155 2344 9215
rect 2396 9155 2400 9215
rect 2030 9080 2400 9155
rect 2430 9215 2800 9225
rect 2430 9155 2434 9215
rect 2486 9155 2744 9215
rect 2796 9155 2800 9215
rect 2430 9080 2800 9155
rect 30 9040 2800 9080
rect 30 8955 400 9040
rect 30 8895 34 8955
rect 86 8895 344 8955
rect 396 8895 400 8955
rect 30 8885 400 8895
rect 430 8955 800 9040
rect 430 8895 434 8955
rect 486 8895 744 8955
rect 796 8895 800 8955
rect 430 8885 800 8895
rect 830 8955 1200 9040
rect 830 8895 834 8955
rect 886 8895 1144 8955
rect 1196 8895 1200 8955
rect 830 8885 1200 8895
rect 1230 8955 1600 9040
rect 1230 8895 1234 8955
rect 1286 8895 1544 8955
rect 1596 8895 1600 8955
rect 1230 8885 1600 8895
rect 1630 8955 2000 9040
rect 1630 8895 1634 8955
rect 1686 8895 1944 8955
rect 1996 8895 2000 8955
rect 1630 8885 2000 8895
rect 2030 8955 2400 9040
rect 2030 8895 2034 8955
rect 2086 8895 2344 8955
rect 2396 8895 2400 8955
rect 2030 8885 2400 8895
rect 2430 8955 2800 9040
rect 2430 8895 2434 8955
rect 2486 8895 2744 8955
rect 2796 8895 2800 8955
rect 2430 8885 2800 8895
rect 2830 9215 3200 9225
rect 2830 9155 2834 9215
rect 2886 9155 3144 9215
rect 3196 9155 3200 9215
rect 2830 9080 3200 9155
rect 3230 9215 3600 9225
rect 3230 9155 3234 9215
rect 3286 9155 3544 9215
rect 3596 9155 3600 9215
rect 3230 9080 3600 9155
rect 3630 9215 4000 9225
rect 3630 9155 3634 9215
rect 3686 9155 3944 9215
rect 3996 9155 4000 9215
rect 3630 9080 4000 9155
rect 4030 9215 4400 9225
rect 4030 9155 4034 9215
rect 4086 9155 4344 9215
rect 4396 9155 4400 9215
rect 4030 9080 4400 9155
rect 4430 9215 4800 9225
rect 4430 9155 4434 9215
rect 4486 9155 4744 9215
rect 4796 9155 4800 9215
rect 4430 9080 4800 9155
rect 4830 9215 5200 9225
rect 4830 9155 4834 9215
rect 4886 9155 5144 9215
rect 5196 9155 5200 9215
rect 4830 9080 5200 9155
rect 5230 9215 5600 9225
rect 5230 9155 5234 9215
rect 5286 9155 5544 9215
rect 5596 9155 5600 9215
rect 5230 9080 5600 9155
rect 5630 9215 6000 9225
rect 5630 9155 5634 9215
rect 5686 9155 5944 9215
rect 5996 9155 6000 9215
rect 5630 9080 6000 9155
rect 2830 9040 6000 9080
rect 2830 8955 3200 9040
rect 2830 8895 2834 8955
rect 2886 8895 3144 8955
rect 3196 8895 3200 8955
rect 2830 8885 3200 8895
rect 3230 8955 3600 9040
rect 3230 8895 3234 8955
rect 3286 8895 3544 8955
rect 3596 8895 3600 8955
rect 3230 8885 3600 8895
rect 3630 8955 4000 9040
rect 3630 8895 3634 8955
rect 3686 8895 3944 8955
rect 3996 8895 4000 8955
rect 3630 8885 4000 8895
rect 4030 8955 4400 9040
rect 4030 8895 4034 8955
rect 4086 8895 4344 8955
rect 4396 8895 4400 8955
rect 4030 8885 4400 8895
rect 4430 8955 4800 9040
rect 4430 8895 4434 8955
rect 4486 8895 4744 8955
rect 4796 8895 4800 8955
rect 4430 8885 4800 8895
rect 4830 8955 5200 9040
rect 4830 8895 4834 8955
rect 4886 8895 5144 8955
rect 5196 8895 5200 8955
rect 4830 8885 5200 8895
rect 5230 8955 5600 9040
rect 5230 8895 5234 8955
rect 5286 8895 5544 8955
rect 5596 8895 5600 8955
rect 5230 8885 5600 8895
rect 5630 8955 6000 9040
rect 5630 8895 5634 8955
rect 5686 8895 5944 8955
rect 5996 8895 6000 8955
rect 5630 8885 6000 8895
rect 6030 9215 6400 9225
rect 6030 9155 6034 9215
rect 6086 9155 6344 9215
rect 6396 9155 6400 9215
rect 6030 9080 6400 9155
rect 6430 9215 6800 9225
rect 6430 9155 6434 9215
rect 6486 9155 6744 9215
rect 6796 9155 6800 9215
rect 6430 9080 6800 9155
rect 6830 9215 7200 9225
rect 6830 9155 6834 9215
rect 6886 9155 7144 9215
rect 7196 9155 7200 9215
rect 6830 9080 7200 9155
rect 7230 9215 7600 9225
rect 7230 9155 7234 9215
rect 7286 9155 7544 9215
rect 7596 9155 7600 9215
rect 7230 9080 7600 9155
rect 6030 9040 7600 9080
rect 6030 8955 6400 9040
rect 6030 8895 6034 8955
rect 6086 8895 6344 8955
rect 6396 8895 6400 8955
rect 6030 8885 6400 8895
rect 6430 8955 6800 9040
rect 6430 8895 6434 8955
rect 6486 8895 6744 8955
rect 6796 8895 6800 8955
rect 6430 8885 6800 8895
rect 6830 8955 7200 9040
rect 6830 8895 6834 8955
rect 6886 8895 7144 8955
rect 7196 8895 7200 8955
rect 6830 8885 7200 8895
rect 7230 8955 7600 9040
rect 7230 8895 7234 8955
rect 7286 8895 7544 8955
rect 7596 8895 7600 8955
rect 7230 8885 7600 8895
rect 7630 9215 8000 9225
rect 7630 9155 7634 9215
rect 7686 9155 7944 9215
rect 7996 9155 8000 9215
rect 7630 9080 8000 9155
rect 8030 9215 8400 9225
rect 8030 9155 8034 9215
rect 8086 9155 8344 9215
rect 8396 9155 8400 9215
rect 8030 9080 8400 9155
rect 8430 9215 8800 9225
rect 8430 9155 8434 9215
rect 8486 9155 8744 9215
rect 8796 9155 8800 9215
rect 8430 9080 8800 9155
rect 8830 9215 9200 9225
rect 8830 9155 8834 9215
rect 8886 9155 9144 9215
rect 9196 9155 9200 9215
rect 8830 9080 9200 9155
rect 9230 9215 9600 9225
rect 9230 9155 9234 9215
rect 9286 9155 9544 9215
rect 9596 9155 9600 9215
rect 9230 9080 9600 9155
rect 9630 9215 10000 9225
rect 9630 9155 9634 9215
rect 9686 9155 9944 9215
rect 9996 9155 10000 9215
rect 9630 9080 10000 9155
rect 10030 9215 10400 9225
rect 10030 9155 10034 9215
rect 10086 9155 10344 9215
rect 10396 9155 10400 9215
rect 10030 9080 10400 9155
rect 10430 9215 10800 9225
rect 10430 9155 10434 9215
rect 10486 9155 10744 9215
rect 10796 9155 10800 9215
rect 10430 9080 10800 9155
rect 10830 9215 11200 9225
rect 10830 9155 10834 9215
rect 10886 9155 11144 9215
rect 11196 9155 11200 9215
rect 10830 9080 11200 9155
rect 11230 9215 11600 9225
rect 11230 9155 11234 9215
rect 11286 9155 11544 9215
rect 11596 9155 11600 9215
rect 11230 9080 11600 9155
rect 11630 9215 12000 9225
rect 11630 9155 11634 9215
rect 11686 9155 11944 9215
rect 11996 9155 12000 9215
rect 11630 9080 12000 9155
rect 12030 9215 12400 9225
rect 12030 9155 12034 9215
rect 12086 9155 12344 9215
rect 12396 9155 12400 9215
rect 12030 9080 12400 9155
rect 12430 9215 12800 9225
rect 12430 9155 12434 9215
rect 12486 9155 12744 9215
rect 12796 9155 12800 9215
rect 12430 9080 12800 9155
rect 12830 9215 13200 9225
rect 12830 9155 12834 9215
rect 12886 9155 13144 9215
rect 13196 9155 13200 9215
rect 12830 9080 13200 9155
rect 7630 9040 13390 9080
rect 7630 8955 8000 9040
rect 7630 8895 7634 8955
rect 7686 8895 7944 8955
rect 7996 8895 8000 8955
rect 7630 8885 8000 8895
rect 8030 8955 8400 9040
rect 8030 8895 8034 8955
rect 8086 8895 8344 8955
rect 8396 8895 8400 8955
rect 8030 8885 8400 8895
rect 8430 8955 8800 9040
rect 8430 8895 8434 8955
rect 8486 8895 8744 8955
rect 8796 8895 8800 8955
rect 8430 8885 8800 8895
rect 8830 8955 9200 9040
rect 8830 8895 8834 8955
rect 8886 8895 9144 8955
rect 9196 8895 9200 8955
rect 8830 8885 9200 8895
rect 9230 8955 9600 9040
rect 9230 8895 9234 8955
rect 9286 8895 9544 8955
rect 9596 8895 9600 8955
rect 9230 8885 9600 8895
rect 9630 8955 10000 9040
rect 9630 8895 9634 8955
rect 9686 8895 9944 8955
rect 9996 8895 10000 8955
rect 9630 8885 10000 8895
rect 10030 8955 10400 9040
rect 10030 8895 10034 8955
rect 10086 8895 10344 8955
rect 10396 8895 10400 8955
rect 10030 8885 10400 8895
rect 10430 8955 10800 9040
rect 10430 8895 10434 8955
rect 10486 8895 10744 8955
rect 10796 8895 10800 8955
rect 10430 8885 10800 8895
rect 10830 8955 11200 9040
rect 10830 8895 10834 8955
rect 10886 8895 11144 8955
rect 11196 8895 11200 8955
rect 10830 8885 11200 8895
rect 11230 8955 11600 9040
rect 11230 8895 11234 8955
rect 11286 8895 11544 8955
rect 11596 8895 11600 8955
rect 11230 8885 11600 8895
rect 11630 8955 12000 9040
rect 11630 8895 11634 8955
rect 11686 8895 11944 8955
rect 11996 8895 12000 8955
rect 11630 8885 12000 8895
rect 12030 8955 12400 9040
rect 12030 8895 12034 8955
rect 12086 8895 12344 8955
rect 12396 8895 12400 8955
rect 12030 8885 12400 8895
rect 12430 8955 12800 9040
rect 12430 8895 12434 8955
rect 12486 8895 12744 8955
rect 12796 8895 12800 8955
rect 12430 8885 12800 8895
rect 12830 8955 13200 9040
rect 12830 8895 12834 8955
rect 12886 8895 13144 8955
rect 13196 8895 13200 8955
rect 12830 8885 13200 8895
rect -330 8855 -324 8885
rect 30 8855 70 8885
rect 430 8855 470 8885
rect 830 8855 870 8885
rect 1230 8855 1270 8885
rect 1630 8855 1670 8885
rect 2030 8855 2070 8885
rect 2430 8855 2470 8885
rect 3230 8855 3270 8885
rect 3630 8855 3670 8885
rect 4030 8855 4070 8885
rect 4430 8855 4470 8885
rect 4830 8855 4870 8885
rect 5230 8855 5270 8885
rect 5630 8855 5670 8885
rect 6030 8855 6070 8885
rect 6430 8855 6470 8885
rect 6830 8855 6870 8885
rect 7230 8855 7270 8885
rect 8030 8855 8070 8885
rect 8430 8855 8470 8885
rect 8830 8855 8870 8885
rect 9230 8855 9270 8885
rect 9630 8855 9670 8885
rect 10030 8855 10070 8885
rect 10430 8855 10470 8885
rect 10830 8855 10870 8885
rect 11230 8855 11270 8885
rect 11630 8855 11670 8885
rect 12030 8855 12070 8885
rect 12430 8855 12470 8885
rect -330 8845 0 8855
rect -314 8785 -56 8845
rect -4 8785 0 8845
rect -330 8585 0 8785
rect -314 8525 -56 8585
rect -4 8525 0 8585
rect -330 8515 0 8525
rect 30 8845 400 8855
rect 30 8785 34 8845
rect 86 8785 344 8845
rect 396 8785 400 8845
rect 30 8710 400 8785
rect 430 8845 800 8855
rect 430 8785 434 8845
rect 486 8785 744 8845
rect 796 8785 800 8845
rect 430 8710 800 8785
rect 830 8845 1200 8855
rect 830 8785 834 8845
rect 886 8785 1144 8845
rect 1196 8785 1200 8845
rect 830 8710 1200 8785
rect 1230 8845 1600 8855
rect 1230 8785 1234 8845
rect 1286 8785 1544 8845
rect 1596 8785 1600 8845
rect 1230 8710 1600 8785
rect 1630 8845 2000 8855
rect 1630 8785 1634 8845
rect 1686 8785 1944 8845
rect 1996 8785 2000 8845
rect 1630 8710 2000 8785
rect 2030 8845 2400 8855
rect 2030 8785 2034 8845
rect 2086 8785 2344 8845
rect 2396 8785 2400 8845
rect 2030 8710 2400 8785
rect 2430 8845 2800 8855
rect 2430 8785 2434 8845
rect 2486 8785 2744 8845
rect 2796 8785 2800 8845
rect 2430 8710 2800 8785
rect 2830 8845 3200 8855
rect 2830 8785 2834 8845
rect 2886 8785 3144 8845
rect 3196 8785 3200 8845
rect 2830 8710 3200 8785
rect 30 8670 3200 8710
rect 30 8585 400 8670
rect 30 8525 34 8585
rect 86 8525 344 8585
rect 396 8525 400 8585
rect 30 8515 400 8525
rect 430 8585 800 8670
rect 430 8525 434 8585
rect 486 8525 744 8585
rect 796 8525 800 8585
rect 430 8515 800 8525
rect 830 8585 1200 8670
rect 830 8525 834 8585
rect 886 8525 1144 8585
rect 1196 8525 1200 8585
rect 830 8515 1200 8525
rect 1230 8585 1600 8670
rect 1230 8525 1234 8585
rect 1286 8525 1544 8585
rect 1596 8525 1600 8585
rect 1230 8515 1600 8525
rect 1630 8585 2000 8670
rect 1630 8525 1634 8585
rect 1686 8525 1944 8585
rect 1996 8525 2000 8585
rect 1630 8515 2000 8525
rect 2030 8585 2400 8670
rect 2030 8525 2034 8585
rect 2086 8525 2344 8585
rect 2396 8525 2400 8585
rect 2030 8515 2400 8525
rect 2430 8585 2800 8670
rect 2430 8525 2434 8585
rect 2486 8525 2744 8585
rect 2796 8525 2800 8585
rect 2430 8515 2800 8525
rect 2830 8585 3200 8670
rect 2830 8525 2834 8585
rect 2886 8525 3144 8585
rect 3196 8525 3200 8585
rect 2830 8515 3200 8525
rect 3230 8845 3600 8855
rect 3230 8785 3234 8845
rect 3286 8785 3544 8845
rect 3596 8785 3600 8845
rect 3230 8710 3600 8785
rect 3630 8845 4000 8855
rect 3630 8785 3634 8845
rect 3686 8785 3944 8845
rect 3996 8785 4000 8845
rect 3630 8710 4000 8785
rect 4030 8845 4400 8855
rect 4030 8785 4034 8845
rect 4086 8785 4344 8845
rect 4396 8785 4400 8845
rect 4030 8710 4400 8785
rect 4430 8845 4800 8855
rect 4430 8785 4434 8845
rect 4486 8785 4744 8845
rect 4796 8785 4800 8845
rect 4430 8710 4800 8785
rect 4830 8845 5200 8855
rect 4830 8785 4834 8845
rect 4886 8785 5144 8845
rect 5196 8785 5200 8845
rect 4830 8710 5200 8785
rect 5230 8845 5600 8855
rect 5230 8785 5234 8845
rect 5286 8785 5544 8845
rect 5596 8785 5600 8845
rect 5230 8710 5600 8785
rect 5630 8845 6000 8855
rect 5630 8785 5634 8845
rect 5686 8785 5944 8845
rect 5996 8785 6000 8845
rect 5630 8710 6000 8785
rect 3230 8670 6000 8710
rect 3230 8585 3600 8670
rect 3230 8525 3234 8585
rect 3286 8525 3544 8585
rect 3596 8525 3600 8585
rect 3230 8515 3600 8525
rect 3630 8585 4000 8670
rect 3630 8525 3634 8585
rect 3686 8525 3944 8585
rect 3996 8525 4000 8585
rect 3630 8515 4000 8525
rect 4030 8585 4400 8670
rect 4030 8525 4034 8585
rect 4086 8525 4344 8585
rect 4396 8525 4400 8585
rect 4030 8515 4400 8525
rect 4430 8585 4800 8670
rect 4430 8525 4434 8585
rect 4486 8525 4744 8585
rect 4796 8525 4800 8585
rect 4430 8515 4800 8525
rect 4830 8585 5200 8670
rect 4830 8525 4834 8585
rect 4886 8525 5144 8585
rect 5196 8525 5200 8585
rect 4830 8515 5200 8525
rect 5230 8585 5600 8670
rect 5230 8525 5234 8585
rect 5286 8525 5544 8585
rect 5596 8525 5600 8585
rect 5230 8515 5600 8525
rect 5630 8585 6000 8670
rect 5630 8525 5634 8585
rect 5686 8525 5944 8585
rect 5996 8525 6000 8585
rect 5630 8515 6000 8525
rect 6030 8845 6400 8855
rect 6030 8785 6034 8845
rect 6086 8785 6344 8845
rect 6396 8785 6400 8845
rect 6030 8710 6400 8785
rect 6430 8845 6800 8855
rect 6430 8785 6434 8845
rect 6486 8785 6744 8845
rect 6796 8785 6800 8845
rect 6430 8710 6800 8785
rect 6830 8845 7200 8855
rect 6830 8785 6834 8845
rect 6886 8785 7144 8845
rect 7196 8785 7200 8845
rect 6830 8710 7200 8785
rect 7230 8845 7600 8855
rect 7230 8785 7234 8845
rect 7286 8785 7544 8845
rect 7596 8785 7600 8845
rect 7230 8710 7600 8785
rect 7630 8845 8000 8855
rect 7630 8785 7634 8845
rect 7686 8785 7944 8845
rect 7996 8785 8000 8845
rect 7630 8710 8000 8785
rect 6030 8670 8000 8710
rect 6030 8585 6400 8670
rect 6030 8525 6034 8585
rect 6086 8525 6344 8585
rect 6396 8525 6400 8585
rect 6030 8515 6400 8525
rect 6430 8585 6800 8670
rect 6430 8525 6434 8585
rect 6486 8525 6744 8585
rect 6796 8525 6800 8585
rect 6430 8515 6800 8525
rect 6830 8585 7200 8670
rect 6830 8525 6834 8585
rect 6886 8525 7144 8585
rect 7196 8525 7200 8585
rect 6830 8515 7200 8525
rect 7230 8585 7600 8670
rect 7230 8525 7234 8585
rect 7286 8525 7544 8585
rect 7596 8525 7600 8585
rect 7230 8515 7600 8525
rect 7630 8585 8000 8670
rect 7630 8525 7634 8585
rect 7686 8525 7944 8585
rect 7996 8525 8000 8585
rect 7630 8515 8000 8525
rect 8030 8845 8400 8855
rect 8030 8785 8034 8845
rect 8086 8785 8344 8845
rect 8396 8785 8400 8845
rect 8030 8710 8400 8785
rect 8430 8845 8800 8855
rect 8430 8785 8434 8845
rect 8486 8785 8744 8845
rect 8796 8785 8800 8845
rect 8430 8710 8800 8785
rect 8830 8845 9200 8855
rect 8830 8785 8834 8845
rect 8886 8785 9144 8845
rect 9196 8785 9200 8845
rect 8830 8710 9200 8785
rect 9230 8845 9600 8855
rect 9230 8785 9234 8845
rect 9286 8785 9544 8845
rect 9596 8785 9600 8845
rect 9230 8710 9600 8785
rect 9630 8845 10000 8855
rect 9630 8785 9634 8845
rect 9686 8785 9944 8845
rect 9996 8785 10000 8845
rect 9630 8710 10000 8785
rect 10030 8845 10400 8855
rect 10030 8785 10034 8845
rect 10086 8785 10344 8845
rect 10396 8785 10400 8845
rect 10030 8710 10400 8785
rect 10430 8845 10800 8855
rect 10430 8785 10434 8845
rect 10486 8785 10744 8845
rect 10796 8785 10800 8845
rect 10430 8710 10800 8785
rect 10830 8845 11200 8855
rect 10830 8785 10834 8845
rect 10886 8785 11144 8845
rect 11196 8785 11200 8845
rect 10830 8710 11200 8785
rect 11230 8845 11600 8855
rect 11230 8785 11234 8845
rect 11286 8785 11544 8845
rect 11596 8785 11600 8845
rect 11230 8710 11600 8785
rect 11630 8845 12000 8855
rect 11630 8785 11634 8845
rect 11686 8785 11944 8845
rect 11996 8785 12000 8845
rect 11630 8710 12000 8785
rect 12030 8845 12400 8855
rect 12030 8785 12034 8845
rect 12086 8785 12344 8845
rect 12396 8785 12400 8845
rect 12030 8710 12400 8785
rect 12430 8845 12800 8855
rect 12430 8785 12434 8845
rect 12486 8785 12744 8845
rect 12796 8785 12800 8845
rect 12430 8710 12800 8785
rect 12830 8845 13200 8855
rect 12830 8785 12834 8845
rect 12886 8785 13144 8845
rect 13196 8785 13200 8845
rect 12830 8710 13200 8785
rect 8030 8670 13200 8710
rect 8030 8585 8400 8670
rect 8030 8525 8034 8585
rect 8086 8525 8344 8585
rect 8396 8525 8400 8585
rect 8030 8515 8400 8525
rect 8430 8585 8800 8670
rect 8430 8525 8434 8585
rect 8486 8525 8744 8585
rect 8796 8525 8800 8585
rect 8430 8515 8800 8525
rect 8830 8585 9200 8670
rect 8830 8525 8834 8585
rect 8886 8525 9144 8585
rect 9196 8525 9200 8585
rect 8830 8515 9200 8525
rect 9230 8585 9600 8670
rect 9230 8525 9234 8585
rect 9286 8525 9544 8585
rect 9596 8525 9600 8585
rect 9230 8515 9600 8525
rect 9630 8585 10000 8670
rect 9630 8525 9634 8585
rect 9686 8525 9944 8585
rect 9996 8525 10000 8585
rect 9630 8515 10000 8525
rect 10030 8585 10400 8670
rect 10030 8525 10034 8585
rect 10086 8525 10344 8585
rect 10396 8525 10400 8585
rect 10030 8515 10400 8525
rect 10430 8585 10800 8670
rect 10430 8525 10434 8585
rect 10486 8525 10744 8585
rect 10796 8525 10800 8585
rect 10430 8515 10800 8525
rect 10830 8585 11200 8670
rect 10830 8525 10834 8585
rect 10886 8525 11144 8585
rect 11196 8525 11200 8585
rect 10830 8515 11200 8525
rect 11230 8585 11600 8670
rect 11230 8525 11234 8585
rect 11286 8525 11544 8585
rect 11596 8525 11600 8585
rect 11230 8515 11600 8525
rect 11630 8585 12000 8670
rect 11630 8525 11634 8585
rect 11686 8525 11944 8585
rect 11996 8525 12000 8585
rect 11630 8515 12000 8525
rect 12030 8585 12400 8670
rect 12030 8525 12034 8585
rect 12086 8525 12344 8585
rect 12396 8525 12400 8585
rect 12030 8515 12400 8525
rect 12430 8585 12800 8670
rect 12430 8525 12434 8585
rect 12486 8525 12744 8585
rect 12796 8525 12800 8585
rect 12430 8515 12800 8525
rect 12830 8585 13200 8670
rect 12830 8525 12834 8585
rect 12886 8525 13144 8585
rect 13196 8525 13200 8585
rect 12830 8515 13200 8525
rect -330 8485 -324 8515
rect 30 8485 70 8515
rect 430 8485 470 8515
rect 830 8485 870 8515
rect 1230 8485 1270 8515
rect 1630 8485 1670 8515
rect 2030 8485 2070 8515
rect 2430 8485 2470 8515
rect 2830 8485 2870 8515
rect 3230 8485 3270 8515
rect 3630 8485 3670 8515
rect 4030 8485 4070 8515
rect 4430 8485 4470 8515
rect 4830 8485 4870 8515
rect 5230 8485 5270 8515
rect 5630 8485 5670 8515
rect 6030 8485 6070 8515
rect 6430 8485 6470 8515
rect 6830 8485 6870 8515
rect 7230 8485 7270 8515
rect 7630 8485 7670 8515
rect 8030 8485 8070 8515
rect 8430 8485 8470 8515
rect 8830 8485 8870 8515
rect 9230 8485 9270 8515
rect 9630 8485 9670 8515
rect 10030 8485 10070 8515
rect 10430 8485 10470 8515
rect 10830 8485 10870 8515
rect 11230 8485 11270 8515
rect 11630 8485 11670 8515
rect 12030 8485 12070 8515
rect 12430 8485 12470 8515
rect -330 8475 0 8485
rect -314 8415 -56 8475
rect -4 8415 0 8475
rect -330 8215 0 8415
rect -314 8155 -56 8215
rect -4 8155 0 8215
rect -330 8145 0 8155
rect 30 8475 400 8485
rect 30 8415 34 8475
rect 86 8415 344 8475
rect 396 8415 400 8475
rect 30 8340 400 8415
rect 430 8475 800 8485
rect 430 8415 434 8475
rect 486 8415 744 8475
rect 796 8415 800 8475
rect 430 8340 800 8415
rect 830 8475 1200 8485
rect 830 8415 834 8475
rect 886 8415 1144 8475
rect 1196 8415 1200 8475
rect 830 8340 1200 8415
rect 1230 8475 1600 8485
rect 1230 8415 1234 8475
rect 1286 8415 1544 8475
rect 1596 8415 1600 8475
rect 1230 8340 1600 8415
rect 1630 8475 2000 8485
rect 1630 8415 1634 8475
rect 1686 8415 1944 8475
rect 1996 8415 2000 8475
rect 1630 8340 2000 8415
rect 2030 8475 2400 8485
rect 2030 8415 2034 8475
rect 2086 8415 2344 8475
rect 2396 8415 2400 8475
rect 2030 8340 2400 8415
rect 2430 8475 2800 8485
rect 2430 8415 2434 8475
rect 2486 8415 2744 8475
rect 2796 8415 2800 8475
rect 2430 8340 2800 8415
rect 2830 8475 3200 8485
rect 2830 8415 2834 8475
rect 2886 8415 3144 8475
rect 3196 8415 3200 8475
rect 2830 8340 3200 8415
rect 30 8300 3200 8340
rect 30 8215 400 8300
rect 30 8155 34 8215
rect 86 8155 344 8215
rect 396 8155 400 8215
rect 30 8145 400 8155
rect 430 8215 800 8300
rect 430 8155 434 8215
rect 486 8155 744 8215
rect 796 8155 800 8215
rect 430 8145 800 8155
rect 830 8215 1200 8300
rect 830 8155 834 8215
rect 886 8155 1144 8215
rect 1196 8155 1200 8215
rect 830 8145 1200 8155
rect 1230 8215 1600 8300
rect 1230 8155 1234 8215
rect 1286 8155 1544 8215
rect 1596 8155 1600 8215
rect 1230 8145 1600 8155
rect 1630 8215 2000 8300
rect 1630 8155 1634 8215
rect 1686 8155 1944 8215
rect 1996 8155 2000 8215
rect 1630 8145 2000 8155
rect 2030 8215 2400 8300
rect 2030 8155 2034 8215
rect 2086 8155 2344 8215
rect 2396 8155 2400 8215
rect 2030 8145 2400 8155
rect 2430 8215 2800 8300
rect 2430 8155 2434 8215
rect 2486 8155 2744 8215
rect 2796 8155 2800 8215
rect 2430 8145 2800 8155
rect 2830 8215 3200 8300
rect 2830 8155 2834 8215
rect 2886 8155 3144 8215
rect 3196 8155 3200 8215
rect 2830 8145 3200 8155
rect 3230 8475 3600 8485
rect 3230 8415 3234 8475
rect 3286 8415 3544 8475
rect 3596 8415 3600 8475
rect 3230 8340 3600 8415
rect 3630 8475 4000 8485
rect 3630 8415 3634 8475
rect 3686 8415 3944 8475
rect 3996 8415 4000 8475
rect 3630 8340 4000 8415
rect 4030 8475 4400 8485
rect 4030 8415 4034 8475
rect 4086 8415 4344 8475
rect 4396 8415 4400 8475
rect 4030 8340 4400 8415
rect 4430 8475 4800 8485
rect 4430 8415 4434 8475
rect 4486 8415 4744 8475
rect 4796 8415 4800 8475
rect 4430 8340 4800 8415
rect 4830 8475 5200 8485
rect 4830 8415 4834 8475
rect 4886 8415 5144 8475
rect 5196 8415 5200 8475
rect 4830 8340 5200 8415
rect 5230 8475 5600 8485
rect 5230 8415 5234 8475
rect 5286 8415 5544 8475
rect 5596 8415 5600 8475
rect 5230 8340 5600 8415
rect 5630 8475 6000 8485
rect 5630 8415 5634 8475
rect 5686 8415 5944 8475
rect 5996 8415 6000 8475
rect 5630 8340 6000 8415
rect 3230 8300 6000 8340
rect 3230 8215 3600 8300
rect 3230 8155 3234 8215
rect 3286 8155 3544 8215
rect 3596 8155 3600 8215
rect 3230 8145 3600 8155
rect 3630 8215 4000 8300
rect 3630 8155 3634 8215
rect 3686 8155 3944 8215
rect 3996 8155 4000 8215
rect 3630 8145 4000 8155
rect 4030 8215 4400 8300
rect 4030 8155 4034 8215
rect 4086 8155 4344 8215
rect 4396 8155 4400 8215
rect 4030 8145 4400 8155
rect 4430 8215 4800 8300
rect 4430 8155 4434 8215
rect 4486 8155 4744 8215
rect 4796 8155 4800 8215
rect 4430 8145 4800 8155
rect 4830 8215 5200 8300
rect 4830 8155 4834 8215
rect 4886 8155 5144 8215
rect 5196 8155 5200 8215
rect 4830 8145 5200 8155
rect 5230 8215 5600 8300
rect 5230 8155 5234 8215
rect 5286 8155 5544 8215
rect 5596 8155 5600 8215
rect 5230 8145 5600 8155
rect 5630 8215 6000 8300
rect 5630 8155 5634 8215
rect 5686 8155 5944 8215
rect 5996 8155 6000 8215
rect 5630 8145 6000 8155
rect 6030 8475 6400 8485
rect 6030 8415 6034 8475
rect 6086 8415 6344 8475
rect 6396 8415 6400 8475
rect 6030 8340 6400 8415
rect 6430 8475 6800 8485
rect 6430 8415 6434 8475
rect 6486 8415 6744 8475
rect 6796 8415 6800 8475
rect 6430 8340 6800 8415
rect 6830 8475 7200 8485
rect 6830 8415 6834 8475
rect 6886 8415 7144 8475
rect 7196 8415 7200 8475
rect 6830 8340 7200 8415
rect 7230 8475 7600 8485
rect 7230 8415 7234 8475
rect 7286 8415 7544 8475
rect 7596 8415 7600 8475
rect 7230 8340 7600 8415
rect 7630 8475 8000 8485
rect 7630 8415 7634 8475
rect 7686 8415 7944 8475
rect 7996 8415 8000 8475
rect 7630 8340 8000 8415
rect 6030 8300 8000 8340
rect 6030 8215 6400 8300
rect 6030 8155 6034 8215
rect 6086 8155 6344 8215
rect 6396 8155 6400 8215
rect 6030 8145 6400 8155
rect 6430 8215 6800 8300
rect 6430 8155 6434 8215
rect 6486 8155 6744 8215
rect 6796 8155 6800 8215
rect 6430 8145 6800 8155
rect 6830 8215 7200 8300
rect 6830 8155 6834 8215
rect 6886 8155 7144 8215
rect 7196 8155 7200 8215
rect 6830 8145 7200 8155
rect 7230 8215 7600 8300
rect 7230 8155 7234 8215
rect 7286 8155 7544 8215
rect 7596 8155 7600 8215
rect 7230 8145 7600 8155
rect 7630 8215 8000 8300
rect 7630 8155 7634 8215
rect 7686 8155 7944 8215
rect 7996 8155 8000 8215
rect 7630 8145 8000 8155
rect 8030 8475 8400 8485
rect 8030 8415 8034 8475
rect 8086 8415 8344 8475
rect 8396 8415 8400 8475
rect 8030 8340 8400 8415
rect 8430 8475 8800 8485
rect 8430 8415 8434 8475
rect 8486 8415 8744 8475
rect 8796 8415 8800 8475
rect 8430 8340 8800 8415
rect 8830 8475 9200 8485
rect 8830 8415 8834 8475
rect 8886 8415 9144 8475
rect 9196 8415 9200 8475
rect 8830 8340 9200 8415
rect 9230 8475 9600 8485
rect 9230 8415 9234 8475
rect 9286 8415 9544 8475
rect 9596 8415 9600 8475
rect 9230 8340 9600 8415
rect 9630 8475 10000 8485
rect 9630 8415 9634 8475
rect 9686 8415 9944 8475
rect 9996 8415 10000 8475
rect 9630 8340 10000 8415
rect 10030 8475 10400 8485
rect 10030 8415 10034 8475
rect 10086 8415 10344 8475
rect 10396 8415 10400 8475
rect 10030 8340 10400 8415
rect 10430 8475 10800 8485
rect 10430 8415 10434 8475
rect 10486 8415 10744 8475
rect 10796 8415 10800 8475
rect 10430 8340 10800 8415
rect 10830 8475 11200 8485
rect 10830 8415 10834 8475
rect 10886 8415 11144 8475
rect 11196 8415 11200 8475
rect 10830 8340 11200 8415
rect 11230 8475 11600 8485
rect 11230 8415 11234 8475
rect 11286 8415 11544 8475
rect 11596 8415 11600 8475
rect 11230 8340 11600 8415
rect 11630 8475 12000 8485
rect 11630 8415 11634 8475
rect 11686 8415 11944 8475
rect 11996 8415 12000 8475
rect 11630 8340 12000 8415
rect 12030 8475 12400 8485
rect 12030 8415 12034 8475
rect 12086 8415 12344 8475
rect 12396 8415 12400 8475
rect 12030 8340 12400 8415
rect 12430 8475 12800 8485
rect 12430 8415 12434 8475
rect 12486 8415 12744 8475
rect 12796 8415 12800 8475
rect 12430 8340 12800 8415
rect 12830 8475 13200 8485
rect 12830 8415 12834 8475
rect 12886 8415 13144 8475
rect 13196 8415 13200 8475
rect 12830 8340 13200 8415
rect 8030 8300 13200 8340
rect 8030 8215 8400 8300
rect 8030 8155 8034 8215
rect 8086 8155 8344 8215
rect 8396 8155 8400 8215
rect 8030 8145 8400 8155
rect 8430 8215 8800 8300
rect 8430 8155 8434 8215
rect 8486 8155 8744 8215
rect 8796 8155 8800 8215
rect 8430 8145 8800 8155
rect 8830 8215 9200 8300
rect 8830 8155 8834 8215
rect 8886 8155 9144 8215
rect 9196 8155 9200 8215
rect 8830 8145 9200 8155
rect 9230 8215 9600 8300
rect 9230 8155 9234 8215
rect 9286 8155 9544 8215
rect 9596 8155 9600 8215
rect 9230 8145 9600 8155
rect 9630 8215 10000 8300
rect 9630 8155 9634 8215
rect 9686 8155 9944 8215
rect 9996 8155 10000 8215
rect 9630 8145 10000 8155
rect 10030 8215 10400 8300
rect 10030 8155 10034 8215
rect 10086 8155 10344 8215
rect 10396 8155 10400 8215
rect 10030 8145 10400 8155
rect 10430 8215 10800 8300
rect 10430 8155 10434 8215
rect 10486 8155 10744 8215
rect 10796 8155 10800 8215
rect 10430 8145 10800 8155
rect 10830 8215 11200 8300
rect 10830 8155 10834 8215
rect 10886 8155 11144 8215
rect 11196 8155 11200 8215
rect 10830 8145 11200 8155
rect 11230 8215 11600 8300
rect 11230 8155 11234 8215
rect 11286 8155 11544 8215
rect 11596 8155 11600 8215
rect 11230 8145 11600 8155
rect 11630 8215 12000 8300
rect 11630 8155 11634 8215
rect 11686 8155 11944 8215
rect 11996 8155 12000 8215
rect 11630 8145 12000 8155
rect 12030 8215 12400 8300
rect 12030 8155 12034 8215
rect 12086 8155 12344 8215
rect 12396 8155 12400 8215
rect 12030 8145 12400 8155
rect 12430 8215 12800 8300
rect 12430 8155 12434 8215
rect 12486 8155 12744 8215
rect 12796 8155 12800 8215
rect 12430 8145 12800 8155
rect 12830 8215 13200 8300
rect 12830 8155 12834 8215
rect 12886 8155 13144 8215
rect 13196 8155 13200 8215
rect 12830 8145 13200 8155
rect -330 8115 -324 8145
rect 30 8115 70 8145
rect 430 8115 470 8145
rect 830 8115 870 8145
rect 1230 8115 1270 8145
rect 1630 8115 1670 8145
rect 2030 8115 2070 8145
rect 2430 8115 2470 8145
rect 2830 8115 2870 8145
rect 3230 8115 3270 8145
rect 3630 8115 3670 8145
rect 4030 8115 4070 8145
rect 4430 8115 4470 8145
rect 4830 8115 4870 8145
rect 5230 8115 5270 8145
rect 5630 8115 5670 8145
rect 6030 8115 6070 8145
rect 6430 8115 6470 8145
rect 6830 8115 6870 8145
rect 7230 8115 7270 8145
rect 7630 8115 7670 8145
rect -330 8105 0 8115
rect -314 8045 -56 8105
rect -4 8045 0 8105
rect -330 7845 0 8045
rect -314 7785 -56 7845
rect -4 7785 0 7845
rect -330 7775 0 7785
rect 30 8105 400 8115
rect 30 8045 34 8105
rect 86 8045 344 8105
rect 396 8045 400 8105
rect 30 7970 400 8045
rect 430 8105 800 8115
rect 430 8045 434 8105
rect 486 8045 744 8105
rect 796 8045 800 8105
rect 430 7970 800 8045
rect 830 8105 1200 8115
rect 830 8045 834 8105
rect 886 8045 1144 8105
rect 1196 8045 1200 8105
rect 830 7970 1200 8045
rect 1230 8105 1600 8115
rect 1230 8045 1234 8105
rect 1286 8045 1544 8105
rect 1596 8045 1600 8105
rect 1230 7970 1600 8045
rect 1630 8105 2000 8115
rect 1630 8045 1634 8105
rect 1686 8045 1944 8105
rect 1996 8045 2000 8105
rect 1630 7970 2000 8045
rect 2030 8105 2400 8115
rect 2030 8045 2034 8105
rect 2086 8045 2344 8105
rect 2396 8045 2400 8105
rect 2030 7970 2400 8045
rect 2430 8105 2800 8115
rect 2430 8045 2434 8105
rect 2486 8045 2744 8105
rect 2796 8045 2800 8105
rect 2430 7970 2800 8045
rect 2830 8105 3200 8115
rect 2830 8045 2834 8105
rect 2886 8045 3144 8105
rect 3196 8045 3200 8105
rect 2830 7970 3200 8045
rect 30 7930 3200 7970
rect 30 7845 400 7930
rect 30 7785 34 7845
rect 86 7785 344 7845
rect 396 7785 400 7845
rect 30 7775 400 7785
rect 430 7845 800 7930
rect 430 7785 434 7845
rect 486 7785 744 7845
rect 796 7785 800 7845
rect 430 7775 800 7785
rect 830 7845 1200 7930
rect 830 7785 834 7845
rect 886 7785 1144 7845
rect 1196 7785 1200 7845
rect 830 7775 1200 7785
rect 1230 7845 1600 7930
rect 1230 7785 1234 7845
rect 1286 7785 1544 7845
rect 1596 7785 1600 7845
rect 1230 7775 1600 7785
rect 1630 7845 2000 7930
rect 1630 7785 1634 7845
rect 1686 7785 1944 7845
rect 1996 7785 2000 7845
rect 1630 7775 2000 7785
rect 2030 7845 2400 7930
rect 2030 7785 2034 7845
rect 2086 7785 2344 7845
rect 2396 7785 2400 7845
rect 2030 7775 2400 7785
rect 2430 7845 2800 7930
rect 2430 7785 2434 7845
rect 2486 7785 2744 7845
rect 2796 7785 2800 7845
rect 2430 7775 2800 7785
rect 2830 7845 3200 7930
rect 2830 7785 2834 7845
rect 2886 7785 3144 7845
rect 3196 7785 3200 7845
rect 2830 7775 3200 7785
rect 3230 8105 3600 8115
rect 3230 8045 3234 8105
rect 3286 8045 3544 8105
rect 3596 8045 3600 8105
rect 3230 7970 3600 8045
rect 3630 8105 4000 8115
rect 3630 8045 3634 8105
rect 3686 8045 3944 8105
rect 3996 8045 4000 8105
rect 3630 7970 4000 8045
rect 4030 8105 4400 8115
rect 4030 8045 4034 8105
rect 4086 8045 4344 8105
rect 4396 8045 4400 8105
rect 4030 7970 4400 8045
rect 4430 8105 4800 8115
rect 4430 8045 4434 8105
rect 4486 8045 4744 8105
rect 4796 8045 4800 8105
rect 4430 7970 4800 8045
rect 4830 8105 5200 8115
rect 4830 8045 4834 8105
rect 4886 8045 5144 8105
rect 5196 8045 5200 8105
rect 4830 7970 5200 8045
rect 5230 8105 5600 8115
rect 5230 8045 5234 8105
rect 5286 8045 5544 8105
rect 5596 8045 5600 8105
rect 5230 7970 5600 8045
rect 5630 8105 6000 8115
rect 5630 8045 5634 8105
rect 5686 8045 5944 8105
rect 5996 8045 6000 8105
rect 5630 7970 6000 8045
rect 3230 7930 6000 7970
rect 3230 7845 3600 7930
rect 3230 7785 3234 7845
rect 3286 7785 3544 7845
rect 3596 7785 3600 7845
rect 3230 7775 3600 7785
rect 3630 7845 4000 7930
rect 3630 7785 3634 7845
rect 3686 7785 3944 7845
rect 3996 7785 4000 7845
rect 3630 7775 4000 7785
rect 4030 7845 4400 7930
rect 4030 7785 4034 7845
rect 4086 7785 4344 7845
rect 4396 7785 4400 7845
rect 4030 7775 4400 7785
rect 4430 7845 4800 7930
rect 4430 7785 4434 7845
rect 4486 7785 4744 7845
rect 4796 7785 4800 7845
rect 4430 7775 4800 7785
rect 4830 7845 5200 7930
rect 4830 7785 4834 7845
rect 4886 7785 5144 7845
rect 5196 7785 5200 7845
rect 4830 7775 5200 7785
rect 5230 7845 5600 7930
rect 5230 7785 5234 7845
rect 5286 7785 5544 7845
rect 5596 7785 5600 7845
rect 5230 7775 5600 7785
rect 5630 7845 6000 7930
rect 5630 7785 5634 7845
rect 5686 7785 5944 7845
rect 5996 7785 6000 7845
rect 5630 7775 6000 7785
rect 6030 8105 6400 8115
rect 6030 8045 6034 8105
rect 6086 8045 6344 8105
rect 6396 8045 6400 8105
rect 6030 7970 6400 8045
rect 6430 8105 6800 8115
rect 6430 8045 6434 8105
rect 6486 8045 6744 8105
rect 6796 8045 6800 8105
rect 6430 7970 6800 8045
rect 6830 8105 7200 8115
rect 6830 8045 6834 8105
rect 6886 8045 7144 8105
rect 7196 8045 7200 8105
rect 6830 7970 7200 8045
rect 7230 8105 7600 8115
rect 7230 8045 7234 8105
rect 7286 8045 7544 8105
rect 7596 8045 7600 8105
rect 7230 7970 7600 8045
rect 7630 8105 8000 8115
rect 7630 8045 7634 8105
rect 7686 8045 7944 8105
rect 7996 8045 8000 8105
rect 7630 7970 8000 8045
rect 8030 8105 8400 8115
rect 8030 8045 8034 8105
rect 8086 8045 8344 8105
rect 8396 8045 8400 8105
rect 8030 7970 8400 8045
rect 8430 8105 8800 8115
rect 8430 8045 8434 8105
rect 8486 8045 8744 8105
rect 8796 8045 8800 8105
rect 8430 7970 8800 8045
rect 8830 8105 9200 8115
rect 8830 8045 8834 8105
rect 8886 8045 9144 8105
rect 9196 8045 9200 8105
rect 8830 7970 9200 8045
rect 9230 8105 9600 8115
rect 9230 8045 9234 8105
rect 9286 8045 9544 8105
rect 9596 8045 9600 8105
rect 9230 7970 9600 8045
rect 9630 8105 10000 8115
rect 9630 8045 9634 8105
rect 9686 8045 9944 8105
rect 9996 8045 10000 8105
rect 9630 7970 10000 8045
rect 10030 8105 10400 8115
rect 10030 8045 10034 8105
rect 10086 8045 10344 8105
rect 10396 8045 10400 8105
rect 10030 7970 10400 8045
rect 10430 8105 10800 8115
rect 10430 8045 10434 8105
rect 10486 8045 10744 8105
rect 10796 8045 10800 8105
rect 10430 7970 10800 8045
rect 10830 8105 11200 8115
rect 10830 8045 10834 8105
rect 10886 8045 11144 8105
rect 11196 8045 11200 8105
rect 10830 7970 11200 8045
rect 11230 8105 11600 8115
rect 11230 8045 11234 8105
rect 11286 8045 11544 8105
rect 11596 8045 11600 8105
rect 11230 7970 11600 8045
rect 11630 8105 12000 8115
rect 11630 8045 11634 8105
rect 11686 8045 11944 8105
rect 11996 8045 12000 8105
rect 11630 7970 12000 8045
rect 12030 8105 12400 8115
rect 12030 8045 12034 8105
rect 12086 8045 12344 8105
rect 12396 8045 12400 8105
rect 12030 7970 12400 8045
rect 12430 8105 12800 8115
rect 12430 8045 12434 8105
rect 12486 8045 12744 8105
rect 12796 8045 12800 8105
rect 12430 7970 12800 8045
rect 12830 8105 13200 8115
rect 12830 8045 12834 8105
rect 12886 8045 13144 8105
rect 13196 8045 13200 8105
rect 12830 7970 13200 8045
rect 6030 7930 13390 7970
rect 6030 7845 6400 7930
rect 6030 7785 6034 7845
rect 6086 7785 6344 7845
rect 6396 7785 6400 7845
rect 6030 7775 6400 7785
rect 6430 7845 6800 7930
rect 6430 7785 6434 7845
rect 6486 7785 6744 7845
rect 6796 7785 6800 7845
rect 6430 7775 6800 7785
rect 6830 7845 7200 7930
rect 6830 7785 6834 7845
rect 6886 7785 7144 7845
rect 7196 7785 7200 7845
rect 6830 7775 7200 7785
rect 7230 7845 7600 7930
rect 7230 7785 7234 7845
rect 7286 7785 7544 7845
rect 7596 7785 7600 7845
rect 7230 7775 7600 7785
rect 7630 7845 8000 7930
rect 7630 7785 7634 7845
rect 7686 7785 7944 7845
rect 7996 7785 8000 7845
rect 7630 7775 8000 7785
rect 8030 7845 8400 7930
rect 8030 7785 8034 7845
rect 8086 7785 8344 7845
rect 8396 7785 8400 7845
rect 8030 7775 8400 7785
rect 8430 7845 8800 7930
rect 8430 7785 8434 7845
rect 8486 7785 8744 7845
rect 8796 7785 8800 7845
rect 8430 7775 8800 7785
rect 8830 7845 9200 7930
rect 8830 7785 8834 7845
rect 8886 7785 9144 7845
rect 9196 7785 9200 7845
rect 8830 7775 9200 7785
rect 9230 7845 9600 7930
rect 9230 7785 9234 7845
rect 9286 7785 9544 7845
rect 9596 7785 9600 7845
rect 9230 7775 9600 7785
rect 9630 7845 10000 7930
rect 9630 7785 9634 7845
rect 9686 7785 9944 7845
rect 9996 7785 10000 7845
rect 9630 7775 10000 7785
rect 10030 7845 10400 7930
rect 10030 7785 10034 7845
rect 10086 7785 10344 7845
rect 10396 7785 10400 7845
rect 10030 7775 10400 7785
rect 10430 7845 10800 7930
rect 10430 7785 10434 7845
rect 10486 7785 10744 7845
rect 10796 7785 10800 7845
rect 10430 7775 10800 7785
rect 10830 7845 11200 7930
rect 10830 7785 10834 7845
rect 10886 7785 11144 7845
rect 11196 7785 11200 7845
rect 10830 7775 11200 7785
rect 11230 7845 11600 7930
rect 11230 7785 11234 7845
rect 11286 7785 11544 7845
rect 11596 7785 11600 7845
rect 11230 7775 11600 7785
rect 11630 7845 12000 7930
rect 11630 7785 11634 7845
rect 11686 7785 11944 7845
rect 11996 7785 12000 7845
rect 11630 7775 12000 7785
rect 12030 7845 12400 7930
rect 12030 7785 12034 7845
rect 12086 7785 12344 7845
rect 12396 7785 12400 7845
rect 12030 7775 12400 7785
rect 12430 7845 12800 7930
rect 12430 7785 12434 7845
rect 12486 7785 12744 7845
rect 12796 7785 12800 7845
rect 12430 7775 12800 7785
rect 12830 7845 13200 7930
rect 12830 7785 12834 7845
rect 12886 7785 13144 7845
rect 13196 7785 13200 7845
rect 12830 7775 13200 7785
rect -330 7745 -324 7775
rect 30 7745 70 7775
rect 430 7745 470 7775
rect 830 7745 870 7775
rect 1230 7745 1270 7775
rect 1630 7745 1670 7775
rect 2030 7745 2070 7775
rect 2430 7745 2470 7775
rect 2830 7745 2870 7775
rect 3230 7745 3270 7775
rect 3630 7745 3670 7775
rect 4030 7745 4070 7775
rect 4430 7745 4470 7775
rect 4830 7745 4870 7775
rect 5230 7745 5270 7775
rect 5630 7745 5670 7775
rect 6030 7745 6070 7775
rect 6430 7745 6470 7775
rect 6830 7745 6870 7775
rect 7230 7745 7270 7775
rect 7630 7745 7670 7775
rect 8030 7745 8070 7775
rect 8430 7745 8470 7775
rect 8830 7745 8870 7775
rect 9230 7745 9270 7775
rect 9630 7745 9670 7775
rect 10030 7745 10070 7775
rect 10430 7745 10470 7775
rect 10830 7745 10870 7775
rect 11230 7745 11270 7775
rect 11630 7745 11670 7775
rect 12030 7745 12070 7775
rect 12430 7745 12470 7775
rect -330 7735 0 7745
rect -314 7675 -56 7735
rect -4 7675 0 7735
rect -330 7475 0 7675
rect -314 7415 -56 7475
rect -4 7415 0 7475
rect -330 7405 0 7415
rect 30 7735 400 7745
rect 30 7675 34 7735
rect 86 7675 344 7735
rect 396 7675 400 7735
rect 30 7600 400 7675
rect 430 7735 800 7745
rect 430 7675 434 7735
rect 486 7675 744 7735
rect 796 7675 800 7735
rect 430 7600 800 7675
rect 830 7735 1200 7745
rect 830 7675 834 7735
rect 886 7675 1144 7735
rect 1196 7675 1200 7735
rect 830 7600 1200 7675
rect 1230 7735 1600 7745
rect 1230 7675 1234 7735
rect 1286 7675 1544 7735
rect 1596 7675 1600 7735
rect 1230 7600 1600 7675
rect 1630 7735 2000 7745
rect 1630 7675 1634 7735
rect 1686 7675 1944 7735
rect 1996 7675 2000 7735
rect 1630 7600 2000 7675
rect 2030 7735 2400 7745
rect 2030 7675 2034 7735
rect 2086 7675 2344 7735
rect 2396 7675 2400 7735
rect 2030 7600 2400 7675
rect 2430 7735 2800 7745
rect 2430 7675 2434 7735
rect 2486 7675 2744 7735
rect 2796 7675 2800 7735
rect 2430 7600 2800 7675
rect 2830 7735 3200 7745
rect 2830 7675 2834 7735
rect 2886 7675 3144 7735
rect 3196 7675 3200 7735
rect 2830 7600 3200 7675
rect 30 7560 3200 7600
rect 30 7475 400 7560
rect 30 7415 34 7475
rect 86 7415 344 7475
rect 396 7415 400 7475
rect 30 7405 400 7415
rect 430 7475 800 7560
rect 430 7415 434 7475
rect 486 7415 744 7475
rect 796 7415 800 7475
rect 430 7405 800 7415
rect 830 7475 1200 7560
rect 830 7415 834 7475
rect 886 7415 1144 7475
rect 1196 7415 1200 7475
rect 830 7405 1200 7415
rect 1230 7475 1600 7560
rect 1230 7415 1234 7475
rect 1286 7415 1544 7475
rect 1596 7415 1600 7475
rect 1230 7405 1600 7415
rect 1630 7475 2000 7560
rect 1630 7415 1634 7475
rect 1686 7415 1944 7475
rect 1996 7415 2000 7475
rect 1630 7405 2000 7415
rect 2030 7475 2400 7560
rect 2030 7415 2034 7475
rect 2086 7415 2344 7475
rect 2396 7415 2400 7475
rect 2030 7405 2400 7415
rect 2430 7475 2800 7560
rect 2430 7415 2434 7475
rect 2486 7415 2744 7475
rect 2796 7415 2800 7475
rect 2430 7405 2800 7415
rect 2830 7475 3200 7560
rect 2830 7415 2834 7475
rect 2886 7415 3144 7475
rect 3196 7415 3200 7475
rect 2830 7405 3200 7415
rect 3230 7735 3600 7745
rect 3230 7675 3234 7735
rect 3286 7675 3544 7735
rect 3596 7675 3600 7735
rect 3230 7600 3600 7675
rect 3630 7735 4000 7745
rect 3630 7675 3634 7735
rect 3686 7675 3944 7735
rect 3996 7675 4000 7735
rect 3630 7600 4000 7675
rect 4030 7735 4400 7745
rect 4030 7675 4034 7735
rect 4086 7675 4344 7735
rect 4396 7675 4400 7735
rect 4030 7600 4400 7675
rect 4430 7735 4800 7745
rect 4430 7675 4434 7735
rect 4486 7675 4744 7735
rect 4796 7675 4800 7735
rect 4430 7600 4800 7675
rect 4830 7735 5200 7745
rect 4830 7675 4834 7735
rect 4886 7675 5144 7735
rect 5196 7675 5200 7735
rect 4830 7600 5200 7675
rect 5230 7735 5600 7745
rect 5230 7675 5234 7735
rect 5286 7675 5544 7735
rect 5596 7675 5600 7735
rect 5230 7600 5600 7675
rect 5630 7735 6000 7745
rect 5630 7675 5634 7735
rect 5686 7675 5944 7735
rect 5996 7675 6000 7735
rect 5630 7600 6000 7675
rect 3230 7560 6000 7600
rect 3230 7475 3600 7560
rect 3230 7415 3234 7475
rect 3286 7415 3544 7475
rect 3596 7415 3600 7475
rect 3230 7405 3600 7415
rect 3630 7475 4000 7560
rect 3630 7415 3634 7475
rect 3686 7415 3944 7475
rect 3996 7415 4000 7475
rect 3630 7405 4000 7415
rect 4030 7475 4400 7560
rect 4030 7415 4034 7475
rect 4086 7415 4344 7475
rect 4396 7415 4400 7475
rect 4030 7405 4400 7415
rect 4430 7475 4800 7560
rect 4430 7415 4434 7475
rect 4486 7415 4744 7475
rect 4796 7415 4800 7475
rect 4430 7405 4800 7415
rect 4830 7475 5200 7560
rect 4830 7415 4834 7475
rect 4886 7415 5144 7475
rect 5196 7415 5200 7475
rect 4830 7405 5200 7415
rect 5230 7475 5600 7560
rect 5230 7415 5234 7475
rect 5286 7415 5544 7475
rect 5596 7415 5600 7475
rect 5230 7405 5600 7415
rect 5630 7475 6000 7560
rect 5630 7415 5634 7475
rect 5686 7415 5944 7475
rect 5996 7415 6000 7475
rect 5630 7405 6000 7415
rect 6030 7735 6400 7745
rect 6030 7675 6034 7735
rect 6086 7675 6344 7735
rect 6396 7675 6400 7735
rect 6030 7600 6400 7675
rect 6430 7735 6800 7745
rect 6430 7675 6434 7735
rect 6486 7675 6744 7735
rect 6796 7675 6800 7735
rect 6430 7600 6800 7675
rect 6830 7735 7200 7745
rect 6830 7675 6834 7735
rect 6886 7675 7144 7735
rect 7196 7675 7200 7735
rect 6830 7600 7200 7675
rect 7230 7735 7600 7745
rect 7230 7675 7234 7735
rect 7286 7675 7544 7735
rect 7596 7675 7600 7735
rect 7230 7600 7600 7675
rect 7630 7735 8000 7745
rect 7630 7675 7634 7735
rect 7686 7675 7944 7735
rect 7996 7675 8000 7735
rect 7630 7600 8000 7675
rect 8030 7735 8400 7745
rect 8030 7675 8034 7735
rect 8086 7675 8344 7735
rect 8396 7675 8400 7735
rect 8030 7600 8400 7675
rect 8430 7735 8800 7745
rect 8430 7675 8434 7735
rect 8486 7675 8744 7735
rect 8796 7675 8800 7735
rect 8430 7600 8800 7675
rect 8830 7735 9200 7745
rect 8830 7675 8834 7735
rect 8886 7675 9144 7735
rect 9196 7675 9200 7735
rect 8830 7600 9200 7675
rect 9230 7735 9600 7745
rect 9230 7675 9234 7735
rect 9286 7675 9544 7735
rect 9596 7675 9600 7735
rect 9230 7600 9600 7675
rect 9630 7735 10000 7745
rect 9630 7675 9634 7735
rect 9686 7675 9944 7735
rect 9996 7675 10000 7735
rect 9630 7600 10000 7675
rect 10030 7735 10400 7745
rect 10030 7675 10034 7735
rect 10086 7675 10344 7735
rect 10396 7675 10400 7735
rect 10030 7600 10400 7675
rect 10430 7735 10800 7745
rect 10430 7675 10434 7735
rect 10486 7675 10744 7735
rect 10796 7675 10800 7735
rect 10430 7600 10800 7675
rect 10830 7735 11200 7745
rect 10830 7675 10834 7735
rect 10886 7675 11144 7735
rect 11196 7675 11200 7735
rect 10830 7600 11200 7675
rect 11230 7735 11600 7745
rect 11230 7675 11234 7735
rect 11286 7675 11544 7735
rect 11596 7675 11600 7735
rect 11230 7600 11600 7675
rect 11630 7735 12000 7745
rect 11630 7675 11634 7735
rect 11686 7675 11944 7735
rect 11996 7675 12000 7735
rect 11630 7600 12000 7675
rect 12030 7735 12400 7745
rect 12030 7675 12034 7735
rect 12086 7675 12344 7735
rect 12396 7675 12400 7735
rect 12030 7600 12400 7675
rect 12430 7735 12800 7745
rect 12430 7675 12434 7735
rect 12486 7675 12744 7735
rect 12796 7675 12800 7735
rect 12430 7600 12800 7675
rect 12830 7735 13200 7745
rect 12830 7675 12834 7735
rect 12886 7675 13144 7735
rect 13196 7675 13200 7735
rect 12830 7600 13200 7675
rect 6030 7560 13200 7600
rect 6030 7475 6400 7560
rect 6030 7415 6034 7475
rect 6086 7415 6344 7475
rect 6396 7415 6400 7475
rect 6030 7405 6400 7415
rect 6430 7475 6800 7560
rect 6430 7415 6434 7475
rect 6486 7415 6744 7475
rect 6796 7415 6800 7475
rect 6430 7405 6800 7415
rect 6830 7475 7200 7560
rect 6830 7415 6834 7475
rect 6886 7415 7144 7475
rect 7196 7415 7200 7475
rect 6830 7405 7200 7415
rect 7230 7475 7600 7560
rect 7230 7415 7234 7475
rect 7286 7415 7544 7475
rect 7596 7415 7600 7475
rect 7230 7405 7600 7415
rect 7630 7475 8000 7560
rect 7630 7415 7634 7475
rect 7686 7415 7944 7475
rect 7996 7415 8000 7475
rect 7630 7405 8000 7415
rect 8030 7475 8400 7560
rect 8030 7415 8034 7475
rect 8086 7415 8344 7475
rect 8396 7415 8400 7475
rect 8030 7405 8400 7415
rect 8430 7475 8800 7560
rect 8430 7415 8434 7475
rect 8486 7415 8744 7475
rect 8796 7415 8800 7475
rect 8430 7405 8800 7415
rect 8830 7475 9200 7560
rect 8830 7415 8834 7475
rect 8886 7415 9144 7475
rect 9196 7415 9200 7475
rect 8830 7405 9200 7415
rect 9230 7475 9600 7560
rect 9230 7415 9234 7475
rect 9286 7415 9544 7475
rect 9596 7415 9600 7475
rect 9230 7405 9600 7415
rect 9630 7475 10000 7560
rect 9630 7415 9634 7475
rect 9686 7415 9944 7475
rect 9996 7415 10000 7475
rect 9630 7405 10000 7415
rect 10030 7475 10400 7560
rect 10030 7415 10034 7475
rect 10086 7415 10344 7475
rect 10396 7415 10400 7475
rect 10030 7405 10400 7415
rect 10430 7475 10800 7560
rect 10430 7415 10434 7475
rect 10486 7415 10744 7475
rect 10796 7415 10800 7475
rect 10430 7405 10800 7415
rect 10830 7475 11200 7560
rect 10830 7415 10834 7475
rect 10886 7415 11144 7475
rect 11196 7415 11200 7475
rect 10830 7405 11200 7415
rect 11230 7475 11600 7560
rect 11230 7415 11234 7475
rect 11286 7415 11544 7475
rect 11596 7415 11600 7475
rect 11230 7405 11600 7415
rect 11630 7475 12000 7560
rect 11630 7415 11634 7475
rect 11686 7415 11944 7475
rect 11996 7415 12000 7475
rect 11630 7405 12000 7415
rect 12030 7475 12400 7560
rect 12030 7415 12034 7475
rect 12086 7415 12344 7475
rect 12396 7415 12400 7475
rect 12030 7405 12400 7415
rect 12430 7475 12800 7560
rect 12430 7415 12434 7475
rect 12486 7415 12744 7475
rect 12796 7415 12800 7475
rect 12430 7405 12800 7415
rect 12830 7475 13200 7560
rect 12830 7415 12834 7475
rect 12886 7415 13144 7475
rect 13196 7415 13200 7475
rect 12830 7405 13200 7415
rect -330 7375 -324 7405
rect 30 7375 70 7405
rect 430 7375 470 7405
rect 830 7375 870 7405
rect 1230 7375 1270 7405
rect 1630 7375 1670 7405
rect 2030 7375 2070 7405
rect 2430 7375 2470 7405
rect 2830 7375 2870 7405
rect 3230 7375 3270 7405
rect 3630 7375 3670 7405
rect 4030 7375 4070 7405
rect 4430 7375 4470 7405
rect 4830 7375 4870 7405
rect 5230 7375 5270 7405
rect 5630 7375 5670 7405
rect 6030 7375 6070 7405
rect 6430 7375 6470 7405
rect 6830 7375 6870 7405
rect 7230 7375 7270 7405
rect 7630 7375 7670 7405
rect 8030 7375 8070 7405
rect 8430 7375 8470 7405
rect 8830 7375 8870 7405
rect 9230 7375 9270 7405
rect 9630 7375 9670 7405
rect 10030 7375 10070 7405
rect 10430 7375 10470 7405
rect 10830 7375 10870 7405
rect 11230 7375 11270 7405
rect 11630 7375 11670 7405
rect 12030 7375 12070 7405
rect 12430 7375 12470 7405
rect -330 7365 0 7375
rect -314 7305 -56 7365
rect -4 7305 0 7365
rect -330 7105 0 7305
rect -314 7045 -56 7105
rect -4 7045 0 7105
rect -330 7035 0 7045
rect 30 7365 400 7375
rect 30 7305 34 7365
rect 86 7305 344 7365
rect 396 7305 400 7365
rect 30 7230 400 7305
rect 430 7365 800 7375
rect 430 7305 434 7365
rect 486 7305 744 7365
rect 796 7305 800 7365
rect 430 7230 800 7305
rect 830 7365 1200 7375
rect 830 7305 834 7365
rect 886 7305 1144 7365
rect 1196 7305 1200 7365
rect 830 7230 1200 7305
rect 1230 7365 1600 7375
rect 1230 7305 1234 7365
rect 1286 7305 1544 7365
rect 1596 7305 1600 7365
rect 1230 7230 1600 7305
rect 1630 7365 2000 7375
rect 1630 7305 1634 7365
rect 1686 7305 1944 7365
rect 1996 7305 2000 7365
rect 1630 7230 2000 7305
rect 2030 7365 2400 7375
rect 2030 7305 2034 7365
rect 2086 7305 2344 7365
rect 2396 7305 2400 7365
rect 2030 7230 2400 7305
rect 2430 7365 2800 7375
rect 2430 7305 2434 7365
rect 2486 7305 2744 7365
rect 2796 7305 2800 7365
rect 2430 7230 2800 7305
rect 2830 7365 3200 7375
rect 2830 7305 2834 7365
rect 2886 7305 3144 7365
rect 3196 7305 3200 7365
rect 2830 7230 3200 7305
rect 30 7190 3200 7230
rect 30 7105 400 7190
rect 30 7045 34 7105
rect 86 7045 344 7105
rect 396 7045 400 7105
rect 30 7035 400 7045
rect 430 7105 800 7190
rect 430 7045 434 7105
rect 486 7045 744 7105
rect 796 7045 800 7105
rect 430 7035 800 7045
rect 830 7105 1200 7190
rect 830 7045 834 7105
rect 886 7045 1144 7105
rect 1196 7045 1200 7105
rect 830 7035 1200 7045
rect 1230 7105 1600 7190
rect 1230 7045 1234 7105
rect 1286 7045 1544 7105
rect 1596 7045 1600 7105
rect 1230 7035 1600 7045
rect 1630 7105 2000 7190
rect 1630 7045 1634 7105
rect 1686 7045 1944 7105
rect 1996 7045 2000 7105
rect 1630 7035 2000 7045
rect 2030 7105 2400 7190
rect 2030 7045 2034 7105
rect 2086 7045 2344 7105
rect 2396 7045 2400 7105
rect 2030 7035 2400 7045
rect 2430 7105 2800 7190
rect 2430 7045 2434 7105
rect 2486 7045 2744 7105
rect 2796 7045 2800 7105
rect 2430 7035 2800 7045
rect 2830 7105 3200 7190
rect 2830 7045 2834 7105
rect 2886 7045 3144 7105
rect 3196 7045 3200 7105
rect 2830 7035 3200 7045
rect 3230 7365 3600 7375
rect 3230 7305 3234 7365
rect 3286 7305 3544 7365
rect 3596 7305 3600 7365
rect 3230 7230 3600 7305
rect 3630 7365 4000 7375
rect 3630 7305 3634 7365
rect 3686 7305 3944 7365
rect 3996 7305 4000 7365
rect 3630 7230 4000 7305
rect 4030 7365 4400 7375
rect 4030 7305 4034 7365
rect 4086 7305 4344 7365
rect 4396 7305 4400 7365
rect 4030 7230 4400 7305
rect 4430 7365 4800 7375
rect 4430 7305 4434 7365
rect 4486 7305 4744 7365
rect 4796 7305 4800 7365
rect 4430 7230 4800 7305
rect 4830 7365 5200 7375
rect 4830 7305 4834 7365
rect 4886 7305 5144 7365
rect 5196 7305 5200 7365
rect 4830 7230 5200 7305
rect 5230 7365 5600 7375
rect 5230 7305 5234 7365
rect 5286 7305 5544 7365
rect 5596 7305 5600 7365
rect 5230 7230 5600 7305
rect 5630 7365 6000 7375
rect 5630 7305 5634 7365
rect 5686 7305 5944 7365
rect 5996 7305 6000 7365
rect 5630 7230 6000 7305
rect 3230 7190 6000 7230
rect 3230 7105 3600 7190
rect 3230 7045 3234 7105
rect 3286 7045 3544 7105
rect 3596 7045 3600 7105
rect 3230 7035 3600 7045
rect 3630 7105 4000 7190
rect 3630 7045 3634 7105
rect 3686 7045 3944 7105
rect 3996 7045 4000 7105
rect 3630 7035 4000 7045
rect 4030 7105 4400 7190
rect 4030 7045 4034 7105
rect 4086 7045 4344 7105
rect 4396 7045 4400 7105
rect 4030 7035 4400 7045
rect 4430 7105 4800 7190
rect 4430 7045 4434 7105
rect 4486 7045 4744 7105
rect 4796 7045 4800 7105
rect 4430 7035 4800 7045
rect 4830 7105 5200 7190
rect 4830 7045 4834 7105
rect 4886 7045 5144 7105
rect 5196 7045 5200 7105
rect 4830 7035 5200 7045
rect 5230 7105 5600 7190
rect 5230 7045 5234 7105
rect 5286 7045 5544 7105
rect 5596 7045 5600 7105
rect 5230 7035 5600 7045
rect 5630 7105 6000 7190
rect 5630 7045 5634 7105
rect 5686 7045 5944 7105
rect 5996 7045 6000 7105
rect 5630 7035 6000 7045
rect 6030 7365 6400 7375
rect 6030 7305 6034 7365
rect 6086 7305 6344 7365
rect 6396 7305 6400 7365
rect 6030 7230 6400 7305
rect 6430 7365 6800 7375
rect 6430 7305 6434 7365
rect 6486 7305 6744 7365
rect 6796 7305 6800 7365
rect 6430 7230 6800 7305
rect 6830 7365 7200 7375
rect 6830 7305 6834 7365
rect 6886 7305 7144 7365
rect 7196 7305 7200 7365
rect 6830 7230 7200 7305
rect 7230 7365 7600 7375
rect 7230 7305 7234 7365
rect 7286 7305 7544 7365
rect 7596 7305 7600 7365
rect 7230 7230 7600 7305
rect 7630 7365 8000 7375
rect 7630 7305 7634 7365
rect 7686 7305 7944 7365
rect 7996 7305 8000 7365
rect 7630 7230 8000 7305
rect 8030 7365 8400 7375
rect 8030 7305 8034 7365
rect 8086 7305 8344 7365
rect 8396 7305 8400 7365
rect 8030 7230 8400 7305
rect 8430 7365 8800 7375
rect 8430 7305 8434 7365
rect 8486 7305 8744 7365
rect 8796 7305 8800 7365
rect 8430 7230 8800 7305
rect 8830 7365 9200 7375
rect 8830 7305 8834 7365
rect 8886 7305 9144 7365
rect 9196 7305 9200 7365
rect 8830 7230 9200 7305
rect 9230 7365 9600 7375
rect 9230 7305 9234 7365
rect 9286 7305 9544 7365
rect 9596 7305 9600 7365
rect 9230 7230 9600 7305
rect 9630 7365 10000 7375
rect 9630 7305 9634 7365
rect 9686 7305 9944 7365
rect 9996 7305 10000 7365
rect 9630 7230 10000 7305
rect 10030 7365 10400 7375
rect 10030 7305 10034 7365
rect 10086 7305 10344 7365
rect 10396 7305 10400 7365
rect 10030 7230 10400 7305
rect 10430 7365 10800 7375
rect 10430 7305 10434 7365
rect 10486 7305 10744 7365
rect 10796 7305 10800 7365
rect 10430 7230 10800 7305
rect 10830 7365 11200 7375
rect 10830 7305 10834 7365
rect 10886 7305 11144 7365
rect 11196 7305 11200 7365
rect 10830 7230 11200 7305
rect 11230 7365 11600 7375
rect 11230 7305 11234 7365
rect 11286 7305 11544 7365
rect 11596 7305 11600 7365
rect 11230 7230 11600 7305
rect 11630 7365 12000 7375
rect 11630 7305 11634 7365
rect 11686 7305 11944 7365
rect 11996 7305 12000 7365
rect 11630 7230 12000 7305
rect 12030 7365 12400 7375
rect 12030 7305 12034 7365
rect 12086 7305 12344 7365
rect 12396 7305 12400 7365
rect 12030 7230 12400 7305
rect 12430 7365 12800 7375
rect 12430 7305 12434 7365
rect 12486 7305 12744 7365
rect 12796 7305 12800 7365
rect 12430 7230 12800 7305
rect 12830 7365 13200 7375
rect 12830 7305 12834 7365
rect 12886 7305 13144 7365
rect 13196 7305 13200 7365
rect 12830 7230 13200 7305
rect 6030 7190 13200 7230
rect 6030 7105 6400 7190
rect 6030 7045 6034 7105
rect 6086 7045 6344 7105
rect 6396 7045 6400 7105
rect 6030 7035 6400 7045
rect 6430 7105 6800 7190
rect 6430 7045 6434 7105
rect 6486 7045 6744 7105
rect 6796 7045 6800 7105
rect 6430 7035 6800 7045
rect 6830 7105 7200 7190
rect 6830 7045 6834 7105
rect 6886 7045 7144 7105
rect 7196 7045 7200 7105
rect 6830 7035 7200 7045
rect 7230 7105 7600 7190
rect 7230 7045 7234 7105
rect 7286 7045 7544 7105
rect 7596 7045 7600 7105
rect 7230 7035 7600 7045
rect 7630 7105 8000 7190
rect 7630 7045 7634 7105
rect 7686 7045 7944 7105
rect 7996 7045 8000 7105
rect 7630 7035 8000 7045
rect 8030 7105 8400 7190
rect 8030 7045 8034 7105
rect 8086 7045 8344 7105
rect 8396 7045 8400 7105
rect 8030 7035 8400 7045
rect 8430 7105 8800 7190
rect 8430 7045 8434 7105
rect 8486 7045 8744 7105
rect 8796 7045 8800 7105
rect 8430 7035 8800 7045
rect 8830 7105 9200 7190
rect 8830 7045 8834 7105
rect 8886 7045 9144 7105
rect 9196 7045 9200 7105
rect 8830 7035 9200 7045
rect 9230 7105 9600 7190
rect 9230 7045 9234 7105
rect 9286 7045 9544 7105
rect 9596 7045 9600 7105
rect 9230 7035 9600 7045
rect 9630 7105 10000 7190
rect 9630 7045 9634 7105
rect 9686 7045 9944 7105
rect 9996 7045 10000 7105
rect 9630 7035 10000 7045
rect 10030 7105 10400 7190
rect 10030 7045 10034 7105
rect 10086 7045 10344 7105
rect 10396 7045 10400 7105
rect 10030 7035 10400 7045
rect 10430 7105 10800 7190
rect 10430 7045 10434 7105
rect 10486 7045 10744 7105
rect 10796 7045 10800 7105
rect 10430 7035 10800 7045
rect 10830 7105 11200 7190
rect 10830 7045 10834 7105
rect 10886 7045 11144 7105
rect 11196 7045 11200 7105
rect 10830 7035 11200 7045
rect 11230 7105 11600 7190
rect 11230 7045 11234 7105
rect 11286 7045 11544 7105
rect 11596 7045 11600 7105
rect 11230 7035 11600 7045
rect 11630 7105 12000 7190
rect 11630 7045 11634 7105
rect 11686 7045 11944 7105
rect 11996 7045 12000 7105
rect 11630 7035 12000 7045
rect 12030 7105 12400 7190
rect 12030 7045 12034 7105
rect 12086 7045 12344 7105
rect 12396 7045 12400 7105
rect 12030 7035 12400 7045
rect 12430 7105 12800 7190
rect 12430 7045 12434 7105
rect 12486 7045 12744 7105
rect 12796 7045 12800 7105
rect 12430 7035 12800 7045
rect 12830 7105 13200 7190
rect 12830 7045 12834 7105
rect 12886 7045 13144 7105
rect 13196 7045 13200 7105
rect 12830 7035 13200 7045
rect -330 7005 -324 7035
rect 30 7005 70 7035
rect 430 7005 470 7035
rect 830 7005 870 7035
rect 1230 7005 1270 7035
rect 1630 7005 1670 7035
rect 2030 7005 2070 7035
rect 2430 7005 2470 7035
rect 2830 7005 2870 7035
rect 3230 7005 3270 7035
rect 3630 7005 3670 7035
rect 4030 7005 4070 7035
rect 4430 7005 4470 7035
rect 4830 7005 4870 7035
rect 5230 7005 5270 7035
rect 5630 7005 5670 7035
rect 6030 7005 6070 7035
rect 6430 7005 6470 7035
rect 6830 7005 6870 7035
rect 7230 7005 7270 7035
rect 7630 7005 7670 7035
rect 8030 7005 8070 7035
rect 8430 7005 8470 7035
rect 8830 7005 8870 7035
rect 9230 7005 9270 7035
rect 9630 7005 9670 7035
rect 10030 7005 10070 7035
rect 10430 7005 10470 7035
rect 10830 7005 10870 7035
rect 11230 7005 11270 7035
rect 11630 7005 11670 7035
rect 12030 7005 12070 7035
rect 12430 7005 12470 7035
rect -330 6995 0 7005
rect -314 6935 -56 6995
rect -4 6935 0 6995
rect -330 6735 0 6935
rect -314 6675 -56 6735
rect -4 6675 0 6735
rect -330 6665 0 6675
rect 30 6995 400 7005
rect 30 6935 34 6995
rect 86 6935 344 6995
rect 396 6935 400 6995
rect 30 6860 400 6935
rect 430 6995 800 7005
rect 430 6935 434 6995
rect 486 6935 744 6995
rect 796 6935 800 6995
rect 430 6860 800 6935
rect 830 6995 1200 7005
rect 830 6935 834 6995
rect 886 6935 1144 6995
rect 1196 6935 1200 6995
rect 830 6860 1200 6935
rect 1230 6995 1600 7005
rect 1230 6935 1234 6995
rect 1286 6935 1544 6995
rect 1596 6935 1600 6995
rect 1230 6860 1600 6935
rect 1630 6995 2000 7005
rect 1630 6935 1634 6995
rect 1686 6935 1944 6995
rect 1996 6935 2000 6995
rect 1630 6860 2000 6935
rect 2030 6995 2400 7005
rect 2030 6935 2034 6995
rect 2086 6935 2344 6995
rect 2396 6935 2400 6995
rect 2030 6860 2400 6935
rect 2430 6995 2800 7005
rect 2430 6935 2434 6995
rect 2486 6935 2744 6995
rect 2796 6935 2800 6995
rect 2430 6860 2800 6935
rect 2830 6995 3200 7005
rect 2830 6935 2834 6995
rect 2886 6935 3144 6995
rect 3196 6935 3200 6995
rect 2830 6860 3200 6935
rect 30 6820 3200 6860
rect 30 6735 400 6820
rect 30 6675 34 6735
rect 86 6675 344 6735
rect 396 6675 400 6735
rect 30 6665 400 6675
rect 430 6735 800 6820
rect 430 6675 434 6735
rect 486 6675 744 6735
rect 796 6675 800 6735
rect 430 6665 800 6675
rect 830 6735 1200 6820
rect 830 6675 834 6735
rect 886 6675 1144 6735
rect 1196 6675 1200 6735
rect 830 6665 1200 6675
rect 1230 6735 1600 6820
rect 1230 6675 1234 6735
rect 1286 6675 1544 6735
rect 1596 6675 1600 6735
rect 1230 6665 1600 6675
rect 1630 6735 2000 6820
rect 1630 6675 1634 6735
rect 1686 6675 1944 6735
rect 1996 6675 2000 6735
rect 1630 6665 2000 6675
rect 2030 6735 2400 6820
rect 2030 6675 2034 6735
rect 2086 6675 2344 6735
rect 2396 6675 2400 6735
rect 2030 6665 2400 6675
rect 2430 6735 2800 6820
rect 2430 6675 2434 6735
rect 2486 6675 2744 6735
rect 2796 6675 2800 6735
rect 2430 6665 2800 6675
rect 2830 6735 3200 6820
rect 2830 6675 2834 6735
rect 2886 6675 3144 6735
rect 3196 6675 3200 6735
rect 2830 6665 3200 6675
rect 3230 6995 3600 7005
rect 3230 6935 3234 6995
rect 3286 6935 3544 6995
rect 3596 6935 3600 6995
rect 3230 6860 3600 6935
rect 3630 6995 4000 7005
rect 3630 6935 3634 6995
rect 3686 6935 3944 6995
rect 3996 6935 4000 6995
rect 3630 6860 4000 6935
rect 4030 6995 4400 7005
rect 4030 6935 4034 6995
rect 4086 6935 4344 6995
rect 4396 6935 4400 6995
rect 4030 6860 4400 6935
rect 4430 6995 4800 7005
rect 4430 6935 4434 6995
rect 4486 6935 4744 6995
rect 4796 6935 4800 6995
rect 4430 6860 4800 6935
rect 4830 6995 5200 7005
rect 4830 6935 4834 6995
rect 4886 6935 5144 6995
rect 5196 6935 5200 6995
rect 4830 6860 5200 6935
rect 5230 6995 5600 7005
rect 5230 6935 5234 6995
rect 5286 6935 5544 6995
rect 5596 6935 5600 6995
rect 5230 6860 5600 6935
rect 5630 6995 6000 7005
rect 5630 6935 5634 6995
rect 5686 6935 5944 6995
rect 5996 6935 6000 6995
rect 5630 6860 6000 6935
rect 3230 6820 6000 6860
rect 3230 6735 3600 6820
rect 3230 6675 3234 6735
rect 3286 6675 3544 6735
rect 3596 6675 3600 6735
rect 3230 6665 3600 6675
rect 3630 6735 4000 6820
rect 3630 6675 3634 6735
rect 3686 6675 3944 6735
rect 3996 6675 4000 6735
rect 3630 6665 4000 6675
rect 4030 6735 4400 6820
rect 4030 6675 4034 6735
rect 4086 6675 4344 6735
rect 4396 6675 4400 6735
rect 4030 6665 4400 6675
rect 4430 6735 4800 6820
rect 4430 6675 4434 6735
rect 4486 6675 4744 6735
rect 4796 6675 4800 6735
rect 4430 6665 4800 6675
rect 4830 6735 5200 6820
rect 4830 6675 4834 6735
rect 4886 6675 5144 6735
rect 5196 6675 5200 6735
rect 4830 6665 5200 6675
rect 5230 6735 5600 6820
rect 5230 6675 5234 6735
rect 5286 6675 5544 6735
rect 5596 6675 5600 6735
rect 5230 6665 5600 6675
rect 5630 6735 6000 6820
rect 5630 6675 5634 6735
rect 5686 6675 5944 6735
rect 5996 6675 6000 6735
rect 5630 6665 6000 6675
rect 6030 6995 6400 7005
rect 6030 6935 6034 6995
rect 6086 6935 6344 6995
rect 6396 6935 6400 6995
rect 6030 6860 6400 6935
rect 6430 6995 6800 7005
rect 6430 6935 6434 6995
rect 6486 6935 6744 6995
rect 6796 6935 6800 6995
rect 6430 6860 6800 6935
rect 6830 6995 7200 7005
rect 6830 6935 6834 6995
rect 6886 6935 7144 6995
rect 7196 6935 7200 6995
rect 6830 6860 7200 6935
rect 7230 6995 7600 7005
rect 7230 6935 7234 6995
rect 7286 6935 7544 6995
rect 7596 6935 7600 6995
rect 7230 6860 7600 6935
rect 7630 6995 8000 7005
rect 7630 6935 7634 6995
rect 7686 6935 7944 6995
rect 7996 6935 8000 6995
rect 7630 6860 8000 6935
rect 8030 6995 8400 7005
rect 8030 6935 8034 6995
rect 8086 6935 8344 6995
rect 8396 6935 8400 6995
rect 8030 6860 8400 6935
rect 8430 6995 8800 7005
rect 8430 6935 8434 6995
rect 8486 6935 8744 6995
rect 8796 6935 8800 6995
rect 8430 6860 8800 6935
rect 8830 6995 9200 7005
rect 8830 6935 8834 6995
rect 8886 6935 9144 6995
rect 9196 6935 9200 6995
rect 8830 6860 9200 6935
rect 9230 6995 9600 7005
rect 9230 6935 9234 6995
rect 9286 6935 9544 6995
rect 9596 6935 9600 6995
rect 9230 6860 9600 6935
rect 9630 6995 10000 7005
rect 9630 6935 9634 6995
rect 9686 6935 9944 6995
rect 9996 6935 10000 6995
rect 9630 6860 10000 6935
rect 10030 6995 10400 7005
rect 10030 6935 10034 6995
rect 10086 6935 10344 6995
rect 10396 6935 10400 6995
rect 10030 6860 10400 6935
rect 10430 6995 10800 7005
rect 10430 6935 10434 6995
rect 10486 6935 10744 6995
rect 10796 6935 10800 6995
rect 10430 6860 10800 6935
rect 10830 6995 11200 7005
rect 10830 6935 10834 6995
rect 10886 6935 11144 6995
rect 11196 6935 11200 6995
rect 10830 6860 11200 6935
rect 11230 6995 11600 7005
rect 11230 6935 11234 6995
rect 11286 6935 11544 6995
rect 11596 6935 11600 6995
rect 11230 6860 11600 6935
rect 11630 6995 12000 7005
rect 11630 6935 11634 6995
rect 11686 6935 11944 6995
rect 11996 6935 12000 6995
rect 11630 6860 12000 6935
rect 12030 6995 12400 7005
rect 12030 6935 12034 6995
rect 12086 6935 12344 6995
rect 12396 6935 12400 6995
rect 12030 6860 12400 6935
rect 12430 6995 12800 7005
rect 12430 6935 12434 6995
rect 12486 6935 12744 6995
rect 12796 6935 12800 6995
rect 12430 6860 12800 6935
rect 12830 6995 13200 7005
rect 12830 6935 12834 6995
rect 12886 6935 13144 6995
rect 13196 6935 13200 6995
rect 12830 6860 13200 6935
rect 6030 6820 13200 6860
rect 6030 6735 6400 6820
rect 6030 6675 6034 6735
rect 6086 6675 6344 6735
rect 6396 6675 6400 6735
rect 6030 6665 6400 6675
rect 6430 6735 6800 6820
rect 6430 6675 6434 6735
rect 6486 6675 6744 6735
rect 6796 6675 6800 6735
rect 6430 6665 6800 6675
rect 6830 6735 7200 6820
rect 6830 6675 6834 6735
rect 6886 6675 7144 6735
rect 7196 6675 7200 6735
rect 6830 6665 7200 6675
rect 7230 6735 7600 6820
rect 7230 6675 7234 6735
rect 7286 6675 7544 6735
rect 7596 6675 7600 6735
rect 7230 6665 7600 6675
rect 7630 6735 8000 6820
rect 7630 6675 7634 6735
rect 7686 6675 7944 6735
rect 7996 6675 8000 6735
rect 7630 6665 8000 6675
rect 8030 6735 8400 6820
rect 8030 6675 8034 6735
rect 8086 6675 8344 6735
rect 8396 6675 8400 6735
rect 8030 6665 8400 6675
rect 8430 6735 8800 6820
rect 8430 6675 8434 6735
rect 8486 6675 8744 6735
rect 8796 6675 8800 6735
rect 8430 6665 8800 6675
rect 8830 6735 9200 6820
rect 8830 6675 8834 6735
rect 8886 6675 9144 6735
rect 9196 6675 9200 6735
rect 8830 6665 9200 6675
rect 9230 6735 9600 6820
rect 9230 6675 9234 6735
rect 9286 6675 9544 6735
rect 9596 6675 9600 6735
rect 9230 6665 9600 6675
rect 9630 6735 10000 6820
rect 9630 6675 9634 6735
rect 9686 6675 9944 6735
rect 9996 6675 10000 6735
rect 9630 6665 10000 6675
rect 10030 6735 10400 6820
rect 10030 6675 10034 6735
rect 10086 6675 10344 6735
rect 10396 6675 10400 6735
rect 10030 6665 10400 6675
rect 10430 6735 10800 6820
rect 10430 6675 10434 6735
rect 10486 6675 10744 6735
rect 10796 6675 10800 6735
rect 10430 6665 10800 6675
rect 10830 6735 11200 6820
rect 10830 6675 10834 6735
rect 10886 6675 11144 6735
rect 11196 6675 11200 6735
rect 10830 6665 11200 6675
rect 11230 6735 11600 6820
rect 11230 6675 11234 6735
rect 11286 6675 11544 6735
rect 11596 6675 11600 6735
rect 11230 6665 11600 6675
rect 11630 6735 12000 6820
rect 11630 6675 11634 6735
rect 11686 6675 11944 6735
rect 11996 6675 12000 6735
rect 11630 6665 12000 6675
rect 12030 6735 12400 6820
rect 12030 6675 12034 6735
rect 12086 6675 12344 6735
rect 12396 6675 12400 6735
rect 12030 6665 12400 6675
rect 12430 6735 12800 6820
rect 12430 6675 12434 6735
rect 12486 6675 12744 6735
rect 12796 6675 12800 6735
rect 12430 6665 12800 6675
rect 12830 6735 13200 6820
rect 12830 6675 12834 6735
rect 12886 6675 13144 6735
rect 13196 6675 13200 6735
rect 12830 6665 13200 6675
rect -330 6635 -324 6665
rect 30 6635 70 6665
rect 430 6635 470 6665
rect 830 6635 870 6665
rect 1230 6635 1270 6665
rect 1630 6635 1670 6665
rect 2030 6635 2070 6665
rect 2430 6635 2470 6665
rect 2830 6635 2870 6665
rect 3230 6635 3270 6665
rect 3630 6635 3670 6665
rect 4030 6635 4070 6665
rect 4430 6635 4470 6665
rect 4830 6635 4870 6665
rect 5230 6635 5270 6665
rect 5630 6635 5670 6665
rect 6030 6635 6070 6665
rect 6430 6635 6470 6665
rect 6830 6635 6870 6665
rect 7230 6635 7270 6665
rect 7630 6635 7670 6665
rect 8030 6635 8070 6665
rect 8430 6635 8470 6665
rect 8830 6635 8870 6665
rect 9230 6635 9270 6665
rect 9630 6635 9670 6665
rect 10030 6635 10070 6665
rect 10430 6635 10470 6665
rect 10830 6635 10870 6665
rect 11230 6635 11270 6665
rect 11630 6635 11670 6665
rect 12030 6635 12070 6665
rect 12430 6635 12470 6665
rect -330 6625 0 6635
rect -314 6565 -56 6625
rect -4 6565 0 6625
rect -330 6365 0 6565
rect -314 6305 -56 6365
rect -4 6305 0 6365
rect -330 6295 0 6305
rect 30 6625 400 6635
rect 30 6565 34 6625
rect 86 6565 344 6625
rect 396 6565 400 6625
rect 30 6490 400 6565
rect 430 6625 800 6635
rect 430 6565 434 6625
rect 486 6565 744 6625
rect 796 6565 800 6625
rect 430 6490 800 6565
rect 830 6625 1200 6635
rect 830 6565 834 6625
rect 886 6565 1144 6625
rect 1196 6565 1200 6625
rect 830 6490 1200 6565
rect 1230 6625 1600 6635
rect 1230 6565 1234 6625
rect 1286 6565 1544 6625
rect 1596 6565 1600 6625
rect 1230 6490 1600 6565
rect 1630 6625 2000 6635
rect 1630 6565 1634 6625
rect 1686 6565 1944 6625
rect 1996 6565 2000 6625
rect 1630 6490 2000 6565
rect 2030 6625 2400 6635
rect 2030 6565 2034 6625
rect 2086 6565 2344 6625
rect 2396 6565 2400 6625
rect 2030 6490 2400 6565
rect 2430 6625 2800 6635
rect 2430 6565 2434 6625
rect 2486 6565 2744 6625
rect 2796 6565 2800 6625
rect 2430 6490 2800 6565
rect 2830 6625 3200 6635
rect 2830 6565 2834 6625
rect 2886 6565 3144 6625
rect 3196 6565 3200 6625
rect 2830 6490 3200 6565
rect 30 6450 3200 6490
rect 30 6365 400 6450
rect 30 6305 34 6365
rect 86 6305 344 6365
rect 396 6305 400 6365
rect 30 6295 400 6305
rect 430 6365 800 6450
rect 430 6305 434 6365
rect 486 6305 744 6365
rect 796 6305 800 6365
rect 430 6295 800 6305
rect 830 6365 1200 6450
rect 830 6305 834 6365
rect 886 6305 1144 6365
rect 1196 6305 1200 6365
rect 830 6295 1200 6305
rect 1230 6365 1600 6450
rect 1230 6305 1234 6365
rect 1286 6305 1544 6365
rect 1596 6305 1600 6365
rect 1230 6295 1600 6305
rect 1630 6365 2000 6450
rect 1630 6305 1634 6365
rect 1686 6305 1944 6365
rect 1996 6305 2000 6365
rect 1630 6295 2000 6305
rect 2030 6365 2400 6450
rect 2030 6305 2034 6365
rect 2086 6305 2344 6365
rect 2396 6305 2400 6365
rect 2030 6295 2400 6305
rect 2430 6365 2800 6450
rect 2430 6305 2434 6365
rect 2486 6305 2744 6365
rect 2796 6305 2800 6365
rect 2430 6295 2800 6305
rect 2830 6365 3200 6450
rect 2830 6305 2834 6365
rect 2886 6305 3144 6365
rect 3196 6305 3200 6365
rect 2830 6295 3200 6305
rect 3230 6625 3600 6635
rect 3230 6565 3234 6625
rect 3286 6565 3544 6625
rect 3596 6565 3600 6625
rect 3230 6490 3600 6565
rect 3630 6625 4000 6635
rect 3630 6565 3634 6625
rect 3686 6565 3944 6625
rect 3996 6565 4000 6625
rect 3630 6490 4000 6565
rect 4030 6625 4400 6635
rect 4030 6565 4034 6625
rect 4086 6565 4344 6625
rect 4396 6565 4400 6625
rect 4030 6490 4400 6565
rect 4430 6625 4800 6635
rect 4430 6565 4434 6625
rect 4486 6565 4744 6625
rect 4796 6565 4800 6625
rect 4430 6490 4800 6565
rect 4830 6625 5200 6635
rect 4830 6565 4834 6625
rect 4886 6565 5144 6625
rect 5196 6565 5200 6625
rect 4830 6490 5200 6565
rect 5230 6625 5600 6635
rect 5230 6565 5234 6625
rect 5286 6565 5544 6625
rect 5596 6565 5600 6625
rect 5230 6490 5600 6565
rect 5630 6625 6000 6635
rect 5630 6565 5634 6625
rect 5686 6565 5944 6625
rect 5996 6565 6000 6625
rect 5630 6490 6000 6565
rect 3230 6450 6000 6490
rect 3230 6365 3600 6450
rect 3230 6305 3234 6365
rect 3286 6305 3544 6365
rect 3596 6305 3600 6365
rect 3230 6295 3600 6305
rect 3630 6365 4000 6450
rect 3630 6305 3634 6365
rect 3686 6305 3944 6365
rect 3996 6305 4000 6365
rect 3630 6295 4000 6305
rect 4030 6365 4400 6450
rect 4030 6305 4034 6365
rect 4086 6305 4344 6365
rect 4396 6305 4400 6365
rect 4030 6295 4400 6305
rect 4430 6365 4800 6450
rect 4430 6305 4434 6365
rect 4486 6305 4744 6365
rect 4796 6305 4800 6365
rect 4430 6295 4800 6305
rect 4830 6365 5200 6450
rect 4830 6305 4834 6365
rect 4886 6305 5144 6365
rect 5196 6305 5200 6365
rect 4830 6295 5200 6305
rect 5230 6365 5600 6450
rect 5230 6305 5234 6365
rect 5286 6305 5544 6365
rect 5596 6305 5600 6365
rect 5230 6295 5600 6305
rect 5630 6365 6000 6450
rect 5630 6305 5634 6365
rect 5686 6305 5944 6365
rect 5996 6305 6000 6365
rect 5630 6295 6000 6305
rect 6030 6625 6400 6635
rect 6030 6565 6034 6625
rect 6086 6565 6344 6625
rect 6396 6565 6400 6625
rect 6030 6490 6400 6565
rect 6430 6625 6800 6635
rect 6430 6565 6434 6625
rect 6486 6565 6744 6625
rect 6796 6565 6800 6625
rect 6430 6490 6800 6565
rect 6830 6625 7200 6635
rect 6830 6565 6834 6625
rect 6886 6565 7144 6625
rect 7196 6565 7200 6625
rect 6830 6490 7200 6565
rect 7230 6625 7600 6635
rect 7230 6565 7234 6625
rect 7286 6565 7544 6625
rect 7596 6565 7600 6625
rect 7230 6490 7600 6565
rect 7630 6625 8000 6635
rect 7630 6565 7634 6625
rect 7686 6565 7944 6625
rect 7996 6565 8000 6625
rect 7630 6490 8000 6565
rect 8030 6625 8400 6635
rect 8030 6565 8034 6625
rect 8086 6565 8344 6625
rect 8396 6565 8400 6625
rect 8030 6490 8400 6565
rect 8430 6625 8800 6635
rect 8430 6565 8434 6625
rect 8486 6565 8744 6625
rect 8796 6565 8800 6625
rect 8430 6490 8800 6565
rect 8830 6625 9200 6635
rect 8830 6565 8834 6625
rect 8886 6565 9144 6625
rect 9196 6565 9200 6625
rect 8830 6490 9200 6565
rect 9230 6625 9600 6635
rect 9230 6565 9234 6625
rect 9286 6565 9544 6625
rect 9596 6565 9600 6625
rect 9230 6490 9600 6565
rect 9630 6625 10000 6635
rect 9630 6565 9634 6625
rect 9686 6565 9944 6625
rect 9996 6565 10000 6625
rect 9630 6490 10000 6565
rect 10030 6625 10400 6635
rect 10030 6565 10034 6625
rect 10086 6565 10344 6625
rect 10396 6565 10400 6625
rect 10030 6490 10400 6565
rect 10430 6625 10800 6635
rect 10430 6565 10434 6625
rect 10486 6565 10744 6625
rect 10796 6565 10800 6625
rect 10430 6490 10800 6565
rect 10830 6625 11200 6635
rect 10830 6565 10834 6625
rect 10886 6565 11144 6625
rect 11196 6565 11200 6625
rect 10830 6490 11200 6565
rect 11230 6625 11600 6635
rect 11230 6565 11234 6625
rect 11286 6565 11544 6625
rect 11596 6565 11600 6625
rect 11230 6490 11600 6565
rect 11630 6625 12000 6635
rect 11630 6565 11634 6625
rect 11686 6565 11944 6625
rect 11996 6565 12000 6625
rect 11630 6490 12000 6565
rect 12030 6625 12400 6635
rect 12030 6565 12034 6625
rect 12086 6565 12344 6625
rect 12396 6565 12400 6625
rect 12030 6490 12400 6565
rect 12430 6625 12800 6635
rect 12430 6565 12434 6625
rect 12486 6565 12744 6625
rect 12796 6565 12800 6625
rect 12430 6490 12800 6565
rect 12830 6625 13200 6635
rect 12830 6565 12834 6625
rect 12886 6565 13144 6625
rect 13196 6565 13200 6625
rect 12830 6490 13200 6565
rect 6030 6450 13200 6490
rect 6030 6365 6400 6450
rect 6030 6305 6034 6365
rect 6086 6305 6344 6365
rect 6396 6305 6400 6365
rect 6030 6295 6400 6305
rect 6430 6365 6800 6450
rect 6430 6305 6434 6365
rect 6486 6305 6744 6365
rect 6796 6305 6800 6365
rect 6430 6295 6800 6305
rect 6830 6365 7200 6450
rect 6830 6305 6834 6365
rect 6886 6305 7144 6365
rect 7196 6305 7200 6365
rect 6830 6295 7200 6305
rect 7230 6365 7600 6450
rect 7230 6305 7234 6365
rect 7286 6305 7544 6365
rect 7596 6305 7600 6365
rect 7230 6295 7600 6305
rect 7630 6365 8000 6450
rect 7630 6305 7634 6365
rect 7686 6305 7944 6365
rect 7996 6305 8000 6365
rect 7630 6295 8000 6305
rect 8030 6365 8400 6450
rect 8030 6305 8034 6365
rect 8086 6305 8344 6365
rect 8396 6305 8400 6365
rect 8030 6295 8400 6305
rect 8430 6365 8800 6450
rect 8430 6305 8434 6365
rect 8486 6305 8744 6365
rect 8796 6305 8800 6365
rect 8430 6295 8800 6305
rect 8830 6365 9200 6450
rect 8830 6305 8834 6365
rect 8886 6305 9144 6365
rect 9196 6305 9200 6365
rect 8830 6295 9200 6305
rect 9230 6365 9600 6450
rect 9230 6305 9234 6365
rect 9286 6305 9544 6365
rect 9596 6305 9600 6365
rect 9230 6295 9600 6305
rect 9630 6365 10000 6450
rect 9630 6305 9634 6365
rect 9686 6305 9944 6365
rect 9996 6305 10000 6365
rect 9630 6295 10000 6305
rect 10030 6365 10400 6450
rect 10030 6305 10034 6365
rect 10086 6305 10344 6365
rect 10396 6305 10400 6365
rect 10030 6295 10400 6305
rect 10430 6365 10800 6450
rect 10430 6305 10434 6365
rect 10486 6305 10744 6365
rect 10796 6305 10800 6365
rect 10430 6295 10800 6305
rect 10830 6365 11200 6450
rect 10830 6305 10834 6365
rect 10886 6305 11144 6365
rect 11196 6305 11200 6365
rect 10830 6295 11200 6305
rect 11230 6365 11600 6450
rect 11230 6305 11234 6365
rect 11286 6305 11544 6365
rect 11596 6305 11600 6365
rect 11230 6295 11600 6305
rect 11630 6365 12000 6450
rect 11630 6305 11634 6365
rect 11686 6305 11944 6365
rect 11996 6305 12000 6365
rect 11630 6295 12000 6305
rect 12030 6365 12400 6450
rect 12030 6305 12034 6365
rect 12086 6305 12344 6365
rect 12396 6305 12400 6365
rect 12030 6295 12400 6305
rect 12430 6365 12800 6450
rect 12430 6305 12434 6365
rect 12486 6305 12744 6365
rect 12796 6305 12800 6365
rect 12430 6295 12800 6305
rect 12830 6365 13200 6450
rect 12830 6305 12834 6365
rect 12886 6305 13144 6365
rect 13196 6305 13200 6365
rect 12830 6295 13200 6305
rect -330 6265 -324 6295
rect 30 6265 70 6295
rect 430 6265 470 6295
rect 830 6265 870 6295
rect 1230 6265 1270 6295
rect 1630 6265 1670 6295
rect 2030 6265 2070 6295
rect 2430 6265 2470 6295
rect 2830 6265 2870 6295
rect 3230 6265 3270 6295
rect 3630 6265 3670 6295
rect 4030 6265 4070 6295
rect 4430 6265 4470 6295
rect 4830 6265 4870 6295
rect 5230 6265 5270 6295
rect 5630 6265 5670 6295
rect -330 6255 0 6265
rect -314 6195 -56 6255
rect -4 6195 0 6255
rect -330 5995 0 6195
rect -314 5935 -56 5995
rect -4 5935 0 5995
rect -330 5925 0 5935
rect 30 6255 400 6265
rect 30 6195 34 6255
rect 86 6195 344 6255
rect 396 6195 400 6255
rect 30 6120 400 6195
rect 430 6255 800 6265
rect 430 6195 434 6255
rect 486 6195 744 6255
rect 796 6195 800 6255
rect 430 6120 800 6195
rect 830 6255 1200 6265
rect 830 6195 834 6255
rect 886 6195 1144 6255
rect 1196 6195 1200 6255
rect 830 6120 1200 6195
rect 1230 6255 1600 6265
rect 1230 6195 1234 6255
rect 1286 6195 1544 6255
rect 1596 6195 1600 6255
rect 1230 6120 1600 6195
rect 1630 6255 2000 6265
rect 1630 6195 1634 6255
rect 1686 6195 1944 6255
rect 1996 6195 2000 6255
rect 1630 6120 2000 6195
rect 2030 6255 2400 6265
rect 2030 6195 2034 6255
rect 2086 6195 2344 6255
rect 2396 6195 2400 6255
rect 2030 6120 2400 6195
rect 2430 6255 2800 6265
rect 2430 6195 2434 6255
rect 2486 6195 2744 6255
rect 2796 6195 2800 6255
rect 2430 6120 2800 6195
rect 2830 6255 3200 6265
rect 2830 6195 2834 6255
rect 2886 6195 3144 6255
rect 3196 6195 3200 6255
rect 2830 6120 3200 6195
rect 30 6080 3200 6120
rect 30 5995 400 6080
rect 30 5935 34 5995
rect 86 5935 344 5995
rect 396 5935 400 5995
rect 30 5925 400 5935
rect 430 5995 800 6080
rect 430 5935 434 5995
rect 486 5935 744 5995
rect 796 5935 800 5995
rect 430 5925 800 5935
rect 830 5995 1200 6080
rect 830 5935 834 5995
rect 886 5935 1144 5995
rect 1196 5935 1200 5995
rect 830 5925 1200 5935
rect 1230 5995 1600 6080
rect 1230 5935 1234 5995
rect 1286 5935 1544 5995
rect 1596 5935 1600 5995
rect 1230 5925 1600 5935
rect 1630 5995 2000 6080
rect 1630 5935 1634 5995
rect 1686 5935 1944 5995
rect 1996 5935 2000 5995
rect 1630 5925 2000 5935
rect 2030 5995 2400 6080
rect 2030 5935 2034 5995
rect 2086 5935 2344 5995
rect 2396 5935 2400 5995
rect 2030 5925 2400 5935
rect 2430 5995 2800 6080
rect 2430 5935 2434 5995
rect 2486 5935 2744 5995
rect 2796 5935 2800 5995
rect 2430 5925 2800 5935
rect 2830 5995 3200 6080
rect 2830 5935 2834 5995
rect 2886 5935 3144 5995
rect 3196 5935 3200 5995
rect 2830 5925 3200 5935
rect 3230 6255 3600 6265
rect 3230 6195 3234 6255
rect 3286 6195 3544 6255
rect 3596 6195 3600 6255
rect 3230 6120 3600 6195
rect 3630 6255 4000 6265
rect 3630 6195 3634 6255
rect 3686 6195 3944 6255
rect 3996 6195 4000 6255
rect 3630 6120 4000 6195
rect 4030 6255 4400 6265
rect 4030 6195 4034 6255
rect 4086 6195 4344 6255
rect 4396 6195 4400 6255
rect 4030 6120 4400 6195
rect 4430 6255 4800 6265
rect 4430 6195 4434 6255
rect 4486 6195 4744 6255
rect 4796 6195 4800 6255
rect 4430 6120 4800 6195
rect 4830 6255 5200 6265
rect 4830 6195 4834 6255
rect 4886 6195 5144 6255
rect 5196 6195 5200 6255
rect 4830 6120 5200 6195
rect 5230 6255 5600 6265
rect 5230 6195 5234 6255
rect 5286 6195 5544 6255
rect 5596 6195 5600 6255
rect 5230 6120 5600 6195
rect 5630 6255 6000 6265
rect 5630 6195 5634 6255
rect 5686 6195 5944 6255
rect 5996 6195 6000 6255
rect 5630 6120 6000 6195
rect 6030 6255 6400 6265
rect 6030 6195 6034 6255
rect 6086 6195 6344 6255
rect 6396 6195 6400 6255
rect 6030 6120 6400 6195
rect 6430 6255 6800 6265
rect 6430 6195 6434 6255
rect 6486 6195 6744 6255
rect 6796 6195 6800 6255
rect 6430 6120 6800 6195
rect 6830 6255 7200 6265
rect 6830 6195 6834 6255
rect 6886 6195 7144 6255
rect 7196 6195 7200 6255
rect 6830 6120 7200 6195
rect 7230 6255 7600 6265
rect 7230 6195 7234 6255
rect 7286 6195 7544 6255
rect 7596 6195 7600 6255
rect 7230 6120 7600 6195
rect 7630 6255 8000 6265
rect 7630 6195 7634 6255
rect 7686 6195 7944 6255
rect 7996 6195 8000 6255
rect 7630 6120 8000 6195
rect 8030 6255 8400 6265
rect 8030 6195 8034 6255
rect 8086 6195 8344 6255
rect 8396 6195 8400 6255
rect 8030 6120 8400 6195
rect 8430 6255 8800 6265
rect 8430 6195 8434 6255
rect 8486 6195 8744 6255
rect 8796 6195 8800 6255
rect 8430 6120 8800 6195
rect 8830 6255 9200 6265
rect 8830 6195 8834 6255
rect 8886 6195 9144 6255
rect 9196 6195 9200 6255
rect 8830 6120 9200 6195
rect 9230 6255 9600 6265
rect 9230 6195 9234 6255
rect 9286 6195 9544 6255
rect 9596 6195 9600 6255
rect 9230 6120 9600 6195
rect 9630 6255 10000 6265
rect 9630 6195 9634 6255
rect 9686 6195 9944 6255
rect 9996 6195 10000 6255
rect 9630 6120 10000 6195
rect 10030 6255 10400 6265
rect 10030 6195 10034 6255
rect 10086 6195 10344 6255
rect 10396 6195 10400 6255
rect 10030 6120 10400 6195
rect 10430 6255 10800 6265
rect 10430 6195 10434 6255
rect 10486 6195 10744 6255
rect 10796 6195 10800 6255
rect 10430 6120 10800 6195
rect 10830 6255 11200 6265
rect 10830 6195 10834 6255
rect 10886 6195 11144 6255
rect 11196 6195 11200 6255
rect 10830 6120 11200 6195
rect 11230 6255 11600 6265
rect 11230 6195 11234 6255
rect 11286 6195 11544 6255
rect 11596 6195 11600 6255
rect 11230 6120 11600 6195
rect 11630 6255 12000 6265
rect 11630 6195 11634 6255
rect 11686 6195 11944 6255
rect 11996 6195 12000 6255
rect 11630 6120 12000 6195
rect 12030 6255 12400 6265
rect 12030 6195 12034 6255
rect 12086 6195 12344 6255
rect 12396 6195 12400 6255
rect 12030 6120 12400 6195
rect 12430 6255 12800 6265
rect 12430 6195 12434 6255
rect 12486 6195 12744 6255
rect 12796 6195 12800 6255
rect 12430 6120 12800 6195
rect 12830 6255 13200 6265
rect 12830 6195 12834 6255
rect 12886 6195 13144 6255
rect 13196 6195 13200 6255
rect 12830 6120 13200 6195
rect 3230 6080 13390 6120
rect 3230 5995 3600 6080
rect 3230 5935 3234 5995
rect 3286 5935 3544 5995
rect 3596 5935 3600 5995
rect 3230 5925 3600 5935
rect 3630 5995 4000 6080
rect 3630 5935 3634 5995
rect 3686 5935 3944 5995
rect 3996 5935 4000 5995
rect 3630 5925 4000 5935
rect 4030 5995 4400 6080
rect 4030 5935 4034 5995
rect 4086 5935 4344 5995
rect 4396 5935 4400 5995
rect 4030 5925 4400 5935
rect 4430 5995 4800 6080
rect 4430 5935 4434 5995
rect 4486 5935 4744 5995
rect 4796 5935 4800 5995
rect 4430 5925 4800 5935
rect 4830 5995 5200 6080
rect 4830 5935 4834 5995
rect 4886 5935 5144 5995
rect 5196 5935 5200 5995
rect 4830 5925 5200 5935
rect 5230 5995 5600 6080
rect 5230 5935 5234 5995
rect 5286 5935 5544 5995
rect 5596 5935 5600 5995
rect 5230 5925 5600 5935
rect 5630 5995 6000 6080
rect 5630 5935 5634 5995
rect 5686 5935 5944 5995
rect 5996 5935 6000 5995
rect 5630 5925 6000 5935
rect 6030 5995 6400 6080
rect 6030 5935 6034 5995
rect 6086 5935 6344 5995
rect 6396 5935 6400 5995
rect 6030 5925 6400 5935
rect 6430 5995 6800 6080
rect 6430 5935 6434 5995
rect 6486 5935 6744 5995
rect 6796 5935 6800 5995
rect 6430 5925 6800 5935
rect 6830 5995 7200 6080
rect 6830 5935 6834 5995
rect 6886 5935 7144 5995
rect 7196 5935 7200 5995
rect 6830 5925 7200 5935
rect 7230 5995 7600 6080
rect 7230 5935 7234 5995
rect 7286 5935 7544 5995
rect 7596 5935 7600 5995
rect 7230 5925 7600 5935
rect 7630 5995 8000 6080
rect 7630 5935 7634 5995
rect 7686 5935 7944 5995
rect 7996 5935 8000 5995
rect 7630 5925 8000 5935
rect 8030 5995 8400 6080
rect 8030 5935 8034 5995
rect 8086 5935 8344 5995
rect 8396 5935 8400 5995
rect 8030 5925 8400 5935
rect 8430 5995 8800 6080
rect 8430 5935 8434 5995
rect 8486 5935 8744 5995
rect 8796 5935 8800 5995
rect 8430 5925 8800 5935
rect 8830 5995 9200 6080
rect 8830 5935 8834 5995
rect 8886 5935 9144 5995
rect 9196 5935 9200 5995
rect 8830 5925 9200 5935
rect 9230 5995 9600 6080
rect 9230 5935 9234 5995
rect 9286 5935 9544 5995
rect 9596 5935 9600 5995
rect 9230 5925 9600 5935
rect 9630 5995 10000 6080
rect 9630 5935 9634 5995
rect 9686 5935 9944 5995
rect 9996 5935 10000 5995
rect 9630 5925 10000 5935
rect 10030 5995 10400 6080
rect 10030 5935 10034 5995
rect 10086 5935 10344 5995
rect 10396 5935 10400 5995
rect 10030 5925 10400 5935
rect 10430 5995 10800 6080
rect 10430 5935 10434 5995
rect 10486 5935 10744 5995
rect 10796 5935 10800 5995
rect 10430 5925 10800 5935
rect 10830 5995 11200 6080
rect 10830 5935 10834 5995
rect 10886 5935 11144 5995
rect 11196 5935 11200 5995
rect 10830 5925 11200 5935
rect 11230 5995 11600 6080
rect 11230 5935 11234 5995
rect 11286 5935 11544 5995
rect 11596 5935 11600 5995
rect 11230 5925 11600 5935
rect 11630 5995 12000 6080
rect 11630 5935 11634 5995
rect 11686 5935 11944 5995
rect 11996 5935 12000 5995
rect 11630 5925 12000 5935
rect 12030 5995 12400 6080
rect 12030 5935 12034 5995
rect 12086 5935 12344 5995
rect 12396 5935 12400 5995
rect 12030 5925 12400 5935
rect 12430 5995 12800 6080
rect 12430 5935 12434 5995
rect 12486 5935 12744 5995
rect 12796 5935 12800 5995
rect 12430 5925 12800 5935
rect 12830 5995 13200 6080
rect 12830 5935 12834 5995
rect 12886 5935 13144 5995
rect 13196 5935 13200 5995
rect 12830 5925 13200 5935
rect -330 5895 -324 5925
rect 30 5895 70 5925
rect 430 5895 470 5925
rect 830 5895 870 5925
rect 1230 5895 1270 5925
rect 1630 5895 1670 5925
rect 2030 5895 2070 5925
rect 2430 5895 2470 5925
rect 2830 5895 2870 5925
rect 3230 5895 3270 5925
rect 3630 5895 3670 5925
rect 4030 5895 4070 5925
rect 4430 5895 4470 5925
rect 4830 5895 4870 5925
rect 5230 5895 5270 5925
rect 5630 5895 5670 5925
rect 6030 5895 6070 5925
rect 6430 5895 6470 5925
rect 6830 5895 6870 5925
rect 7230 5895 7270 5925
rect 7630 5895 7670 5925
rect 8030 5895 8070 5925
rect 8430 5895 8470 5925
rect 8830 5895 8870 5925
rect 9230 5895 9270 5925
rect 9630 5895 9670 5925
rect 10030 5895 10070 5925
rect 10430 5895 10470 5925
rect 10830 5895 10870 5925
rect 11230 5895 11270 5925
rect 11630 5895 11670 5925
rect 12030 5895 12070 5925
rect 12430 5895 12470 5925
rect -330 5885 0 5895
rect -314 5825 -56 5885
rect -4 5825 0 5885
rect -330 5625 0 5825
rect -314 5565 -56 5625
rect -4 5565 0 5625
rect -330 5555 0 5565
rect 30 5885 400 5895
rect 30 5825 34 5885
rect 86 5825 344 5885
rect 396 5825 400 5885
rect 30 5750 400 5825
rect 430 5885 800 5895
rect 430 5825 434 5885
rect 486 5825 744 5885
rect 796 5825 800 5885
rect 430 5750 800 5825
rect 830 5885 1200 5895
rect 830 5825 834 5885
rect 886 5825 1144 5885
rect 1196 5825 1200 5885
rect 830 5750 1200 5825
rect 1230 5885 1600 5895
rect 1230 5825 1234 5885
rect 1286 5825 1544 5885
rect 1596 5825 1600 5885
rect 1230 5750 1600 5825
rect 1630 5885 2000 5895
rect 1630 5825 1634 5885
rect 1686 5825 1944 5885
rect 1996 5825 2000 5885
rect 1630 5750 2000 5825
rect 2030 5885 2400 5895
rect 2030 5825 2034 5885
rect 2086 5825 2344 5885
rect 2396 5825 2400 5885
rect 2030 5750 2400 5825
rect 2430 5885 2800 5895
rect 2430 5825 2434 5885
rect 2486 5825 2744 5885
rect 2796 5825 2800 5885
rect 2430 5750 2800 5825
rect 2830 5885 3200 5895
rect 2830 5825 2834 5885
rect 2886 5825 3144 5885
rect 3196 5825 3200 5885
rect 2830 5750 3200 5825
rect 30 5710 3200 5750
rect 30 5625 400 5710
rect 30 5565 34 5625
rect 86 5565 344 5625
rect 396 5565 400 5625
rect 30 5555 400 5565
rect 430 5625 800 5710
rect 430 5565 434 5625
rect 486 5565 744 5625
rect 796 5565 800 5625
rect 430 5555 800 5565
rect 830 5625 1200 5710
rect 830 5565 834 5625
rect 886 5565 1144 5625
rect 1196 5565 1200 5625
rect 830 5555 1200 5565
rect 1230 5625 1600 5710
rect 1230 5565 1234 5625
rect 1286 5565 1544 5625
rect 1596 5565 1600 5625
rect 1230 5555 1600 5565
rect 1630 5625 2000 5710
rect 1630 5565 1634 5625
rect 1686 5565 1944 5625
rect 1996 5565 2000 5625
rect 1630 5555 2000 5565
rect 2030 5625 2400 5710
rect 2030 5565 2034 5625
rect 2086 5565 2344 5625
rect 2396 5565 2400 5625
rect 2030 5555 2400 5565
rect 2430 5625 2800 5710
rect 2430 5565 2434 5625
rect 2486 5565 2744 5625
rect 2796 5565 2800 5625
rect 2430 5555 2800 5565
rect 2830 5625 3200 5710
rect 2830 5565 2834 5625
rect 2886 5565 3144 5625
rect 3196 5565 3200 5625
rect 2830 5555 3200 5565
rect 3230 5885 3600 5895
rect 3230 5825 3234 5885
rect 3286 5825 3544 5885
rect 3596 5825 3600 5885
rect 3230 5750 3600 5825
rect 3630 5885 4000 5895
rect 3630 5825 3634 5885
rect 3686 5825 3944 5885
rect 3996 5825 4000 5885
rect 3630 5750 4000 5825
rect 4030 5885 4400 5895
rect 4030 5825 4034 5885
rect 4086 5825 4344 5885
rect 4396 5825 4400 5885
rect 4030 5750 4400 5825
rect 4430 5885 4800 5895
rect 4430 5825 4434 5885
rect 4486 5825 4744 5885
rect 4796 5825 4800 5885
rect 4430 5750 4800 5825
rect 4830 5885 5200 5895
rect 4830 5825 4834 5885
rect 4886 5825 5144 5885
rect 5196 5825 5200 5885
rect 4830 5750 5200 5825
rect 5230 5885 5600 5895
rect 5230 5825 5234 5885
rect 5286 5825 5544 5885
rect 5596 5825 5600 5885
rect 5230 5750 5600 5825
rect 5630 5885 6000 5895
rect 5630 5825 5634 5885
rect 5686 5825 5944 5885
rect 5996 5825 6000 5885
rect 5630 5750 6000 5825
rect 6030 5885 6400 5895
rect 6030 5825 6034 5885
rect 6086 5825 6344 5885
rect 6396 5825 6400 5885
rect 6030 5750 6400 5825
rect 6430 5885 6800 5895
rect 6430 5825 6434 5885
rect 6486 5825 6744 5885
rect 6796 5825 6800 5885
rect 6430 5750 6800 5825
rect 6830 5885 7200 5895
rect 6830 5825 6834 5885
rect 6886 5825 7144 5885
rect 7196 5825 7200 5885
rect 6830 5750 7200 5825
rect 7230 5885 7600 5895
rect 7230 5825 7234 5885
rect 7286 5825 7544 5885
rect 7596 5825 7600 5885
rect 7230 5750 7600 5825
rect 7630 5885 8000 5895
rect 7630 5825 7634 5885
rect 7686 5825 7944 5885
rect 7996 5825 8000 5885
rect 7630 5750 8000 5825
rect 8030 5885 8400 5895
rect 8030 5825 8034 5885
rect 8086 5825 8344 5885
rect 8396 5825 8400 5885
rect 8030 5750 8400 5825
rect 8430 5885 8800 5895
rect 8430 5825 8434 5885
rect 8486 5825 8744 5885
rect 8796 5825 8800 5885
rect 8430 5750 8800 5825
rect 8830 5885 9200 5895
rect 8830 5825 8834 5885
rect 8886 5825 9144 5885
rect 9196 5825 9200 5885
rect 8830 5750 9200 5825
rect 9230 5885 9600 5895
rect 9230 5825 9234 5885
rect 9286 5825 9544 5885
rect 9596 5825 9600 5885
rect 9230 5750 9600 5825
rect 9630 5885 10000 5895
rect 9630 5825 9634 5885
rect 9686 5825 9944 5885
rect 9996 5825 10000 5885
rect 9630 5750 10000 5825
rect 10030 5885 10400 5895
rect 10030 5825 10034 5885
rect 10086 5825 10344 5885
rect 10396 5825 10400 5885
rect 10030 5750 10400 5825
rect 10430 5885 10800 5895
rect 10430 5825 10434 5885
rect 10486 5825 10744 5885
rect 10796 5825 10800 5885
rect 10430 5750 10800 5825
rect 10830 5885 11200 5895
rect 10830 5825 10834 5885
rect 10886 5825 11144 5885
rect 11196 5825 11200 5885
rect 10830 5750 11200 5825
rect 11230 5885 11600 5895
rect 11230 5825 11234 5885
rect 11286 5825 11544 5885
rect 11596 5825 11600 5885
rect 11230 5750 11600 5825
rect 11630 5885 12000 5895
rect 11630 5825 11634 5885
rect 11686 5825 11944 5885
rect 11996 5825 12000 5885
rect 11630 5750 12000 5825
rect 12030 5885 12400 5895
rect 12030 5825 12034 5885
rect 12086 5825 12344 5885
rect 12396 5825 12400 5885
rect 12030 5750 12400 5825
rect 12430 5885 12800 5895
rect 12430 5825 12434 5885
rect 12486 5825 12744 5885
rect 12796 5825 12800 5885
rect 12430 5750 12800 5825
rect 12830 5885 13200 5895
rect 12830 5825 12834 5885
rect 12886 5825 13144 5885
rect 13196 5825 13200 5885
rect 12830 5750 13200 5825
rect 3230 5710 13200 5750
rect 3230 5625 3600 5710
rect 3230 5565 3234 5625
rect 3286 5565 3544 5625
rect 3596 5565 3600 5625
rect 3230 5555 3600 5565
rect 3630 5625 4000 5710
rect 3630 5565 3634 5625
rect 3686 5565 3944 5625
rect 3996 5565 4000 5625
rect 3630 5555 4000 5565
rect 4030 5625 4400 5710
rect 4030 5565 4034 5625
rect 4086 5565 4344 5625
rect 4396 5565 4400 5625
rect 4030 5555 4400 5565
rect 4430 5625 4800 5710
rect 4430 5565 4434 5625
rect 4486 5565 4744 5625
rect 4796 5565 4800 5625
rect 4430 5555 4800 5565
rect 4830 5625 5200 5710
rect 4830 5565 4834 5625
rect 4886 5565 5144 5625
rect 5196 5565 5200 5625
rect 4830 5555 5200 5565
rect 5230 5625 5600 5710
rect 5230 5565 5234 5625
rect 5286 5565 5544 5625
rect 5596 5565 5600 5625
rect 5230 5555 5600 5565
rect 5630 5625 6000 5710
rect 5630 5565 5634 5625
rect 5686 5565 5944 5625
rect 5996 5565 6000 5625
rect 5630 5555 6000 5565
rect 6030 5625 6400 5710
rect 6030 5565 6034 5625
rect 6086 5565 6344 5625
rect 6396 5565 6400 5625
rect 6030 5555 6400 5565
rect 6430 5625 6800 5710
rect 6430 5565 6434 5625
rect 6486 5565 6744 5625
rect 6796 5565 6800 5625
rect 6430 5555 6800 5565
rect 6830 5625 7200 5710
rect 6830 5565 6834 5625
rect 6886 5565 7144 5625
rect 7196 5565 7200 5625
rect 6830 5555 7200 5565
rect 7230 5625 7600 5710
rect 7230 5565 7234 5625
rect 7286 5565 7544 5625
rect 7596 5565 7600 5625
rect 7230 5555 7600 5565
rect 7630 5625 8000 5710
rect 7630 5565 7634 5625
rect 7686 5565 7944 5625
rect 7996 5565 8000 5625
rect 7630 5555 8000 5565
rect 8030 5625 8400 5710
rect 8030 5565 8034 5625
rect 8086 5565 8344 5625
rect 8396 5565 8400 5625
rect 8030 5555 8400 5565
rect 8430 5625 8800 5710
rect 8430 5565 8434 5625
rect 8486 5565 8744 5625
rect 8796 5565 8800 5625
rect 8430 5555 8800 5565
rect 8830 5625 9200 5710
rect 8830 5565 8834 5625
rect 8886 5565 9144 5625
rect 9196 5565 9200 5625
rect 8830 5555 9200 5565
rect 9230 5625 9600 5710
rect 9230 5565 9234 5625
rect 9286 5565 9544 5625
rect 9596 5565 9600 5625
rect 9230 5555 9600 5565
rect 9630 5625 10000 5710
rect 9630 5565 9634 5625
rect 9686 5565 9944 5625
rect 9996 5565 10000 5625
rect 9630 5555 10000 5565
rect 10030 5625 10400 5710
rect 10030 5565 10034 5625
rect 10086 5565 10344 5625
rect 10396 5565 10400 5625
rect 10030 5555 10400 5565
rect 10430 5625 10800 5710
rect 10430 5565 10434 5625
rect 10486 5565 10744 5625
rect 10796 5565 10800 5625
rect 10430 5555 10800 5565
rect 10830 5625 11200 5710
rect 10830 5565 10834 5625
rect 10886 5565 11144 5625
rect 11196 5565 11200 5625
rect 10830 5555 11200 5565
rect 11230 5625 11600 5710
rect 11230 5565 11234 5625
rect 11286 5565 11544 5625
rect 11596 5565 11600 5625
rect 11230 5555 11600 5565
rect 11630 5625 12000 5710
rect 11630 5565 11634 5625
rect 11686 5565 11944 5625
rect 11996 5565 12000 5625
rect 11630 5555 12000 5565
rect 12030 5625 12400 5710
rect 12030 5565 12034 5625
rect 12086 5565 12344 5625
rect 12396 5565 12400 5625
rect 12030 5555 12400 5565
rect 12430 5625 12800 5710
rect 12430 5565 12434 5625
rect 12486 5565 12744 5625
rect 12796 5565 12800 5625
rect 12430 5555 12800 5565
rect 12830 5625 13200 5710
rect 12830 5565 12834 5625
rect 12886 5565 13144 5625
rect 13196 5565 13200 5625
rect 12830 5555 13200 5565
rect -330 5525 -324 5555
rect 30 5525 70 5555
rect 430 5525 470 5555
rect 830 5525 870 5555
rect 1230 5525 1270 5555
rect 1630 5525 1670 5555
rect 2030 5525 2070 5555
rect 2430 5525 2470 5555
rect 2830 5525 2870 5555
rect 3230 5525 3270 5555
rect 3630 5525 3670 5555
rect 4030 5525 4070 5555
rect 4430 5525 4470 5555
rect 4830 5525 4870 5555
rect 5230 5525 5270 5555
rect 5630 5525 5670 5555
rect 6030 5525 6070 5555
rect 6430 5525 6470 5555
rect 6830 5525 6870 5555
rect 7230 5525 7270 5555
rect 7630 5525 7670 5555
rect 8030 5525 8070 5555
rect 8430 5525 8470 5555
rect 8830 5525 8870 5555
rect 9230 5525 9270 5555
rect 9630 5525 9670 5555
rect 10030 5525 10070 5555
rect 10430 5525 10470 5555
rect 10830 5525 10870 5555
rect 11230 5525 11270 5555
rect 11630 5525 11670 5555
rect 12030 5525 12070 5555
rect 12430 5525 12470 5555
rect -330 5515 0 5525
rect -314 5455 -56 5515
rect -4 5455 0 5515
rect -330 5255 0 5455
rect -314 5195 -56 5255
rect -4 5195 0 5255
rect -330 5185 0 5195
rect 30 5515 400 5525
rect 30 5455 34 5515
rect 86 5455 344 5515
rect 396 5455 400 5515
rect 30 5380 400 5455
rect 430 5515 800 5525
rect 430 5455 434 5515
rect 486 5455 744 5515
rect 796 5455 800 5515
rect 430 5380 800 5455
rect 830 5515 1200 5525
rect 830 5455 834 5515
rect 886 5455 1144 5515
rect 1196 5455 1200 5515
rect 830 5380 1200 5455
rect 1230 5515 1600 5525
rect 1230 5455 1234 5515
rect 1286 5455 1544 5515
rect 1596 5455 1600 5515
rect 1230 5380 1600 5455
rect 1630 5515 2000 5525
rect 1630 5455 1634 5515
rect 1686 5455 1944 5515
rect 1996 5455 2000 5515
rect 1630 5380 2000 5455
rect 2030 5515 2400 5525
rect 2030 5455 2034 5515
rect 2086 5455 2344 5515
rect 2396 5455 2400 5515
rect 2030 5380 2400 5455
rect 2430 5515 2800 5525
rect 2430 5455 2434 5515
rect 2486 5455 2744 5515
rect 2796 5455 2800 5515
rect 2430 5380 2800 5455
rect 2830 5515 3200 5525
rect 2830 5455 2834 5515
rect 2886 5455 3144 5515
rect 3196 5455 3200 5515
rect 2830 5380 3200 5455
rect 30 5340 3200 5380
rect 30 5255 400 5340
rect 30 5195 34 5255
rect 86 5195 344 5255
rect 396 5195 400 5255
rect 30 5185 400 5195
rect 430 5255 800 5340
rect 430 5195 434 5255
rect 486 5195 744 5255
rect 796 5195 800 5255
rect 430 5185 800 5195
rect 830 5255 1200 5340
rect 830 5195 834 5255
rect 886 5195 1144 5255
rect 1196 5195 1200 5255
rect 830 5185 1200 5195
rect 1230 5255 1600 5340
rect 1230 5195 1234 5255
rect 1286 5195 1544 5255
rect 1596 5195 1600 5255
rect 1230 5185 1600 5195
rect 1630 5255 2000 5340
rect 1630 5195 1634 5255
rect 1686 5195 1944 5255
rect 1996 5195 2000 5255
rect 1630 5185 2000 5195
rect 2030 5255 2400 5340
rect 2030 5195 2034 5255
rect 2086 5195 2344 5255
rect 2396 5195 2400 5255
rect 2030 5185 2400 5195
rect 2430 5255 2800 5340
rect 2430 5195 2434 5255
rect 2486 5195 2744 5255
rect 2796 5195 2800 5255
rect 2430 5185 2800 5195
rect 2830 5255 3200 5340
rect 2830 5195 2834 5255
rect 2886 5195 3144 5255
rect 3196 5195 3200 5255
rect 2830 5185 3200 5195
rect 3230 5515 3600 5525
rect 3230 5455 3234 5515
rect 3286 5455 3544 5515
rect 3596 5455 3600 5515
rect 3230 5380 3600 5455
rect 3630 5515 4000 5525
rect 3630 5455 3634 5515
rect 3686 5455 3944 5515
rect 3996 5455 4000 5515
rect 3630 5380 4000 5455
rect 4030 5515 4400 5525
rect 4030 5455 4034 5515
rect 4086 5455 4344 5515
rect 4396 5455 4400 5515
rect 4030 5380 4400 5455
rect 4430 5515 4800 5525
rect 4430 5455 4434 5515
rect 4486 5455 4744 5515
rect 4796 5455 4800 5515
rect 4430 5380 4800 5455
rect 4830 5515 5200 5525
rect 4830 5455 4834 5515
rect 4886 5455 5144 5515
rect 5196 5455 5200 5515
rect 4830 5380 5200 5455
rect 5230 5515 5600 5525
rect 5230 5455 5234 5515
rect 5286 5455 5544 5515
rect 5596 5455 5600 5515
rect 5230 5380 5600 5455
rect 5630 5515 6000 5525
rect 5630 5455 5634 5515
rect 5686 5455 5944 5515
rect 5996 5455 6000 5515
rect 5630 5380 6000 5455
rect 6030 5515 6400 5525
rect 6030 5455 6034 5515
rect 6086 5455 6344 5515
rect 6396 5455 6400 5515
rect 6030 5380 6400 5455
rect 6430 5515 6800 5525
rect 6430 5455 6434 5515
rect 6486 5455 6744 5515
rect 6796 5455 6800 5515
rect 6430 5380 6800 5455
rect 6830 5515 7200 5525
rect 6830 5455 6834 5515
rect 6886 5455 7144 5515
rect 7196 5455 7200 5515
rect 6830 5380 7200 5455
rect 7230 5515 7600 5525
rect 7230 5455 7234 5515
rect 7286 5455 7544 5515
rect 7596 5455 7600 5515
rect 7230 5380 7600 5455
rect 7630 5515 8000 5525
rect 7630 5455 7634 5515
rect 7686 5455 7944 5515
rect 7996 5455 8000 5515
rect 7630 5380 8000 5455
rect 8030 5515 8400 5525
rect 8030 5455 8034 5515
rect 8086 5455 8344 5515
rect 8396 5455 8400 5515
rect 8030 5380 8400 5455
rect 8430 5515 8800 5525
rect 8430 5455 8434 5515
rect 8486 5455 8744 5515
rect 8796 5455 8800 5515
rect 8430 5380 8800 5455
rect 8830 5515 9200 5525
rect 8830 5455 8834 5515
rect 8886 5455 9144 5515
rect 9196 5455 9200 5515
rect 8830 5380 9200 5455
rect 9230 5515 9600 5525
rect 9230 5455 9234 5515
rect 9286 5455 9544 5515
rect 9596 5455 9600 5515
rect 9230 5380 9600 5455
rect 9630 5515 10000 5525
rect 9630 5455 9634 5515
rect 9686 5455 9944 5515
rect 9996 5455 10000 5515
rect 9630 5380 10000 5455
rect 10030 5515 10400 5525
rect 10030 5455 10034 5515
rect 10086 5455 10344 5515
rect 10396 5455 10400 5515
rect 10030 5380 10400 5455
rect 10430 5515 10800 5525
rect 10430 5455 10434 5515
rect 10486 5455 10744 5515
rect 10796 5455 10800 5515
rect 10430 5380 10800 5455
rect 10830 5515 11200 5525
rect 10830 5455 10834 5515
rect 10886 5455 11144 5515
rect 11196 5455 11200 5515
rect 10830 5380 11200 5455
rect 11230 5515 11600 5525
rect 11230 5455 11234 5515
rect 11286 5455 11544 5515
rect 11596 5455 11600 5515
rect 11230 5380 11600 5455
rect 11630 5515 12000 5525
rect 11630 5455 11634 5515
rect 11686 5455 11944 5515
rect 11996 5455 12000 5515
rect 11630 5380 12000 5455
rect 12030 5515 12400 5525
rect 12030 5455 12034 5515
rect 12086 5455 12344 5515
rect 12396 5455 12400 5515
rect 12030 5380 12400 5455
rect 12430 5515 12800 5525
rect 12430 5455 12434 5515
rect 12486 5455 12744 5515
rect 12796 5455 12800 5515
rect 12430 5380 12800 5455
rect 12830 5515 13200 5525
rect 12830 5455 12834 5515
rect 12886 5455 13144 5515
rect 13196 5455 13200 5515
rect 12830 5380 13200 5455
rect 3230 5340 13200 5380
rect 3230 5255 3600 5340
rect 3230 5195 3234 5255
rect 3286 5195 3544 5255
rect 3596 5195 3600 5255
rect 3230 5185 3600 5195
rect 3630 5255 4000 5340
rect 3630 5195 3634 5255
rect 3686 5195 3944 5255
rect 3996 5195 4000 5255
rect 3630 5185 4000 5195
rect 4030 5255 4400 5340
rect 4030 5195 4034 5255
rect 4086 5195 4344 5255
rect 4396 5195 4400 5255
rect 4030 5185 4400 5195
rect 4430 5255 4800 5340
rect 4430 5195 4434 5255
rect 4486 5195 4744 5255
rect 4796 5195 4800 5255
rect 4430 5185 4800 5195
rect 4830 5255 5200 5340
rect 4830 5195 4834 5255
rect 4886 5195 5144 5255
rect 5196 5195 5200 5255
rect 4830 5185 5200 5195
rect 5230 5255 5600 5340
rect 5230 5195 5234 5255
rect 5286 5195 5544 5255
rect 5596 5195 5600 5255
rect 5230 5185 5600 5195
rect 5630 5255 6000 5340
rect 5630 5195 5634 5255
rect 5686 5195 5944 5255
rect 5996 5195 6000 5255
rect 5630 5185 6000 5195
rect 6030 5255 6400 5340
rect 6030 5195 6034 5255
rect 6086 5195 6344 5255
rect 6396 5195 6400 5255
rect 6030 5185 6400 5195
rect 6430 5255 6800 5340
rect 6430 5195 6434 5255
rect 6486 5195 6744 5255
rect 6796 5195 6800 5255
rect 6430 5185 6800 5195
rect 6830 5255 7200 5340
rect 6830 5195 6834 5255
rect 6886 5195 7144 5255
rect 7196 5195 7200 5255
rect 6830 5185 7200 5195
rect 7230 5255 7600 5340
rect 7230 5195 7234 5255
rect 7286 5195 7544 5255
rect 7596 5195 7600 5255
rect 7230 5185 7600 5195
rect 7630 5255 8000 5340
rect 7630 5195 7634 5255
rect 7686 5195 7944 5255
rect 7996 5195 8000 5255
rect 7630 5185 8000 5195
rect 8030 5255 8400 5340
rect 8030 5195 8034 5255
rect 8086 5195 8344 5255
rect 8396 5195 8400 5255
rect 8030 5185 8400 5195
rect 8430 5255 8800 5340
rect 8430 5195 8434 5255
rect 8486 5195 8744 5255
rect 8796 5195 8800 5255
rect 8430 5185 8800 5195
rect 8830 5255 9200 5340
rect 8830 5195 8834 5255
rect 8886 5195 9144 5255
rect 9196 5195 9200 5255
rect 8830 5185 9200 5195
rect 9230 5255 9600 5340
rect 9230 5195 9234 5255
rect 9286 5195 9544 5255
rect 9596 5195 9600 5255
rect 9230 5185 9600 5195
rect 9630 5255 10000 5340
rect 9630 5195 9634 5255
rect 9686 5195 9944 5255
rect 9996 5195 10000 5255
rect 9630 5185 10000 5195
rect 10030 5255 10400 5340
rect 10030 5195 10034 5255
rect 10086 5195 10344 5255
rect 10396 5195 10400 5255
rect 10030 5185 10400 5195
rect 10430 5255 10800 5340
rect 10430 5195 10434 5255
rect 10486 5195 10744 5255
rect 10796 5195 10800 5255
rect 10430 5185 10800 5195
rect 10830 5255 11200 5340
rect 10830 5195 10834 5255
rect 10886 5195 11144 5255
rect 11196 5195 11200 5255
rect 10830 5185 11200 5195
rect 11230 5255 11600 5340
rect 11230 5195 11234 5255
rect 11286 5195 11544 5255
rect 11596 5195 11600 5255
rect 11230 5185 11600 5195
rect 11630 5255 12000 5340
rect 11630 5195 11634 5255
rect 11686 5195 11944 5255
rect 11996 5195 12000 5255
rect 11630 5185 12000 5195
rect 12030 5255 12400 5340
rect 12030 5195 12034 5255
rect 12086 5195 12344 5255
rect 12396 5195 12400 5255
rect 12030 5185 12400 5195
rect 12430 5255 12800 5340
rect 12430 5195 12434 5255
rect 12486 5195 12744 5255
rect 12796 5195 12800 5255
rect 12430 5185 12800 5195
rect 12830 5255 13200 5340
rect 12830 5195 12834 5255
rect 12886 5195 13144 5255
rect 13196 5195 13200 5255
rect 12830 5185 13200 5195
rect -330 5155 -324 5185
rect 30 5155 70 5185
rect 430 5155 470 5185
rect 830 5155 870 5185
rect 1230 5155 1270 5185
rect 1630 5155 1670 5185
rect 2030 5155 2070 5185
rect 2430 5155 2470 5185
rect 2830 5155 2870 5185
rect 3230 5155 3270 5185
rect 3630 5155 3670 5185
rect 4030 5155 4070 5185
rect 4430 5155 4470 5185
rect 4830 5155 4870 5185
rect 5230 5155 5270 5185
rect 5630 5155 5670 5185
rect 6030 5155 6070 5185
rect 6430 5155 6470 5185
rect 6830 5155 6870 5185
rect 7230 5155 7270 5185
rect 7630 5155 7670 5185
rect 8030 5155 8070 5185
rect 8430 5155 8470 5185
rect 8830 5155 8870 5185
rect 9230 5155 9270 5185
rect 9630 5155 9670 5185
rect 10030 5155 10070 5185
rect 10430 5155 10470 5185
rect 10830 5155 10870 5185
rect 11230 5155 11270 5185
rect 11630 5155 11670 5185
rect 12030 5155 12070 5185
rect 12430 5155 12470 5185
rect -330 5145 0 5155
rect -314 5085 -56 5145
rect -4 5085 0 5145
rect -330 4885 0 5085
rect -314 4825 -56 4885
rect -4 4825 0 4885
rect -330 4815 0 4825
rect 30 5145 400 5155
rect 30 5085 34 5145
rect 86 5085 344 5145
rect 396 5085 400 5145
rect 30 5010 400 5085
rect 430 5145 800 5155
rect 430 5085 434 5145
rect 486 5085 744 5145
rect 796 5085 800 5145
rect 430 5010 800 5085
rect 830 5145 1200 5155
rect 830 5085 834 5145
rect 886 5085 1144 5145
rect 1196 5085 1200 5145
rect 830 5010 1200 5085
rect 1230 5145 1600 5155
rect 1230 5085 1234 5145
rect 1286 5085 1544 5145
rect 1596 5085 1600 5145
rect 1230 5010 1600 5085
rect 1630 5145 2000 5155
rect 1630 5085 1634 5145
rect 1686 5085 1944 5145
rect 1996 5085 2000 5145
rect 1630 5010 2000 5085
rect 2030 5145 2400 5155
rect 2030 5085 2034 5145
rect 2086 5085 2344 5145
rect 2396 5085 2400 5145
rect 2030 5010 2400 5085
rect 2430 5145 2800 5155
rect 2430 5085 2434 5145
rect 2486 5085 2744 5145
rect 2796 5085 2800 5145
rect 2430 5010 2800 5085
rect 2830 5145 3200 5155
rect 2830 5085 2834 5145
rect 2886 5085 3144 5145
rect 3196 5085 3200 5145
rect 2830 5010 3200 5085
rect 30 4970 3200 5010
rect 30 4885 400 4970
rect 30 4825 34 4885
rect 86 4825 344 4885
rect 396 4825 400 4885
rect 30 4815 400 4825
rect 430 4885 800 4970
rect 430 4825 434 4885
rect 486 4825 744 4885
rect 796 4825 800 4885
rect 430 4815 800 4825
rect 830 4885 1200 4970
rect 830 4825 834 4885
rect 886 4825 1144 4885
rect 1196 4825 1200 4885
rect 830 4815 1200 4825
rect 1230 4885 1600 4970
rect 1230 4825 1234 4885
rect 1286 4825 1544 4885
rect 1596 4825 1600 4885
rect 1230 4815 1600 4825
rect 1630 4885 2000 4970
rect 1630 4825 1634 4885
rect 1686 4825 1944 4885
rect 1996 4825 2000 4885
rect 1630 4815 2000 4825
rect 2030 4885 2400 4970
rect 2030 4825 2034 4885
rect 2086 4825 2344 4885
rect 2396 4825 2400 4885
rect 2030 4815 2400 4825
rect 2430 4885 2800 4970
rect 2430 4825 2434 4885
rect 2486 4825 2744 4885
rect 2796 4825 2800 4885
rect 2430 4815 2800 4825
rect 2830 4885 3200 4970
rect 2830 4825 2834 4885
rect 2886 4825 3144 4885
rect 3196 4825 3200 4885
rect 2830 4815 3200 4825
rect 3230 5145 3600 5155
rect 3230 5085 3234 5145
rect 3286 5085 3544 5145
rect 3596 5085 3600 5145
rect 3230 5010 3600 5085
rect 3630 5145 4000 5155
rect 3630 5085 3634 5145
rect 3686 5085 3944 5145
rect 3996 5085 4000 5145
rect 3630 5010 4000 5085
rect 4030 5145 4400 5155
rect 4030 5085 4034 5145
rect 4086 5085 4344 5145
rect 4396 5085 4400 5145
rect 4030 5010 4400 5085
rect 4430 5145 4800 5155
rect 4430 5085 4434 5145
rect 4486 5085 4744 5145
rect 4796 5085 4800 5145
rect 4430 5010 4800 5085
rect 4830 5145 5200 5155
rect 4830 5085 4834 5145
rect 4886 5085 5144 5145
rect 5196 5085 5200 5145
rect 4830 5010 5200 5085
rect 5230 5145 5600 5155
rect 5230 5085 5234 5145
rect 5286 5085 5544 5145
rect 5596 5085 5600 5145
rect 5230 5010 5600 5085
rect 5630 5145 6000 5155
rect 5630 5085 5634 5145
rect 5686 5085 5944 5145
rect 5996 5085 6000 5145
rect 5630 5010 6000 5085
rect 6030 5145 6400 5155
rect 6030 5085 6034 5145
rect 6086 5085 6344 5145
rect 6396 5085 6400 5145
rect 6030 5010 6400 5085
rect 6430 5145 6800 5155
rect 6430 5085 6434 5145
rect 6486 5085 6744 5145
rect 6796 5085 6800 5145
rect 6430 5010 6800 5085
rect 6830 5145 7200 5155
rect 6830 5085 6834 5145
rect 6886 5085 7144 5145
rect 7196 5085 7200 5145
rect 6830 5010 7200 5085
rect 7230 5145 7600 5155
rect 7230 5085 7234 5145
rect 7286 5085 7544 5145
rect 7596 5085 7600 5145
rect 7230 5010 7600 5085
rect 7630 5145 8000 5155
rect 7630 5085 7634 5145
rect 7686 5085 7944 5145
rect 7996 5085 8000 5145
rect 7630 5010 8000 5085
rect 8030 5145 8400 5155
rect 8030 5085 8034 5145
rect 8086 5085 8344 5145
rect 8396 5085 8400 5145
rect 8030 5010 8400 5085
rect 8430 5145 8800 5155
rect 8430 5085 8434 5145
rect 8486 5085 8744 5145
rect 8796 5085 8800 5145
rect 8430 5010 8800 5085
rect 8830 5145 9200 5155
rect 8830 5085 8834 5145
rect 8886 5085 9144 5145
rect 9196 5085 9200 5145
rect 8830 5010 9200 5085
rect 9230 5145 9600 5155
rect 9230 5085 9234 5145
rect 9286 5085 9544 5145
rect 9596 5085 9600 5145
rect 9230 5010 9600 5085
rect 9630 5145 10000 5155
rect 9630 5085 9634 5145
rect 9686 5085 9944 5145
rect 9996 5085 10000 5145
rect 9630 5010 10000 5085
rect 10030 5145 10400 5155
rect 10030 5085 10034 5145
rect 10086 5085 10344 5145
rect 10396 5085 10400 5145
rect 10030 5010 10400 5085
rect 10430 5145 10800 5155
rect 10430 5085 10434 5145
rect 10486 5085 10744 5145
rect 10796 5085 10800 5145
rect 10430 5010 10800 5085
rect 10830 5145 11200 5155
rect 10830 5085 10834 5145
rect 10886 5085 11144 5145
rect 11196 5085 11200 5145
rect 10830 5010 11200 5085
rect 11230 5145 11600 5155
rect 11230 5085 11234 5145
rect 11286 5085 11544 5145
rect 11596 5085 11600 5145
rect 11230 5010 11600 5085
rect 11630 5145 12000 5155
rect 11630 5085 11634 5145
rect 11686 5085 11944 5145
rect 11996 5085 12000 5145
rect 11630 5010 12000 5085
rect 12030 5145 12400 5155
rect 12030 5085 12034 5145
rect 12086 5085 12344 5145
rect 12396 5085 12400 5145
rect 12030 5010 12400 5085
rect 12430 5145 12800 5155
rect 12430 5085 12434 5145
rect 12486 5085 12744 5145
rect 12796 5085 12800 5145
rect 12430 5010 12800 5085
rect 12830 5145 13200 5155
rect 12830 5085 12834 5145
rect 12886 5085 13144 5145
rect 13196 5085 13200 5145
rect 12830 5010 13200 5085
rect 3230 4970 13200 5010
rect 3230 4885 3600 4970
rect 3230 4825 3234 4885
rect 3286 4825 3544 4885
rect 3596 4825 3600 4885
rect 3230 4815 3600 4825
rect 3630 4885 4000 4970
rect 3630 4825 3634 4885
rect 3686 4825 3944 4885
rect 3996 4825 4000 4885
rect 3630 4815 4000 4825
rect 4030 4885 4400 4970
rect 4030 4825 4034 4885
rect 4086 4825 4344 4885
rect 4396 4825 4400 4885
rect 4030 4815 4400 4825
rect 4430 4885 4800 4970
rect 4430 4825 4434 4885
rect 4486 4825 4744 4885
rect 4796 4825 4800 4885
rect 4430 4815 4800 4825
rect 4830 4885 5200 4970
rect 4830 4825 4834 4885
rect 4886 4825 5144 4885
rect 5196 4825 5200 4885
rect 4830 4815 5200 4825
rect 5230 4885 5600 4970
rect 5230 4825 5234 4885
rect 5286 4825 5544 4885
rect 5596 4825 5600 4885
rect 5230 4815 5600 4825
rect 5630 4885 6000 4970
rect 5630 4825 5634 4885
rect 5686 4825 5944 4885
rect 5996 4825 6000 4885
rect 5630 4815 6000 4825
rect 6030 4885 6400 4970
rect 6030 4825 6034 4885
rect 6086 4825 6344 4885
rect 6396 4825 6400 4885
rect 6030 4815 6400 4825
rect 6430 4885 6800 4970
rect 6430 4825 6434 4885
rect 6486 4825 6744 4885
rect 6796 4825 6800 4885
rect 6430 4815 6800 4825
rect 6830 4885 7200 4970
rect 6830 4825 6834 4885
rect 6886 4825 7144 4885
rect 7196 4825 7200 4885
rect 6830 4815 7200 4825
rect 7230 4885 7600 4970
rect 7230 4825 7234 4885
rect 7286 4825 7544 4885
rect 7596 4825 7600 4885
rect 7230 4815 7600 4825
rect 7630 4885 8000 4970
rect 7630 4825 7634 4885
rect 7686 4825 7944 4885
rect 7996 4825 8000 4885
rect 7630 4815 8000 4825
rect 8030 4885 8400 4970
rect 8030 4825 8034 4885
rect 8086 4825 8344 4885
rect 8396 4825 8400 4885
rect 8030 4815 8400 4825
rect 8430 4885 8800 4970
rect 8430 4825 8434 4885
rect 8486 4825 8744 4885
rect 8796 4825 8800 4885
rect 8430 4815 8800 4825
rect 8830 4885 9200 4970
rect 8830 4825 8834 4885
rect 8886 4825 9144 4885
rect 9196 4825 9200 4885
rect 8830 4815 9200 4825
rect 9230 4885 9600 4970
rect 9230 4825 9234 4885
rect 9286 4825 9544 4885
rect 9596 4825 9600 4885
rect 9230 4815 9600 4825
rect 9630 4885 10000 4970
rect 9630 4825 9634 4885
rect 9686 4825 9944 4885
rect 9996 4825 10000 4885
rect 9630 4815 10000 4825
rect 10030 4885 10400 4970
rect 10030 4825 10034 4885
rect 10086 4825 10344 4885
rect 10396 4825 10400 4885
rect 10030 4815 10400 4825
rect 10430 4885 10800 4970
rect 10430 4825 10434 4885
rect 10486 4825 10744 4885
rect 10796 4825 10800 4885
rect 10430 4815 10800 4825
rect 10830 4885 11200 4970
rect 10830 4825 10834 4885
rect 10886 4825 11144 4885
rect 11196 4825 11200 4885
rect 10830 4815 11200 4825
rect 11230 4885 11600 4970
rect 11230 4825 11234 4885
rect 11286 4825 11544 4885
rect 11596 4825 11600 4885
rect 11230 4815 11600 4825
rect 11630 4885 12000 4970
rect 11630 4825 11634 4885
rect 11686 4825 11944 4885
rect 11996 4825 12000 4885
rect 11630 4815 12000 4825
rect 12030 4885 12400 4970
rect 12030 4825 12034 4885
rect 12086 4825 12344 4885
rect 12396 4825 12400 4885
rect 12030 4815 12400 4825
rect 12430 4885 12800 4970
rect 12430 4825 12434 4885
rect 12486 4825 12744 4885
rect 12796 4825 12800 4885
rect 12430 4815 12800 4825
rect 12830 4885 13200 4970
rect 12830 4825 12834 4885
rect 12886 4825 13144 4885
rect 13196 4825 13200 4885
rect 12830 4815 13200 4825
rect -330 4785 -324 4815
rect 30 4785 70 4815
rect 430 4785 470 4815
rect 830 4785 870 4815
rect 1230 4785 1270 4815
rect 1630 4785 1670 4815
rect 2030 4785 2070 4815
rect 2430 4785 2470 4815
rect 2830 4785 2870 4815
rect 3230 4785 3270 4815
rect 3630 4785 3670 4815
rect 4030 4785 4070 4815
rect 4430 4785 4470 4815
rect 4830 4785 4870 4815
rect 5230 4785 5270 4815
rect 5630 4785 5670 4815
rect 6030 4785 6070 4815
rect 6430 4785 6470 4815
rect 6830 4785 6870 4815
rect 7230 4785 7270 4815
rect 7630 4785 7670 4815
rect 8030 4785 8070 4815
rect 8430 4785 8470 4815
rect 8830 4785 8870 4815
rect 9230 4785 9270 4815
rect 9630 4785 9670 4815
rect 10030 4785 10070 4815
rect 10430 4785 10470 4815
rect 10830 4785 10870 4815
rect 11230 4785 11270 4815
rect 11630 4785 11670 4815
rect 12030 4785 12070 4815
rect 12430 4785 12470 4815
rect -330 4775 0 4785
rect -314 4715 -56 4775
rect -4 4715 0 4775
rect -330 4515 0 4715
rect -314 4455 -56 4515
rect -4 4455 0 4515
rect -330 4445 0 4455
rect 30 4775 400 4785
rect 30 4715 34 4775
rect 86 4715 344 4775
rect 396 4715 400 4775
rect 30 4640 400 4715
rect 430 4775 800 4785
rect 430 4715 434 4775
rect 486 4715 744 4775
rect 796 4715 800 4775
rect 430 4640 800 4715
rect 830 4775 1200 4785
rect 830 4715 834 4775
rect 886 4715 1144 4775
rect 1196 4715 1200 4775
rect 830 4640 1200 4715
rect 1230 4775 1600 4785
rect 1230 4715 1234 4775
rect 1286 4715 1544 4775
rect 1596 4715 1600 4775
rect 1230 4640 1600 4715
rect 1630 4775 2000 4785
rect 1630 4715 1634 4775
rect 1686 4715 1944 4775
rect 1996 4715 2000 4775
rect 1630 4640 2000 4715
rect 2030 4775 2400 4785
rect 2030 4715 2034 4775
rect 2086 4715 2344 4775
rect 2396 4715 2400 4775
rect 2030 4640 2400 4715
rect 2430 4775 2800 4785
rect 2430 4715 2434 4775
rect 2486 4715 2744 4775
rect 2796 4715 2800 4775
rect 2430 4640 2800 4715
rect 2830 4775 3200 4785
rect 2830 4715 2834 4775
rect 2886 4715 3144 4775
rect 3196 4715 3200 4775
rect 2830 4640 3200 4715
rect 30 4600 3200 4640
rect 30 4515 400 4600
rect 30 4455 34 4515
rect 86 4455 344 4515
rect 396 4455 400 4515
rect 30 4445 400 4455
rect 430 4515 800 4600
rect 430 4455 434 4515
rect 486 4455 744 4515
rect 796 4455 800 4515
rect 430 4445 800 4455
rect 830 4515 1200 4600
rect 830 4455 834 4515
rect 886 4455 1144 4515
rect 1196 4455 1200 4515
rect 830 4445 1200 4455
rect 1230 4515 1600 4600
rect 1230 4455 1234 4515
rect 1286 4455 1544 4515
rect 1596 4455 1600 4515
rect 1230 4445 1600 4455
rect 1630 4515 2000 4600
rect 1630 4455 1634 4515
rect 1686 4455 1944 4515
rect 1996 4455 2000 4515
rect 1630 4445 2000 4455
rect 2030 4515 2400 4600
rect 2030 4455 2034 4515
rect 2086 4455 2344 4515
rect 2396 4455 2400 4515
rect 2030 4445 2400 4455
rect 2430 4515 2800 4600
rect 2430 4455 2434 4515
rect 2486 4455 2744 4515
rect 2796 4455 2800 4515
rect 2430 4445 2800 4455
rect 2830 4515 3200 4600
rect 2830 4455 2834 4515
rect 2886 4455 3144 4515
rect 3196 4455 3200 4515
rect 2830 4445 3200 4455
rect 3230 4775 3600 4785
rect 3230 4715 3234 4775
rect 3286 4715 3544 4775
rect 3596 4715 3600 4775
rect 3230 4640 3600 4715
rect 3630 4775 4000 4785
rect 3630 4715 3634 4775
rect 3686 4715 3944 4775
rect 3996 4715 4000 4775
rect 3630 4640 4000 4715
rect 4030 4775 4400 4785
rect 4030 4715 4034 4775
rect 4086 4715 4344 4775
rect 4396 4715 4400 4775
rect 4030 4640 4400 4715
rect 4430 4775 4800 4785
rect 4430 4715 4434 4775
rect 4486 4715 4744 4775
rect 4796 4715 4800 4775
rect 4430 4640 4800 4715
rect 4830 4775 5200 4785
rect 4830 4715 4834 4775
rect 4886 4715 5144 4775
rect 5196 4715 5200 4775
rect 4830 4640 5200 4715
rect 5230 4775 5600 4785
rect 5230 4715 5234 4775
rect 5286 4715 5544 4775
rect 5596 4715 5600 4775
rect 5230 4640 5600 4715
rect 5630 4775 6000 4785
rect 5630 4715 5634 4775
rect 5686 4715 5944 4775
rect 5996 4715 6000 4775
rect 5630 4640 6000 4715
rect 6030 4775 6400 4785
rect 6030 4715 6034 4775
rect 6086 4715 6344 4775
rect 6396 4715 6400 4775
rect 6030 4640 6400 4715
rect 6430 4775 6800 4785
rect 6430 4715 6434 4775
rect 6486 4715 6744 4775
rect 6796 4715 6800 4775
rect 6430 4640 6800 4715
rect 6830 4775 7200 4785
rect 6830 4715 6834 4775
rect 6886 4715 7144 4775
rect 7196 4715 7200 4775
rect 6830 4640 7200 4715
rect 7230 4775 7600 4785
rect 7230 4715 7234 4775
rect 7286 4715 7544 4775
rect 7596 4715 7600 4775
rect 7230 4640 7600 4715
rect 7630 4775 8000 4785
rect 7630 4715 7634 4775
rect 7686 4715 7944 4775
rect 7996 4715 8000 4775
rect 7630 4640 8000 4715
rect 8030 4775 8400 4785
rect 8030 4715 8034 4775
rect 8086 4715 8344 4775
rect 8396 4715 8400 4775
rect 8030 4640 8400 4715
rect 8430 4775 8800 4785
rect 8430 4715 8434 4775
rect 8486 4715 8744 4775
rect 8796 4715 8800 4775
rect 8430 4640 8800 4715
rect 8830 4775 9200 4785
rect 8830 4715 8834 4775
rect 8886 4715 9144 4775
rect 9196 4715 9200 4775
rect 8830 4640 9200 4715
rect 9230 4775 9600 4785
rect 9230 4715 9234 4775
rect 9286 4715 9544 4775
rect 9596 4715 9600 4775
rect 9230 4640 9600 4715
rect 9630 4775 10000 4785
rect 9630 4715 9634 4775
rect 9686 4715 9944 4775
rect 9996 4715 10000 4775
rect 9630 4640 10000 4715
rect 10030 4775 10400 4785
rect 10030 4715 10034 4775
rect 10086 4715 10344 4775
rect 10396 4715 10400 4775
rect 10030 4640 10400 4715
rect 10430 4775 10800 4785
rect 10430 4715 10434 4775
rect 10486 4715 10744 4775
rect 10796 4715 10800 4775
rect 10430 4640 10800 4715
rect 10830 4775 11200 4785
rect 10830 4715 10834 4775
rect 10886 4715 11144 4775
rect 11196 4715 11200 4775
rect 10830 4640 11200 4715
rect 11230 4775 11600 4785
rect 11230 4715 11234 4775
rect 11286 4715 11544 4775
rect 11596 4715 11600 4775
rect 11230 4640 11600 4715
rect 11630 4775 12000 4785
rect 11630 4715 11634 4775
rect 11686 4715 11944 4775
rect 11996 4715 12000 4775
rect 11630 4640 12000 4715
rect 12030 4775 12400 4785
rect 12030 4715 12034 4775
rect 12086 4715 12344 4775
rect 12396 4715 12400 4775
rect 12030 4640 12400 4715
rect 12430 4775 12800 4785
rect 12430 4715 12434 4775
rect 12486 4715 12744 4775
rect 12796 4715 12800 4775
rect 12430 4640 12800 4715
rect 12830 4775 13200 4785
rect 12830 4715 12834 4775
rect 12886 4715 13144 4775
rect 13196 4715 13200 4775
rect 12830 4640 13200 4715
rect 3230 4600 13200 4640
rect 3230 4515 3600 4600
rect 3230 4455 3234 4515
rect 3286 4455 3544 4515
rect 3596 4455 3600 4515
rect 3230 4445 3600 4455
rect 3630 4515 4000 4600
rect 3630 4455 3634 4515
rect 3686 4455 3944 4515
rect 3996 4455 4000 4515
rect 3630 4445 4000 4455
rect 4030 4515 4400 4600
rect 4030 4455 4034 4515
rect 4086 4455 4344 4515
rect 4396 4455 4400 4515
rect 4030 4445 4400 4455
rect 4430 4515 4800 4600
rect 4430 4455 4434 4515
rect 4486 4455 4744 4515
rect 4796 4455 4800 4515
rect 4430 4445 4800 4455
rect 4830 4515 5200 4600
rect 4830 4455 4834 4515
rect 4886 4455 5144 4515
rect 5196 4455 5200 4515
rect 4830 4445 5200 4455
rect 5230 4515 5600 4600
rect 5230 4455 5234 4515
rect 5286 4455 5544 4515
rect 5596 4455 5600 4515
rect 5230 4445 5600 4455
rect 5630 4515 6000 4600
rect 5630 4455 5634 4515
rect 5686 4455 5944 4515
rect 5996 4455 6000 4515
rect 5630 4445 6000 4455
rect 6030 4515 6400 4600
rect 6030 4455 6034 4515
rect 6086 4455 6344 4515
rect 6396 4455 6400 4515
rect 6030 4445 6400 4455
rect 6430 4515 6800 4600
rect 6430 4455 6434 4515
rect 6486 4455 6744 4515
rect 6796 4455 6800 4515
rect 6430 4445 6800 4455
rect 6830 4515 7200 4600
rect 6830 4455 6834 4515
rect 6886 4455 7144 4515
rect 7196 4455 7200 4515
rect 6830 4445 7200 4455
rect 7230 4515 7600 4600
rect 7230 4455 7234 4515
rect 7286 4455 7544 4515
rect 7596 4455 7600 4515
rect 7230 4445 7600 4455
rect 7630 4515 8000 4600
rect 7630 4455 7634 4515
rect 7686 4455 7944 4515
rect 7996 4455 8000 4515
rect 7630 4445 8000 4455
rect 8030 4515 8400 4600
rect 8030 4455 8034 4515
rect 8086 4455 8344 4515
rect 8396 4455 8400 4515
rect 8030 4445 8400 4455
rect 8430 4515 8800 4600
rect 8430 4455 8434 4515
rect 8486 4455 8744 4515
rect 8796 4455 8800 4515
rect 8430 4445 8800 4455
rect 8830 4515 9200 4600
rect 8830 4455 8834 4515
rect 8886 4455 9144 4515
rect 9196 4455 9200 4515
rect 8830 4445 9200 4455
rect 9230 4515 9600 4600
rect 9230 4455 9234 4515
rect 9286 4455 9544 4515
rect 9596 4455 9600 4515
rect 9230 4445 9600 4455
rect 9630 4515 10000 4600
rect 9630 4455 9634 4515
rect 9686 4455 9944 4515
rect 9996 4455 10000 4515
rect 9630 4445 10000 4455
rect 10030 4515 10400 4600
rect 10030 4455 10034 4515
rect 10086 4455 10344 4515
rect 10396 4455 10400 4515
rect 10030 4445 10400 4455
rect 10430 4515 10800 4600
rect 10430 4455 10434 4515
rect 10486 4455 10744 4515
rect 10796 4455 10800 4515
rect 10430 4445 10800 4455
rect 10830 4515 11200 4600
rect 10830 4455 10834 4515
rect 10886 4455 11144 4515
rect 11196 4455 11200 4515
rect 10830 4445 11200 4455
rect 11230 4515 11600 4600
rect 11230 4455 11234 4515
rect 11286 4455 11544 4515
rect 11596 4455 11600 4515
rect 11230 4445 11600 4455
rect 11630 4515 12000 4600
rect 11630 4455 11634 4515
rect 11686 4455 11944 4515
rect 11996 4455 12000 4515
rect 11630 4445 12000 4455
rect 12030 4515 12400 4600
rect 12030 4455 12034 4515
rect 12086 4455 12344 4515
rect 12396 4455 12400 4515
rect 12030 4445 12400 4455
rect 12430 4515 12800 4600
rect 12430 4455 12434 4515
rect 12486 4455 12744 4515
rect 12796 4455 12800 4515
rect 12430 4445 12800 4455
rect 12830 4515 13200 4600
rect 12830 4455 12834 4515
rect 12886 4455 13144 4515
rect 13196 4455 13200 4515
rect 12830 4445 13200 4455
rect -330 4415 -324 4445
rect 30 4415 70 4445
rect 430 4415 470 4445
rect 830 4415 870 4445
rect 1230 4415 1270 4445
rect 1630 4415 1670 4445
rect 2030 4415 2070 4445
rect 2430 4415 2470 4445
rect 2830 4415 2870 4445
rect 3230 4415 3270 4445
rect 3630 4415 3670 4445
rect 4030 4415 4070 4445
rect 4430 4415 4470 4445
rect 4830 4415 4870 4445
rect 5230 4415 5270 4445
rect 5630 4415 5670 4445
rect 6030 4415 6070 4445
rect 6430 4415 6470 4445
rect 6830 4415 6870 4445
rect 7230 4415 7270 4445
rect 7630 4415 7670 4445
rect 8030 4415 8070 4445
rect 8430 4415 8470 4445
rect 8830 4415 8870 4445
rect 9230 4415 9270 4445
rect 9630 4415 9670 4445
rect 10030 4415 10070 4445
rect 10430 4415 10470 4445
rect 10830 4415 10870 4445
rect 11230 4415 11270 4445
rect 11630 4415 11670 4445
rect 12030 4415 12070 4445
rect 12430 4415 12470 4445
rect -330 4405 0 4415
rect -314 4345 -56 4405
rect -4 4345 0 4405
rect -330 4145 0 4345
rect -314 4085 -56 4145
rect -4 4085 0 4145
rect -330 4075 0 4085
rect 30 4405 400 4415
rect 30 4345 34 4405
rect 86 4345 344 4405
rect 396 4345 400 4405
rect 30 4270 400 4345
rect 430 4405 800 4415
rect 430 4345 434 4405
rect 486 4345 744 4405
rect 796 4345 800 4405
rect 430 4270 800 4345
rect 830 4405 1200 4415
rect 830 4345 834 4405
rect 886 4345 1144 4405
rect 1196 4345 1200 4405
rect 830 4270 1200 4345
rect 1230 4405 1600 4415
rect 1230 4345 1234 4405
rect 1286 4345 1544 4405
rect 1596 4345 1600 4405
rect 1230 4270 1600 4345
rect 1630 4405 2000 4415
rect 1630 4345 1634 4405
rect 1686 4345 1944 4405
rect 1996 4345 2000 4405
rect 1630 4270 2000 4345
rect 2030 4405 2400 4415
rect 2030 4345 2034 4405
rect 2086 4345 2344 4405
rect 2396 4345 2400 4405
rect 2030 4270 2400 4345
rect 2430 4405 2800 4415
rect 2430 4345 2434 4405
rect 2486 4345 2744 4405
rect 2796 4345 2800 4405
rect 2430 4270 2800 4345
rect 2830 4405 3200 4415
rect 2830 4345 2834 4405
rect 2886 4345 3144 4405
rect 3196 4345 3200 4405
rect 2830 4270 3200 4345
rect 30 4230 3200 4270
rect 30 4145 400 4230
rect 30 4085 34 4145
rect 86 4085 344 4145
rect 396 4085 400 4145
rect 30 4075 400 4085
rect 430 4145 800 4230
rect 430 4085 434 4145
rect 486 4085 744 4145
rect 796 4085 800 4145
rect 430 4075 800 4085
rect 830 4145 1200 4230
rect 830 4085 834 4145
rect 886 4085 1144 4145
rect 1196 4085 1200 4145
rect 830 4075 1200 4085
rect 1230 4145 1600 4230
rect 1230 4085 1234 4145
rect 1286 4085 1544 4145
rect 1596 4085 1600 4145
rect 1230 4075 1600 4085
rect 1630 4145 2000 4230
rect 1630 4085 1634 4145
rect 1686 4085 1944 4145
rect 1996 4085 2000 4145
rect 1630 4075 2000 4085
rect 2030 4145 2400 4230
rect 2030 4085 2034 4145
rect 2086 4085 2344 4145
rect 2396 4085 2400 4145
rect 2030 4075 2400 4085
rect 2430 4145 2800 4230
rect 2430 4085 2434 4145
rect 2486 4085 2744 4145
rect 2796 4085 2800 4145
rect 2430 4075 2800 4085
rect 2830 4145 3200 4230
rect 2830 4085 2834 4145
rect 2886 4085 3144 4145
rect 3196 4085 3200 4145
rect 2830 4075 3200 4085
rect 3230 4405 3600 4415
rect 3230 4345 3234 4405
rect 3286 4345 3544 4405
rect 3596 4345 3600 4405
rect 3230 4270 3600 4345
rect 3630 4405 4000 4415
rect 3630 4345 3634 4405
rect 3686 4345 3944 4405
rect 3996 4345 4000 4405
rect 3630 4270 4000 4345
rect 4030 4405 4400 4415
rect 4030 4345 4034 4405
rect 4086 4345 4344 4405
rect 4396 4345 4400 4405
rect 4030 4270 4400 4345
rect 4430 4405 4800 4415
rect 4430 4345 4434 4405
rect 4486 4345 4744 4405
rect 4796 4345 4800 4405
rect 4430 4270 4800 4345
rect 4830 4405 5200 4415
rect 4830 4345 4834 4405
rect 4886 4345 5144 4405
rect 5196 4345 5200 4405
rect 4830 4270 5200 4345
rect 5230 4405 5600 4415
rect 5230 4345 5234 4405
rect 5286 4345 5544 4405
rect 5596 4345 5600 4405
rect 5230 4270 5600 4345
rect 5630 4405 6000 4415
rect 5630 4345 5634 4405
rect 5686 4345 5944 4405
rect 5996 4345 6000 4405
rect 5630 4270 6000 4345
rect 6030 4405 6400 4415
rect 6030 4345 6034 4405
rect 6086 4345 6344 4405
rect 6396 4345 6400 4405
rect 6030 4270 6400 4345
rect 6430 4405 6800 4415
rect 6430 4345 6434 4405
rect 6486 4345 6744 4405
rect 6796 4345 6800 4405
rect 6430 4270 6800 4345
rect 6830 4405 7200 4415
rect 6830 4345 6834 4405
rect 6886 4345 7144 4405
rect 7196 4345 7200 4405
rect 6830 4270 7200 4345
rect 7230 4405 7600 4415
rect 7230 4345 7234 4405
rect 7286 4345 7544 4405
rect 7596 4345 7600 4405
rect 7230 4270 7600 4345
rect 7630 4405 8000 4415
rect 7630 4345 7634 4405
rect 7686 4345 7944 4405
rect 7996 4345 8000 4405
rect 7630 4270 8000 4345
rect 8030 4405 8400 4415
rect 8030 4345 8034 4405
rect 8086 4345 8344 4405
rect 8396 4345 8400 4405
rect 8030 4270 8400 4345
rect 8430 4405 8800 4415
rect 8430 4345 8434 4405
rect 8486 4345 8744 4405
rect 8796 4345 8800 4405
rect 8430 4270 8800 4345
rect 8830 4405 9200 4415
rect 8830 4345 8834 4405
rect 8886 4345 9144 4405
rect 9196 4345 9200 4405
rect 8830 4270 9200 4345
rect 9230 4405 9600 4415
rect 9230 4345 9234 4405
rect 9286 4345 9544 4405
rect 9596 4345 9600 4405
rect 9230 4270 9600 4345
rect 9630 4405 10000 4415
rect 9630 4345 9634 4405
rect 9686 4345 9944 4405
rect 9996 4345 10000 4405
rect 9630 4270 10000 4345
rect 10030 4405 10400 4415
rect 10030 4345 10034 4405
rect 10086 4345 10344 4405
rect 10396 4345 10400 4405
rect 10030 4270 10400 4345
rect 10430 4405 10800 4415
rect 10430 4345 10434 4405
rect 10486 4345 10744 4405
rect 10796 4345 10800 4405
rect 10430 4270 10800 4345
rect 10830 4405 11200 4415
rect 10830 4345 10834 4405
rect 10886 4345 11144 4405
rect 11196 4345 11200 4405
rect 10830 4270 11200 4345
rect 11230 4405 11600 4415
rect 11230 4345 11234 4405
rect 11286 4345 11544 4405
rect 11596 4345 11600 4405
rect 11230 4270 11600 4345
rect 11630 4405 12000 4415
rect 11630 4345 11634 4405
rect 11686 4345 11944 4405
rect 11996 4345 12000 4405
rect 11630 4270 12000 4345
rect 12030 4405 12400 4415
rect 12030 4345 12034 4405
rect 12086 4345 12344 4405
rect 12396 4345 12400 4405
rect 12030 4270 12400 4345
rect 12430 4405 12800 4415
rect 12430 4345 12434 4405
rect 12486 4345 12744 4405
rect 12796 4345 12800 4405
rect 12430 4270 12800 4345
rect 12830 4405 13200 4415
rect 12830 4345 12834 4405
rect 12886 4345 13144 4405
rect 13196 4345 13200 4405
rect 12830 4270 13200 4345
rect 3230 4230 13200 4270
rect 3230 4145 3600 4230
rect 3230 4085 3234 4145
rect 3286 4085 3544 4145
rect 3596 4085 3600 4145
rect 3230 4075 3600 4085
rect 3630 4145 4000 4230
rect 3630 4085 3634 4145
rect 3686 4085 3944 4145
rect 3996 4085 4000 4145
rect 3630 4075 4000 4085
rect 4030 4145 4400 4230
rect 4030 4085 4034 4145
rect 4086 4085 4344 4145
rect 4396 4085 4400 4145
rect 4030 4075 4400 4085
rect 4430 4145 4800 4230
rect 4430 4085 4434 4145
rect 4486 4085 4744 4145
rect 4796 4085 4800 4145
rect 4430 4075 4800 4085
rect 4830 4145 5200 4230
rect 4830 4085 4834 4145
rect 4886 4085 5144 4145
rect 5196 4085 5200 4145
rect 4830 4075 5200 4085
rect 5230 4145 5600 4230
rect 5230 4085 5234 4145
rect 5286 4085 5544 4145
rect 5596 4085 5600 4145
rect 5230 4075 5600 4085
rect 5630 4145 6000 4230
rect 5630 4085 5634 4145
rect 5686 4085 5944 4145
rect 5996 4085 6000 4145
rect 5630 4075 6000 4085
rect 6030 4145 6400 4230
rect 6030 4085 6034 4145
rect 6086 4085 6344 4145
rect 6396 4085 6400 4145
rect 6030 4075 6400 4085
rect 6430 4145 6800 4230
rect 6430 4085 6434 4145
rect 6486 4085 6744 4145
rect 6796 4085 6800 4145
rect 6430 4075 6800 4085
rect 6830 4145 7200 4230
rect 6830 4085 6834 4145
rect 6886 4085 7144 4145
rect 7196 4085 7200 4145
rect 6830 4075 7200 4085
rect 7230 4145 7600 4230
rect 7230 4085 7234 4145
rect 7286 4085 7544 4145
rect 7596 4085 7600 4145
rect 7230 4075 7600 4085
rect 7630 4145 8000 4230
rect 7630 4085 7634 4145
rect 7686 4085 7944 4145
rect 7996 4085 8000 4145
rect 7630 4075 8000 4085
rect 8030 4145 8400 4230
rect 8030 4085 8034 4145
rect 8086 4085 8344 4145
rect 8396 4085 8400 4145
rect 8030 4075 8400 4085
rect 8430 4145 8800 4230
rect 8430 4085 8434 4145
rect 8486 4085 8744 4145
rect 8796 4085 8800 4145
rect 8430 4075 8800 4085
rect 8830 4145 9200 4230
rect 8830 4085 8834 4145
rect 8886 4085 9144 4145
rect 9196 4085 9200 4145
rect 8830 4075 9200 4085
rect 9230 4145 9600 4230
rect 9230 4085 9234 4145
rect 9286 4085 9544 4145
rect 9596 4085 9600 4145
rect 9230 4075 9600 4085
rect 9630 4145 10000 4230
rect 9630 4085 9634 4145
rect 9686 4085 9944 4145
rect 9996 4085 10000 4145
rect 9630 4075 10000 4085
rect 10030 4145 10400 4230
rect 10030 4085 10034 4145
rect 10086 4085 10344 4145
rect 10396 4085 10400 4145
rect 10030 4075 10400 4085
rect 10430 4145 10800 4230
rect 10430 4085 10434 4145
rect 10486 4085 10744 4145
rect 10796 4085 10800 4145
rect 10430 4075 10800 4085
rect 10830 4145 11200 4230
rect 10830 4085 10834 4145
rect 10886 4085 11144 4145
rect 11196 4085 11200 4145
rect 10830 4075 11200 4085
rect 11230 4145 11600 4230
rect 11230 4085 11234 4145
rect 11286 4085 11544 4145
rect 11596 4085 11600 4145
rect 11230 4075 11600 4085
rect 11630 4145 12000 4230
rect 11630 4085 11634 4145
rect 11686 4085 11944 4145
rect 11996 4085 12000 4145
rect 11630 4075 12000 4085
rect 12030 4145 12400 4230
rect 12030 4085 12034 4145
rect 12086 4085 12344 4145
rect 12396 4085 12400 4145
rect 12030 4075 12400 4085
rect 12430 4145 12800 4230
rect 12430 4085 12434 4145
rect 12486 4085 12744 4145
rect 12796 4085 12800 4145
rect 12430 4075 12800 4085
rect 12830 4145 13200 4230
rect 12830 4085 12834 4145
rect 12886 4085 13144 4145
rect 13196 4085 13200 4145
rect 12830 4075 13200 4085
rect -330 4045 -324 4075
rect 30 4045 70 4075
rect 430 4045 470 4075
rect 830 4045 870 4075
rect 1230 4045 1270 4075
rect 1630 4045 1670 4075
rect 2030 4045 2070 4075
rect 2430 4045 2470 4075
rect 2830 4045 2870 4075
rect -330 4035 0 4045
rect -314 3975 -56 4035
rect -4 3975 0 4035
rect -330 3775 0 3975
rect -314 3715 -56 3775
rect -4 3715 0 3775
rect -330 3705 0 3715
rect 30 4035 400 4045
rect 30 3975 34 4035
rect 86 3975 344 4035
rect 396 3975 400 4035
rect 30 3900 400 3975
rect 430 4035 800 4045
rect 430 3975 434 4035
rect 486 3975 744 4035
rect 796 3975 800 4035
rect 430 3900 800 3975
rect 830 4035 1200 4045
rect 830 3975 834 4035
rect 886 3975 1144 4035
rect 1196 3975 1200 4035
rect 830 3900 1200 3975
rect 1230 4035 1600 4045
rect 1230 3975 1234 4035
rect 1286 3975 1544 4035
rect 1596 3975 1600 4035
rect 1230 3900 1600 3975
rect 1630 4035 2000 4045
rect 1630 3975 1634 4035
rect 1686 3975 1944 4035
rect 1996 3975 2000 4035
rect 1630 3900 2000 3975
rect 2030 4035 2400 4045
rect 2030 3975 2034 4035
rect 2086 3975 2344 4035
rect 2396 3975 2400 4035
rect 2030 3900 2400 3975
rect 2430 4035 2800 4045
rect 2430 3975 2434 4035
rect 2486 3975 2744 4035
rect 2796 3975 2800 4035
rect 2430 3900 2800 3975
rect 2830 4035 3200 4045
rect 2830 3975 2834 4035
rect 2886 3975 3144 4035
rect 3196 3975 3200 4035
rect 2830 3900 3200 3975
rect 3230 4035 3600 4045
rect 3230 3975 3234 4035
rect 3286 3975 3544 4035
rect 3596 3975 3600 4035
rect 3230 3900 3600 3975
rect 3630 4035 4000 4045
rect 3630 3975 3634 4035
rect 3686 3975 3944 4035
rect 3996 3975 4000 4035
rect 3630 3900 4000 3975
rect 4030 4035 4400 4045
rect 4030 3975 4034 4035
rect 4086 3975 4344 4035
rect 4396 3975 4400 4035
rect 4030 3900 4400 3975
rect 4430 4035 4800 4045
rect 4430 3975 4434 4035
rect 4486 3975 4744 4035
rect 4796 3975 4800 4035
rect 4430 3900 4800 3975
rect 4830 4035 5200 4045
rect 4830 3975 4834 4035
rect 4886 3975 5144 4035
rect 5196 3975 5200 4035
rect 4830 3900 5200 3975
rect 5230 4035 5600 4045
rect 5230 3975 5234 4035
rect 5286 3975 5544 4035
rect 5596 3975 5600 4035
rect 5230 3900 5600 3975
rect 5630 4035 6000 4045
rect 5630 3975 5634 4035
rect 5686 3975 5944 4035
rect 5996 3975 6000 4035
rect 5630 3900 6000 3975
rect 6030 4035 6400 4045
rect 6030 3975 6034 4035
rect 6086 3975 6344 4035
rect 6396 3975 6400 4035
rect 6030 3900 6400 3975
rect 6430 4035 6800 4045
rect 6430 3975 6434 4035
rect 6486 3975 6744 4035
rect 6796 3975 6800 4035
rect 6430 3900 6800 3975
rect 6830 4035 7200 4045
rect 6830 3975 6834 4035
rect 6886 3975 7144 4035
rect 7196 3975 7200 4035
rect 6830 3900 7200 3975
rect 7230 4035 7600 4045
rect 7230 3975 7234 4035
rect 7286 3975 7544 4035
rect 7596 3975 7600 4035
rect 7230 3900 7600 3975
rect 7630 4035 8000 4045
rect 7630 3975 7634 4035
rect 7686 3975 7944 4035
rect 7996 3975 8000 4035
rect 7630 3900 8000 3975
rect 8030 4035 8400 4045
rect 8030 3975 8034 4035
rect 8086 3975 8344 4035
rect 8396 3975 8400 4035
rect 8030 3900 8400 3975
rect 8430 4035 8800 4045
rect 8430 3975 8434 4035
rect 8486 3975 8744 4035
rect 8796 3975 8800 4035
rect 8430 3900 8800 3975
rect 8830 4035 9200 4045
rect 8830 3975 8834 4035
rect 8886 3975 9144 4035
rect 9196 3975 9200 4035
rect 8830 3900 9200 3975
rect 9230 4035 9600 4045
rect 9230 3975 9234 4035
rect 9286 3975 9544 4035
rect 9596 3975 9600 4035
rect 9230 3900 9600 3975
rect 9630 4035 10000 4045
rect 9630 3975 9634 4035
rect 9686 3975 9944 4035
rect 9996 3975 10000 4035
rect 9630 3900 10000 3975
rect 10030 4035 10400 4045
rect 10030 3975 10034 4035
rect 10086 3975 10344 4035
rect 10396 3975 10400 4035
rect 10030 3900 10400 3975
rect 10430 4035 10800 4045
rect 10430 3975 10434 4035
rect 10486 3975 10744 4035
rect 10796 3975 10800 4035
rect 10430 3900 10800 3975
rect 10830 4035 11200 4045
rect 10830 3975 10834 4035
rect 10886 3975 11144 4035
rect 11196 3975 11200 4035
rect 10830 3900 11200 3975
rect 11230 4035 11600 4045
rect 11230 3975 11234 4035
rect 11286 3975 11544 4035
rect 11596 3975 11600 4035
rect 11230 3900 11600 3975
rect 11630 4035 12000 4045
rect 11630 3975 11634 4035
rect 11686 3975 11944 4035
rect 11996 3975 12000 4035
rect 11630 3900 12000 3975
rect 12030 4035 12400 4045
rect 12030 3975 12034 4035
rect 12086 3975 12344 4035
rect 12396 3975 12400 4035
rect 12030 3900 12400 3975
rect 12430 4035 12800 4045
rect 12430 3975 12434 4035
rect 12486 3975 12744 4035
rect 12796 3975 12800 4035
rect 12430 3900 12800 3975
rect 12830 4035 13200 4045
rect 12830 3975 12834 4035
rect 12886 3975 13144 4035
rect 13196 3975 13200 4035
rect 12830 3900 13200 3975
rect 30 3860 13390 3900
rect 30 3775 400 3860
rect 30 3715 34 3775
rect 86 3715 344 3775
rect 396 3715 400 3775
rect 30 3705 400 3715
rect 430 3775 800 3860
rect 430 3715 434 3775
rect 486 3715 744 3775
rect 796 3715 800 3775
rect 430 3705 800 3715
rect 830 3775 1200 3860
rect 830 3715 834 3775
rect 886 3715 1144 3775
rect 1196 3715 1200 3775
rect 830 3705 1200 3715
rect 1230 3775 1600 3860
rect 1230 3715 1234 3775
rect 1286 3715 1544 3775
rect 1596 3715 1600 3775
rect 1230 3705 1600 3715
rect 1630 3775 2000 3860
rect 1630 3715 1634 3775
rect 1686 3715 1944 3775
rect 1996 3715 2000 3775
rect 1630 3705 2000 3715
rect 2030 3775 2400 3860
rect 2030 3715 2034 3775
rect 2086 3715 2344 3775
rect 2396 3715 2400 3775
rect 2030 3705 2400 3715
rect 2430 3775 2800 3860
rect 2430 3715 2434 3775
rect 2486 3715 2744 3775
rect 2796 3715 2800 3775
rect 2430 3705 2800 3715
rect 2830 3775 3200 3860
rect 2830 3715 2834 3775
rect 2886 3715 3144 3775
rect 3196 3715 3200 3775
rect 2830 3705 3200 3715
rect 3230 3775 3600 3860
rect 3230 3715 3234 3775
rect 3286 3715 3544 3775
rect 3596 3715 3600 3775
rect 3230 3705 3600 3715
rect 3630 3775 4000 3860
rect 3630 3715 3634 3775
rect 3686 3715 3944 3775
rect 3996 3715 4000 3775
rect 3630 3705 4000 3715
rect 4030 3775 4400 3860
rect 4030 3715 4034 3775
rect 4086 3715 4344 3775
rect 4396 3715 4400 3775
rect 4030 3705 4400 3715
rect 4430 3775 4800 3860
rect 4430 3715 4434 3775
rect 4486 3715 4744 3775
rect 4796 3715 4800 3775
rect 4430 3705 4800 3715
rect 4830 3775 5200 3860
rect 4830 3715 4834 3775
rect 4886 3715 5144 3775
rect 5196 3715 5200 3775
rect 4830 3705 5200 3715
rect 5230 3775 5600 3860
rect 5230 3715 5234 3775
rect 5286 3715 5544 3775
rect 5596 3715 5600 3775
rect 5230 3705 5600 3715
rect 5630 3775 6000 3860
rect 5630 3715 5634 3775
rect 5686 3715 5944 3775
rect 5996 3715 6000 3775
rect 5630 3705 6000 3715
rect 6030 3775 6400 3860
rect 6030 3715 6034 3775
rect 6086 3715 6344 3775
rect 6396 3715 6400 3775
rect 6030 3705 6400 3715
rect 6430 3775 6800 3860
rect 6430 3715 6434 3775
rect 6486 3715 6744 3775
rect 6796 3715 6800 3775
rect 6430 3705 6800 3715
rect 6830 3775 7200 3860
rect 6830 3715 6834 3775
rect 6886 3715 7144 3775
rect 7196 3715 7200 3775
rect 6830 3705 7200 3715
rect 7230 3775 7600 3860
rect 7230 3715 7234 3775
rect 7286 3715 7544 3775
rect 7596 3715 7600 3775
rect 7230 3705 7600 3715
rect 7630 3775 8000 3860
rect 7630 3715 7634 3775
rect 7686 3715 7944 3775
rect 7996 3715 8000 3775
rect 7630 3705 8000 3715
rect 8030 3775 8400 3860
rect 8030 3715 8034 3775
rect 8086 3715 8344 3775
rect 8396 3715 8400 3775
rect 8030 3705 8400 3715
rect 8430 3775 8800 3860
rect 8430 3715 8434 3775
rect 8486 3715 8744 3775
rect 8796 3715 8800 3775
rect 8430 3705 8800 3715
rect 8830 3775 9200 3860
rect 8830 3715 8834 3775
rect 8886 3715 9144 3775
rect 9196 3715 9200 3775
rect 8830 3705 9200 3715
rect 9230 3775 9600 3860
rect 9230 3715 9234 3775
rect 9286 3715 9544 3775
rect 9596 3715 9600 3775
rect 9230 3705 9600 3715
rect 9630 3775 10000 3860
rect 9630 3715 9634 3775
rect 9686 3715 9944 3775
rect 9996 3715 10000 3775
rect 9630 3705 10000 3715
rect 10030 3775 10400 3860
rect 10030 3715 10034 3775
rect 10086 3715 10344 3775
rect 10396 3715 10400 3775
rect 10030 3705 10400 3715
rect 10430 3775 10800 3860
rect 10430 3715 10434 3775
rect 10486 3715 10744 3775
rect 10796 3715 10800 3775
rect 10430 3705 10800 3715
rect 10830 3775 11200 3860
rect 10830 3715 10834 3775
rect 10886 3715 11144 3775
rect 11196 3715 11200 3775
rect 10830 3705 11200 3715
rect 11230 3775 11600 3860
rect 11230 3715 11234 3775
rect 11286 3715 11544 3775
rect 11596 3715 11600 3775
rect 11230 3705 11600 3715
rect 11630 3775 12000 3860
rect 11630 3715 11634 3775
rect 11686 3715 11944 3775
rect 11996 3715 12000 3775
rect 11630 3705 12000 3715
rect 12030 3775 12400 3860
rect 12030 3715 12034 3775
rect 12086 3715 12344 3775
rect 12396 3715 12400 3775
rect 12030 3705 12400 3715
rect 12430 3775 12800 3860
rect 12430 3715 12434 3775
rect 12486 3715 12744 3775
rect 12796 3715 12800 3775
rect 12430 3705 12800 3715
rect 12830 3775 13200 3860
rect 12830 3715 12834 3775
rect 12886 3715 13144 3775
rect 13196 3715 13200 3775
rect 12830 3705 13200 3715
rect -330 3675 -324 3705
rect 30 3675 70 3705
rect 430 3675 470 3705
rect 830 3675 870 3705
rect 1230 3675 1270 3705
rect 1630 3675 1670 3705
rect 2030 3675 2070 3705
rect 2430 3675 2470 3705
rect 2830 3675 2870 3705
rect 3230 3675 3270 3705
rect 3630 3675 3670 3705
rect 4030 3675 4070 3705
rect 4430 3675 4470 3705
rect 4830 3675 4870 3705
rect 5230 3675 5270 3705
rect 5630 3675 5670 3705
rect 6030 3675 6070 3705
rect 6430 3675 6470 3705
rect 6830 3675 6870 3705
rect 7230 3675 7270 3705
rect 7630 3675 7670 3705
rect 8030 3675 8070 3705
rect 8430 3675 8470 3705
rect 8830 3675 8870 3705
rect 9230 3675 9270 3705
rect 9630 3675 9670 3705
rect 10030 3675 10070 3705
rect 10430 3675 10470 3705
rect 10830 3675 10870 3705
rect 11230 3675 11270 3705
rect 11630 3675 11670 3705
rect 12030 3675 12070 3705
rect 12430 3675 12470 3705
rect -330 3665 0 3675
rect -314 3605 -56 3665
rect -4 3605 0 3665
rect -330 3405 0 3605
rect -314 3345 -56 3405
rect -4 3345 0 3405
rect -330 3335 0 3345
rect 30 3665 400 3675
rect 30 3605 34 3665
rect 86 3605 344 3665
rect 396 3605 400 3665
rect 30 3530 400 3605
rect 430 3665 800 3675
rect 430 3605 434 3665
rect 486 3605 744 3665
rect 796 3605 800 3665
rect 430 3530 800 3605
rect 830 3665 1200 3675
rect 830 3605 834 3665
rect 886 3605 1144 3665
rect 1196 3605 1200 3665
rect 830 3530 1200 3605
rect 1230 3665 1600 3675
rect 1230 3605 1234 3665
rect 1286 3605 1544 3665
rect 1596 3605 1600 3665
rect 1230 3530 1600 3605
rect 1630 3665 2000 3675
rect 1630 3605 1634 3665
rect 1686 3605 1944 3665
rect 1996 3605 2000 3665
rect 1630 3530 2000 3605
rect 2030 3665 2400 3675
rect 2030 3605 2034 3665
rect 2086 3605 2344 3665
rect 2396 3605 2400 3665
rect 2030 3530 2400 3605
rect 2430 3665 2800 3675
rect 2430 3605 2434 3665
rect 2486 3605 2744 3665
rect 2796 3605 2800 3665
rect 2430 3530 2800 3605
rect 2830 3665 3200 3675
rect 2830 3605 2834 3665
rect 2886 3605 3144 3665
rect 3196 3605 3200 3665
rect 2830 3530 3200 3605
rect 3230 3665 3600 3675
rect 3230 3605 3234 3665
rect 3286 3605 3544 3665
rect 3596 3605 3600 3665
rect 3230 3530 3600 3605
rect 3630 3665 4000 3675
rect 3630 3605 3634 3665
rect 3686 3605 3944 3665
rect 3996 3605 4000 3665
rect 3630 3530 4000 3605
rect 4030 3665 4400 3675
rect 4030 3605 4034 3665
rect 4086 3605 4344 3665
rect 4396 3605 4400 3665
rect 4030 3530 4400 3605
rect 4430 3665 4800 3675
rect 4430 3605 4434 3665
rect 4486 3605 4744 3665
rect 4796 3605 4800 3665
rect 4430 3530 4800 3605
rect 4830 3665 5200 3675
rect 4830 3605 4834 3665
rect 4886 3605 5144 3665
rect 5196 3605 5200 3665
rect 4830 3530 5200 3605
rect 5230 3665 5600 3675
rect 5230 3605 5234 3665
rect 5286 3605 5544 3665
rect 5596 3605 5600 3665
rect 5230 3530 5600 3605
rect 5630 3665 6000 3675
rect 5630 3605 5634 3665
rect 5686 3605 5944 3665
rect 5996 3605 6000 3665
rect 5630 3530 6000 3605
rect 6030 3665 6400 3675
rect 6030 3605 6034 3665
rect 6086 3605 6344 3665
rect 6396 3605 6400 3665
rect 6030 3530 6400 3605
rect 6430 3665 6800 3675
rect 6430 3605 6434 3665
rect 6486 3605 6744 3665
rect 6796 3605 6800 3665
rect 6430 3530 6800 3605
rect 6830 3665 7200 3675
rect 6830 3605 6834 3665
rect 6886 3605 7144 3665
rect 7196 3605 7200 3665
rect 6830 3530 7200 3605
rect 7230 3665 7600 3675
rect 7230 3605 7234 3665
rect 7286 3605 7544 3665
rect 7596 3605 7600 3665
rect 7230 3530 7600 3605
rect 7630 3665 8000 3675
rect 7630 3605 7634 3665
rect 7686 3605 7944 3665
rect 7996 3605 8000 3665
rect 7630 3530 8000 3605
rect 8030 3665 8400 3675
rect 8030 3605 8034 3665
rect 8086 3605 8344 3665
rect 8396 3605 8400 3665
rect 8030 3530 8400 3605
rect 8430 3665 8800 3675
rect 8430 3605 8434 3665
rect 8486 3605 8744 3665
rect 8796 3605 8800 3665
rect 8430 3530 8800 3605
rect 8830 3665 9200 3675
rect 8830 3605 8834 3665
rect 8886 3605 9144 3665
rect 9196 3605 9200 3665
rect 8830 3530 9200 3605
rect 9230 3665 9600 3675
rect 9230 3605 9234 3665
rect 9286 3605 9544 3665
rect 9596 3605 9600 3665
rect 9230 3530 9600 3605
rect 9630 3665 10000 3675
rect 9630 3605 9634 3665
rect 9686 3605 9944 3665
rect 9996 3605 10000 3665
rect 9630 3530 10000 3605
rect 10030 3665 10400 3675
rect 10030 3605 10034 3665
rect 10086 3605 10344 3665
rect 10396 3605 10400 3665
rect 10030 3530 10400 3605
rect 10430 3665 10800 3675
rect 10430 3605 10434 3665
rect 10486 3605 10744 3665
rect 10796 3605 10800 3665
rect 10430 3530 10800 3605
rect 10830 3665 11200 3675
rect 10830 3605 10834 3665
rect 10886 3605 11144 3665
rect 11196 3605 11200 3665
rect 10830 3530 11200 3605
rect 11230 3665 11600 3675
rect 11230 3605 11234 3665
rect 11286 3605 11544 3665
rect 11596 3605 11600 3665
rect 11230 3530 11600 3605
rect 11630 3665 12000 3675
rect 11630 3605 11634 3665
rect 11686 3605 11944 3665
rect 11996 3605 12000 3665
rect 11630 3530 12000 3605
rect 12030 3665 12400 3675
rect 12030 3605 12034 3665
rect 12086 3605 12344 3665
rect 12396 3605 12400 3665
rect 12030 3530 12400 3605
rect 12430 3665 12800 3675
rect 12430 3605 12434 3665
rect 12486 3605 12744 3665
rect 12796 3605 12800 3665
rect 12430 3530 12800 3605
rect 12830 3665 13200 3675
rect 12830 3605 12834 3665
rect 12886 3605 13144 3665
rect 13196 3605 13200 3665
rect 12830 3530 13200 3605
rect 30 3490 13200 3530
rect 30 3405 400 3490
rect 30 3345 34 3405
rect 86 3345 344 3405
rect 396 3345 400 3405
rect 30 3335 400 3345
rect 430 3405 800 3490
rect 430 3345 434 3405
rect 486 3345 744 3405
rect 796 3345 800 3405
rect 430 3335 800 3345
rect 830 3405 1200 3490
rect 830 3345 834 3405
rect 886 3345 1144 3405
rect 1196 3345 1200 3405
rect 830 3335 1200 3345
rect 1230 3405 1600 3490
rect 1230 3345 1234 3405
rect 1286 3345 1544 3405
rect 1596 3345 1600 3405
rect 1230 3335 1600 3345
rect 1630 3405 2000 3490
rect 1630 3345 1634 3405
rect 1686 3345 1944 3405
rect 1996 3345 2000 3405
rect 1630 3335 2000 3345
rect 2030 3405 2400 3490
rect 2030 3345 2034 3405
rect 2086 3345 2344 3405
rect 2396 3345 2400 3405
rect 2030 3335 2400 3345
rect 2430 3405 2800 3490
rect 2430 3345 2434 3405
rect 2486 3345 2744 3405
rect 2796 3345 2800 3405
rect 2430 3335 2800 3345
rect 2830 3405 3200 3490
rect 2830 3345 2834 3405
rect 2886 3345 3144 3405
rect 3196 3345 3200 3405
rect 2830 3335 3200 3345
rect 3230 3405 3600 3490
rect 3230 3345 3234 3405
rect 3286 3345 3544 3405
rect 3596 3345 3600 3405
rect 3230 3335 3600 3345
rect 3630 3405 4000 3490
rect 3630 3345 3634 3405
rect 3686 3345 3944 3405
rect 3996 3345 4000 3405
rect 3630 3335 4000 3345
rect 4030 3405 4400 3490
rect 4030 3345 4034 3405
rect 4086 3345 4344 3405
rect 4396 3345 4400 3405
rect 4030 3335 4400 3345
rect 4430 3405 4800 3490
rect 4430 3345 4434 3405
rect 4486 3345 4744 3405
rect 4796 3345 4800 3405
rect 4430 3335 4800 3345
rect 4830 3405 5200 3490
rect 4830 3345 4834 3405
rect 4886 3345 5144 3405
rect 5196 3345 5200 3405
rect 4830 3335 5200 3345
rect 5230 3405 5600 3490
rect 5230 3345 5234 3405
rect 5286 3345 5544 3405
rect 5596 3345 5600 3405
rect 5230 3335 5600 3345
rect 5630 3405 6000 3490
rect 5630 3345 5634 3405
rect 5686 3345 5944 3405
rect 5996 3345 6000 3405
rect 5630 3335 6000 3345
rect 6030 3405 6400 3490
rect 6030 3345 6034 3405
rect 6086 3345 6344 3405
rect 6396 3345 6400 3405
rect 6030 3335 6400 3345
rect 6430 3405 6800 3490
rect 6430 3345 6434 3405
rect 6486 3345 6744 3405
rect 6796 3345 6800 3405
rect 6430 3335 6800 3345
rect 6830 3405 7200 3490
rect 6830 3345 6834 3405
rect 6886 3345 7144 3405
rect 7196 3345 7200 3405
rect 6830 3335 7200 3345
rect 7230 3405 7600 3490
rect 7230 3345 7234 3405
rect 7286 3345 7544 3405
rect 7596 3345 7600 3405
rect 7230 3335 7600 3345
rect 7630 3405 8000 3490
rect 7630 3345 7634 3405
rect 7686 3345 7944 3405
rect 7996 3345 8000 3405
rect 7630 3335 8000 3345
rect 8030 3405 8400 3490
rect 8030 3345 8034 3405
rect 8086 3345 8344 3405
rect 8396 3345 8400 3405
rect 8030 3335 8400 3345
rect 8430 3405 8800 3490
rect 8430 3345 8434 3405
rect 8486 3345 8744 3405
rect 8796 3345 8800 3405
rect 8430 3335 8800 3345
rect 8830 3405 9200 3490
rect 8830 3345 8834 3405
rect 8886 3345 9144 3405
rect 9196 3345 9200 3405
rect 8830 3335 9200 3345
rect 9230 3405 9600 3490
rect 9230 3345 9234 3405
rect 9286 3345 9544 3405
rect 9596 3345 9600 3405
rect 9230 3335 9600 3345
rect 9630 3405 10000 3490
rect 9630 3345 9634 3405
rect 9686 3345 9944 3405
rect 9996 3345 10000 3405
rect 9630 3335 10000 3345
rect 10030 3405 10400 3490
rect 10030 3345 10034 3405
rect 10086 3345 10344 3405
rect 10396 3345 10400 3405
rect 10030 3335 10400 3345
rect 10430 3405 10800 3490
rect 10430 3345 10434 3405
rect 10486 3345 10744 3405
rect 10796 3345 10800 3405
rect 10430 3335 10800 3345
rect 10830 3405 11200 3490
rect 10830 3345 10834 3405
rect 10886 3345 11144 3405
rect 11196 3345 11200 3405
rect 10830 3335 11200 3345
rect 11230 3405 11600 3490
rect 11230 3345 11234 3405
rect 11286 3345 11544 3405
rect 11596 3345 11600 3405
rect 11230 3335 11600 3345
rect 11630 3405 12000 3490
rect 11630 3345 11634 3405
rect 11686 3345 11944 3405
rect 11996 3345 12000 3405
rect 11630 3335 12000 3345
rect 12030 3405 12400 3490
rect 12030 3345 12034 3405
rect 12086 3345 12344 3405
rect 12396 3345 12400 3405
rect 12030 3335 12400 3345
rect 12430 3405 12800 3490
rect 12430 3345 12434 3405
rect 12486 3345 12744 3405
rect 12796 3345 12800 3405
rect 12430 3335 12800 3345
rect 12830 3405 13200 3490
rect 12830 3345 12834 3405
rect 12886 3345 13144 3405
rect 13196 3345 13200 3405
rect 12830 3335 13200 3345
rect -330 3305 -324 3335
rect 30 3305 70 3335
rect 430 3305 470 3335
rect 830 3305 870 3335
rect 1230 3305 1270 3335
rect 1630 3305 1670 3335
rect 2030 3305 2070 3335
rect 2430 3305 2470 3335
rect 2830 3305 2870 3335
rect 3230 3305 3270 3335
rect 3630 3305 3670 3335
rect 4030 3305 4070 3335
rect 4430 3305 4470 3335
rect 4830 3305 4870 3335
rect 5230 3305 5270 3335
rect 5630 3305 5670 3335
rect 6030 3305 6070 3335
rect 6430 3305 6470 3335
rect 6830 3305 6870 3335
rect 7230 3305 7270 3335
rect 7630 3305 7670 3335
rect 8030 3305 8070 3335
rect 8430 3305 8470 3335
rect 8830 3305 8870 3335
rect 9230 3305 9270 3335
rect 9630 3305 9670 3335
rect 10030 3305 10070 3335
rect 10430 3305 10470 3335
rect 10830 3305 10870 3335
rect 11230 3305 11270 3335
rect 11630 3305 11670 3335
rect 12030 3305 12070 3335
rect 12430 3305 12470 3335
rect -330 3295 0 3305
rect -314 3235 -56 3295
rect -4 3235 0 3295
rect -330 3035 0 3235
rect -314 2975 -56 3035
rect -4 2975 0 3035
rect -330 2965 0 2975
rect 30 3295 400 3305
rect 30 3235 34 3295
rect 86 3235 344 3295
rect 396 3235 400 3295
rect 30 3160 400 3235
rect 430 3295 800 3305
rect 430 3235 434 3295
rect 486 3235 744 3295
rect 796 3235 800 3295
rect 430 3160 800 3235
rect 830 3295 1200 3305
rect 830 3235 834 3295
rect 886 3235 1144 3295
rect 1196 3235 1200 3295
rect 830 3160 1200 3235
rect 1230 3295 1600 3305
rect 1230 3235 1234 3295
rect 1286 3235 1544 3295
rect 1596 3235 1600 3295
rect 1230 3160 1600 3235
rect 1630 3295 2000 3305
rect 1630 3235 1634 3295
rect 1686 3235 1944 3295
rect 1996 3235 2000 3295
rect 1630 3160 2000 3235
rect 2030 3295 2400 3305
rect 2030 3235 2034 3295
rect 2086 3235 2344 3295
rect 2396 3235 2400 3295
rect 2030 3160 2400 3235
rect 2430 3295 2800 3305
rect 2430 3235 2434 3295
rect 2486 3235 2744 3295
rect 2796 3235 2800 3295
rect 2430 3160 2800 3235
rect 2830 3295 3200 3305
rect 2830 3235 2834 3295
rect 2886 3235 3144 3295
rect 3196 3235 3200 3295
rect 2830 3160 3200 3235
rect 3230 3295 3600 3305
rect 3230 3235 3234 3295
rect 3286 3235 3544 3295
rect 3596 3235 3600 3295
rect 3230 3160 3600 3235
rect 3630 3295 4000 3305
rect 3630 3235 3634 3295
rect 3686 3235 3944 3295
rect 3996 3235 4000 3295
rect 3630 3160 4000 3235
rect 4030 3295 4400 3305
rect 4030 3235 4034 3295
rect 4086 3235 4344 3295
rect 4396 3235 4400 3295
rect 4030 3160 4400 3235
rect 4430 3295 4800 3305
rect 4430 3235 4434 3295
rect 4486 3235 4744 3295
rect 4796 3235 4800 3295
rect 4430 3160 4800 3235
rect 4830 3295 5200 3305
rect 4830 3235 4834 3295
rect 4886 3235 5144 3295
rect 5196 3235 5200 3295
rect 4830 3160 5200 3235
rect 5230 3295 5600 3305
rect 5230 3235 5234 3295
rect 5286 3235 5544 3295
rect 5596 3235 5600 3295
rect 5230 3160 5600 3235
rect 5630 3295 6000 3305
rect 5630 3235 5634 3295
rect 5686 3235 5944 3295
rect 5996 3235 6000 3295
rect 5630 3160 6000 3235
rect 6030 3295 6400 3305
rect 6030 3235 6034 3295
rect 6086 3235 6344 3295
rect 6396 3235 6400 3295
rect 6030 3160 6400 3235
rect 6430 3295 6800 3305
rect 6430 3235 6434 3295
rect 6486 3235 6744 3295
rect 6796 3235 6800 3295
rect 6430 3160 6800 3235
rect 6830 3295 7200 3305
rect 6830 3235 6834 3295
rect 6886 3235 7144 3295
rect 7196 3235 7200 3295
rect 6830 3160 7200 3235
rect 7230 3295 7600 3305
rect 7230 3235 7234 3295
rect 7286 3235 7544 3295
rect 7596 3235 7600 3295
rect 7230 3160 7600 3235
rect 7630 3295 8000 3305
rect 7630 3235 7634 3295
rect 7686 3235 7944 3295
rect 7996 3235 8000 3295
rect 7630 3160 8000 3235
rect 8030 3295 8400 3305
rect 8030 3235 8034 3295
rect 8086 3235 8344 3295
rect 8396 3235 8400 3295
rect 8030 3160 8400 3235
rect 8430 3295 8800 3305
rect 8430 3235 8434 3295
rect 8486 3235 8744 3295
rect 8796 3235 8800 3295
rect 8430 3160 8800 3235
rect 8830 3295 9200 3305
rect 8830 3235 8834 3295
rect 8886 3235 9144 3295
rect 9196 3235 9200 3295
rect 8830 3160 9200 3235
rect 9230 3295 9600 3305
rect 9230 3235 9234 3295
rect 9286 3235 9544 3295
rect 9596 3235 9600 3295
rect 9230 3160 9600 3235
rect 9630 3295 10000 3305
rect 9630 3235 9634 3295
rect 9686 3235 9944 3295
rect 9996 3235 10000 3295
rect 9630 3160 10000 3235
rect 10030 3295 10400 3305
rect 10030 3235 10034 3295
rect 10086 3235 10344 3295
rect 10396 3235 10400 3295
rect 10030 3160 10400 3235
rect 10430 3295 10800 3305
rect 10430 3235 10434 3295
rect 10486 3235 10744 3295
rect 10796 3235 10800 3295
rect 10430 3160 10800 3235
rect 10830 3295 11200 3305
rect 10830 3235 10834 3295
rect 10886 3235 11144 3295
rect 11196 3235 11200 3295
rect 10830 3160 11200 3235
rect 11230 3295 11600 3305
rect 11230 3235 11234 3295
rect 11286 3235 11544 3295
rect 11596 3235 11600 3295
rect 11230 3160 11600 3235
rect 11630 3295 12000 3305
rect 11630 3235 11634 3295
rect 11686 3235 11944 3295
rect 11996 3235 12000 3295
rect 11630 3160 12000 3235
rect 12030 3295 12400 3305
rect 12030 3235 12034 3295
rect 12086 3235 12344 3295
rect 12396 3235 12400 3295
rect 12030 3160 12400 3235
rect 12430 3295 12800 3305
rect 12430 3235 12434 3295
rect 12486 3235 12744 3295
rect 12796 3235 12800 3295
rect 12430 3160 12800 3235
rect 12830 3295 13200 3305
rect 12830 3235 12834 3295
rect 12886 3235 13144 3295
rect 13196 3235 13200 3295
rect 12830 3160 13200 3235
rect 30 3120 13200 3160
rect 30 3035 400 3120
rect 30 2975 34 3035
rect 86 2975 344 3035
rect 396 2975 400 3035
rect 30 2965 400 2975
rect 430 3035 800 3120
rect 430 2975 434 3035
rect 486 2975 744 3035
rect 796 2975 800 3035
rect 430 2965 800 2975
rect 830 3035 1200 3120
rect 830 2975 834 3035
rect 886 2975 1144 3035
rect 1196 2975 1200 3035
rect 830 2965 1200 2975
rect 1230 3035 1600 3120
rect 1230 2975 1234 3035
rect 1286 2975 1544 3035
rect 1596 2975 1600 3035
rect 1230 2965 1600 2975
rect 1630 3035 2000 3120
rect 1630 2975 1634 3035
rect 1686 2975 1944 3035
rect 1996 2975 2000 3035
rect 1630 2965 2000 2975
rect 2030 3035 2400 3120
rect 2030 2975 2034 3035
rect 2086 2975 2344 3035
rect 2396 2975 2400 3035
rect 2030 2965 2400 2975
rect 2430 3035 2800 3120
rect 2430 2975 2434 3035
rect 2486 2975 2744 3035
rect 2796 2975 2800 3035
rect 2430 2965 2800 2975
rect 2830 3035 3200 3120
rect 2830 2975 2834 3035
rect 2886 2975 3144 3035
rect 3196 2975 3200 3035
rect 2830 2965 3200 2975
rect 3230 3035 3600 3120
rect 3230 2975 3234 3035
rect 3286 2975 3544 3035
rect 3596 2975 3600 3035
rect 3230 2965 3600 2975
rect 3630 3035 4000 3120
rect 3630 2975 3634 3035
rect 3686 2975 3944 3035
rect 3996 2975 4000 3035
rect 3630 2965 4000 2975
rect 4030 3035 4400 3120
rect 4030 2975 4034 3035
rect 4086 2975 4344 3035
rect 4396 2975 4400 3035
rect 4030 2965 4400 2975
rect 4430 3035 4800 3120
rect 4430 2975 4434 3035
rect 4486 2975 4744 3035
rect 4796 2975 4800 3035
rect 4430 2965 4800 2975
rect 4830 3035 5200 3120
rect 4830 2975 4834 3035
rect 4886 2975 5144 3035
rect 5196 2975 5200 3035
rect 4830 2965 5200 2975
rect 5230 3035 5600 3120
rect 5230 2975 5234 3035
rect 5286 2975 5544 3035
rect 5596 2975 5600 3035
rect 5230 2965 5600 2975
rect 5630 3035 6000 3120
rect 5630 2975 5634 3035
rect 5686 2975 5944 3035
rect 5996 2975 6000 3035
rect 5630 2965 6000 2975
rect 6030 3035 6400 3120
rect 6030 2975 6034 3035
rect 6086 2975 6344 3035
rect 6396 2975 6400 3035
rect 6030 2965 6400 2975
rect 6430 3035 6800 3120
rect 6430 2975 6434 3035
rect 6486 2975 6744 3035
rect 6796 2975 6800 3035
rect 6430 2965 6800 2975
rect 6830 3035 7200 3120
rect 6830 2975 6834 3035
rect 6886 2975 7144 3035
rect 7196 2975 7200 3035
rect 6830 2965 7200 2975
rect 7230 3035 7600 3120
rect 7230 2975 7234 3035
rect 7286 2975 7544 3035
rect 7596 2975 7600 3035
rect 7230 2965 7600 2975
rect 7630 3035 8000 3120
rect 7630 2975 7634 3035
rect 7686 2975 7944 3035
rect 7996 2975 8000 3035
rect 7630 2965 8000 2975
rect 8030 3035 8400 3120
rect 8030 2975 8034 3035
rect 8086 2975 8344 3035
rect 8396 2975 8400 3035
rect 8030 2965 8400 2975
rect 8430 3035 8800 3120
rect 8430 2975 8434 3035
rect 8486 2975 8744 3035
rect 8796 2975 8800 3035
rect 8430 2965 8800 2975
rect 8830 3035 9200 3120
rect 8830 2975 8834 3035
rect 8886 2975 9144 3035
rect 9196 2975 9200 3035
rect 8830 2965 9200 2975
rect 9230 3035 9600 3120
rect 9230 2975 9234 3035
rect 9286 2975 9544 3035
rect 9596 2975 9600 3035
rect 9230 2965 9600 2975
rect 9630 3035 10000 3120
rect 9630 2975 9634 3035
rect 9686 2975 9944 3035
rect 9996 2975 10000 3035
rect 9630 2965 10000 2975
rect 10030 3035 10400 3120
rect 10030 2975 10034 3035
rect 10086 2975 10344 3035
rect 10396 2975 10400 3035
rect 10030 2965 10400 2975
rect 10430 3035 10800 3120
rect 10430 2975 10434 3035
rect 10486 2975 10744 3035
rect 10796 2975 10800 3035
rect 10430 2965 10800 2975
rect 10830 3035 11200 3120
rect 10830 2975 10834 3035
rect 10886 2975 11144 3035
rect 11196 2975 11200 3035
rect 10830 2965 11200 2975
rect 11230 3035 11600 3120
rect 11230 2975 11234 3035
rect 11286 2975 11544 3035
rect 11596 2975 11600 3035
rect 11230 2965 11600 2975
rect 11630 3035 12000 3120
rect 11630 2975 11634 3035
rect 11686 2975 11944 3035
rect 11996 2975 12000 3035
rect 11630 2965 12000 2975
rect 12030 3035 12400 3120
rect 12030 2975 12034 3035
rect 12086 2975 12344 3035
rect 12396 2975 12400 3035
rect 12030 2965 12400 2975
rect 12430 3035 12800 3120
rect 12430 2975 12434 3035
rect 12486 2975 12744 3035
rect 12796 2975 12800 3035
rect 12430 2965 12800 2975
rect 12830 3035 13200 3120
rect 12830 2975 12834 3035
rect 12886 2975 13144 3035
rect 13196 2975 13200 3035
rect 12830 2965 13200 2975
rect -330 2935 -324 2965
rect 30 2935 70 2965
rect 430 2935 470 2965
rect 830 2935 870 2965
rect 1230 2935 1270 2965
rect 1630 2935 1670 2965
rect 2030 2935 2070 2965
rect 2430 2935 2470 2965
rect 2830 2935 2870 2965
rect 3230 2935 3270 2965
rect 3630 2935 3670 2965
rect 4030 2935 4070 2965
rect 4430 2935 4470 2965
rect 4830 2935 4870 2965
rect 5230 2935 5270 2965
rect 5630 2935 5670 2965
rect 6030 2935 6070 2965
rect 6430 2935 6470 2965
rect 6830 2935 6870 2965
rect 7230 2935 7270 2965
rect 7630 2935 7670 2965
rect 8030 2935 8070 2965
rect 8430 2935 8470 2965
rect 8830 2935 8870 2965
rect 9230 2935 9270 2965
rect 9630 2935 9670 2965
rect 10030 2935 10070 2965
rect 10430 2935 10470 2965
rect 10830 2935 10870 2965
rect 11230 2935 11270 2965
rect 11630 2935 11670 2965
rect 12030 2935 12070 2965
rect 12430 2935 12470 2965
rect -330 2925 0 2935
rect -314 2865 -56 2925
rect -4 2865 0 2925
rect -330 2665 0 2865
rect -314 2605 -56 2665
rect -4 2605 0 2665
rect -330 2595 0 2605
rect 30 2925 400 2935
rect 30 2865 34 2925
rect 86 2865 344 2925
rect 396 2865 400 2925
rect 30 2790 400 2865
rect 430 2925 800 2935
rect 430 2865 434 2925
rect 486 2865 744 2925
rect 796 2865 800 2925
rect 430 2790 800 2865
rect 830 2925 1200 2935
rect 830 2865 834 2925
rect 886 2865 1144 2925
rect 1196 2865 1200 2925
rect 830 2790 1200 2865
rect 1230 2925 1600 2935
rect 1230 2865 1234 2925
rect 1286 2865 1544 2925
rect 1596 2865 1600 2925
rect 1230 2790 1600 2865
rect 1630 2925 2000 2935
rect 1630 2865 1634 2925
rect 1686 2865 1944 2925
rect 1996 2865 2000 2925
rect 1630 2790 2000 2865
rect 2030 2925 2400 2935
rect 2030 2865 2034 2925
rect 2086 2865 2344 2925
rect 2396 2865 2400 2925
rect 2030 2790 2400 2865
rect 2430 2925 2800 2935
rect 2430 2865 2434 2925
rect 2486 2865 2744 2925
rect 2796 2865 2800 2925
rect 2430 2790 2800 2865
rect 2830 2925 3200 2935
rect 2830 2865 2834 2925
rect 2886 2865 3144 2925
rect 3196 2865 3200 2925
rect 2830 2790 3200 2865
rect 3230 2925 3600 2935
rect 3230 2865 3234 2925
rect 3286 2865 3544 2925
rect 3596 2865 3600 2925
rect 3230 2790 3600 2865
rect 3630 2925 4000 2935
rect 3630 2865 3634 2925
rect 3686 2865 3944 2925
rect 3996 2865 4000 2925
rect 3630 2790 4000 2865
rect 4030 2925 4400 2935
rect 4030 2865 4034 2925
rect 4086 2865 4344 2925
rect 4396 2865 4400 2925
rect 4030 2790 4400 2865
rect 4430 2925 4800 2935
rect 4430 2865 4434 2925
rect 4486 2865 4744 2925
rect 4796 2865 4800 2925
rect 4430 2790 4800 2865
rect 4830 2925 5200 2935
rect 4830 2865 4834 2925
rect 4886 2865 5144 2925
rect 5196 2865 5200 2925
rect 4830 2790 5200 2865
rect 5230 2925 5600 2935
rect 5230 2865 5234 2925
rect 5286 2865 5544 2925
rect 5596 2865 5600 2925
rect 5230 2790 5600 2865
rect 5630 2925 6000 2935
rect 5630 2865 5634 2925
rect 5686 2865 5944 2925
rect 5996 2865 6000 2925
rect 5630 2790 6000 2865
rect 6030 2925 6400 2935
rect 6030 2865 6034 2925
rect 6086 2865 6344 2925
rect 6396 2865 6400 2925
rect 6030 2790 6400 2865
rect 6430 2925 6800 2935
rect 6430 2865 6434 2925
rect 6486 2865 6744 2925
rect 6796 2865 6800 2925
rect 6430 2790 6800 2865
rect 6830 2925 7200 2935
rect 6830 2865 6834 2925
rect 6886 2865 7144 2925
rect 7196 2865 7200 2925
rect 6830 2790 7200 2865
rect 7230 2925 7600 2935
rect 7230 2865 7234 2925
rect 7286 2865 7544 2925
rect 7596 2865 7600 2925
rect 7230 2790 7600 2865
rect 7630 2925 8000 2935
rect 7630 2865 7634 2925
rect 7686 2865 7944 2925
rect 7996 2865 8000 2925
rect 7630 2790 8000 2865
rect 8030 2925 8400 2935
rect 8030 2865 8034 2925
rect 8086 2865 8344 2925
rect 8396 2865 8400 2925
rect 8030 2790 8400 2865
rect 8430 2925 8800 2935
rect 8430 2865 8434 2925
rect 8486 2865 8744 2925
rect 8796 2865 8800 2925
rect 8430 2790 8800 2865
rect 8830 2925 9200 2935
rect 8830 2865 8834 2925
rect 8886 2865 9144 2925
rect 9196 2865 9200 2925
rect 8830 2790 9200 2865
rect 9230 2925 9600 2935
rect 9230 2865 9234 2925
rect 9286 2865 9544 2925
rect 9596 2865 9600 2925
rect 9230 2790 9600 2865
rect 9630 2925 10000 2935
rect 9630 2865 9634 2925
rect 9686 2865 9944 2925
rect 9996 2865 10000 2925
rect 9630 2790 10000 2865
rect 10030 2925 10400 2935
rect 10030 2865 10034 2925
rect 10086 2865 10344 2925
rect 10396 2865 10400 2925
rect 10030 2790 10400 2865
rect 10430 2925 10800 2935
rect 10430 2865 10434 2925
rect 10486 2865 10744 2925
rect 10796 2865 10800 2925
rect 10430 2790 10800 2865
rect 10830 2925 11200 2935
rect 10830 2865 10834 2925
rect 10886 2865 11144 2925
rect 11196 2865 11200 2925
rect 10830 2790 11200 2865
rect 11230 2925 11600 2935
rect 11230 2865 11234 2925
rect 11286 2865 11544 2925
rect 11596 2865 11600 2925
rect 11230 2790 11600 2865
rect 11630 2925 12000 2935
rect 11630 2865 11634 2925
rect 11686 2865 11944 2925
rect 11996 2865 12000 2925
rect 11630 2790 12000 2865
rect 12030 2925 12400 2935
rect 12030 2865 12034 2925
rect 12086 2865 12344 2925
rect 12396 2865 12400 2925
rect 12030 2790 12400 2865
rect 12430 2925 12800 2935
rect 12430 2865 12434 2925
rect 12486 2865 12744 2925
rect 12796 2865 12800 2925
rect 12430 2790 12800 2865
rect 12830 2925 13200 2935
rect 12830 2865 12834 2925
rect 12886 2865 13144 2925
rect 13196 2865 13200 2925
rect 12830 2790 13200 2865
rect 30 2750 13200 2790
rect 30 2665 400 2750
rect 30 2605 34 2665
rect 86 2605 344 2665
rect 396 2605 400 2665
rect 30 2595 400 2605
rect 430 2665 800 2750
rect 430 2605 434 2665
rect 486 2605 744 2665
rect 796 2605 800 2665
rect 430 2595 800 2605
rect 830 2665 1200 2750
rect 830 2605 834 2665
rect 886 2605 1144 2665
rect 1196 2605 1200 2665
rect 830 2595 1200 2605
rect 1230 2665 1600 2750
rect 1230 2605 1234 2665
rect 1286 2605 1544 2665
rect 1596 2605 1600 2665
rect 1230 2595 1600 2605
rect 1630 2665 2000 2750
rect 1630 2605 1634 2665
rect 1686 2605 1944 2665
rect 1996 2605 2000 2665
rect 1630 2595 2000 2605
rect 2030 2665 2400 2750
rect 2030 2605 2034 2665
rect 2086 2605 2344 2665
rect 2396 2605 2400 2665
rect 2030 2595 2400 2605
rect 2430 2665 2800 2750
rect 2430 2605 2434 2665
rect 2486 2605 2744 2665
rect 2796 2605 2800 2665
rect 2430 2595 2800 2605
rect 2830 2665 3200 2750
rect 2830 2605 2834 2665
rect 2886 2605 3144 2665
rect 3196 2605 3200 2665
rect 2830 2595 3200 2605
rect 3230 2665 3600 2750
rect 3230 2605 3234 2665
rect 3286 2605 3544 2665
rect 3596 2605 3600 2665
rect 3230 2595 3600 2605
rect 3630 2665 4000 2750
rect 3630 2605 3634 2665
rect 3686 2605 3944 2665
rect 3996 2605 4000 2665
rect 3630 2595 4000 2605
rect 4030 2665 4400 2750
rect 4030 2605 4034 2665
rect 4086 2605 4344 2665
rect 4396 2605 4400 2665
rect 4030 2595 4400 2605
rect 4430 2665 4800 2750
rect 4430 2605 4434 2665
rect 4486 2605 4744 2665
rect 4796 2605 4800 2665
rect 4430 2595 4800 2605
rect 4830 2665 5200 2750
rect 4830 2605 4834 2665
rect 4886 2605 5144 2665
rect 5196 2605 5200 2665
rect 4830 2595 5200 2605
rect 5230 2665 5600 2750
rect 5230 2605 5234 2665
rect 5286 2605 5544 2665
rect 5596 2605 5600 2665
rect 5230 2595 5600 2605
rect 5630 2665 6000 2750
rect 5630 2605 5634 2665
rect 5686 2605 5944 2665
rect 5996 2605 6000 2665
rect 5630 2595 6000 2605
rect 6030 2665 6400 2750
rect 6030 2605 6034 2665
rect 6086 2605 6344 2665
rect 6396 2605 6400 2665
rect 6030 2595 6400 2605
rect 6430 2665 6800 2750
rect 6430 2605 6434 2665
rect 6486 2605 6744 2665
rect 6796 2605 6800 2665
rect 6430 2595 6800 2605
rect 6830 2665 7200 2750
rect 6830 2605 6834 2665
rect 6886 2605 7144 2665
rect 7196 2605 7200 2665
rect 6830 2595 7200 2605
rect 7230 2665 7600 2750
rect 7230 2605 7234 2665
rect 7286 2605 7544 2665
rect 7596 2605 7600 2665
rect 7230 2595 7600 2605
rect 7630 2665 8000 2750
rect 7630 2605 7634 2665
rect 7686 2605 7944 2665
rect 7996 2605 8000 2665
rect 7630 2595 8000 2605
rect 8030 2665 8400 2750
rect 8030 2605 8034 2665
rect 8086 2605 8344 2665
rect 8396 2605 8400 2665
rect 8030 2595 8400 2605
rect 8430 2665 8800 2750
rect 8430 2605 8434 2665
rect 8486 2605 8744 2665
rect 8796 2605 8800 2665
rect 8430 2595 8800 2605
rect 8830 2665 9200 2750
rect 8830 2605 8834 2665
rect 8886 2605 9144 2665
rect 9196 2605 9200 2665
rect 8830 2595 9200 2605
rect 9230 2665 9600 2750
rect 9230 2605 9234 2665
rect 9286 2605 9544 2665
rect 9596 2605 9600 2665
rect 9230 2595 9600 2605
rect 9630 2665 10000 2750
rect 9630 2605 9634 2665
rect 9686 2605 9944 2665
rect 9996 2605 10000 2665
rect 9630 2595 10000 2605
rect 10030 2665 10400 2750
rect 10030 2605 10034 2665
rect 10086 2605 10344 2665
rect 10396 2605 10400 2665
rect 10030 2595 10400 2605
rect 10430 2665 10800 2750
rect 10430 2605 10434 2665
rect 10486 2605 10744 2665
rect 10796 2605 10800 2665
rect 10430 2595 10800 2605
rect 10830 2665 11200 2750
rect 10830 2605 10834 2665
rect 10886 2605 11144 2665
rect 11196 2605 11200 2665
rect 10830 2595 11200 2605
rect 11230 2665 11600 2750
rect 11230 2605 11234 2665
rect 11286 2605 11544 2665
rect 11596 2605 11600 2665
rect 11230 2595 11600 2605
rect 11630 2665 12000 2750
rect 11630 2605 11634 2665
rect 11686 2605 11944 2665
rect 11996 2605 12000 2665
rect 11630 2595 12000 2605
rect 12030 2665 12400 2750
rect 12030 2605 12034 2665
rect 12086 2605 12344 2665
rect 12396 2605 12400 2665
rect 12030 2595 12400 2605
rect 12430 2665 12800 2750
rect 12430 2605 12434 2665
rect 12486 2605 12744 2665
rect 12796 2605 12800 2665
rect 12430 2595 12800 2605
rect 12830 2665 13200 2750
rect 12830 2605 12834 2665
rect 12886 2605 13144 2665
rect 13196 2605 13200 2665
rect 12830 2595 13200 2605
rect -330 2565 -324 2595
rect 30 2565 70 2595
rect 430 2565 470 2595
rect 830 2565 870 2595
rect 1230 2565 1270 2595
rect 1630 2565 1670 2595
rect 2030 2565 2070 2595
rect 2430 2565 2470 2595
rect 2830 2565 2870 2595
rect 3230 2565 3270 2595
rect 3630 2565 3670 2595
rect 4030 2565 4070 2595
rect 4430 2565 4470 2595
rect 4830 2565 4870 2595
rect 5230 2565 5270 2595
rect 5630 2565 5670 2595
rect 6030 2565 6070 2595
rect 6430 2565 6470 2595
rect 6830 2565 6870 2595
rect 7230 2565 7270 2595
rect 7630 2565 7670 2595
rect 8030 2565 8070 2595
rect 8430 2565 8470 2595
rect 8830 2565 8870 2595
rect 9230 2565 9270 2595
rect 9630 2565 9670 2595
rect 10030 2565 10070 2595
rect 10430 2565 10470 2595
rect 10830 2565 10870 2595
rect 11230 2565 11270 2595
rect 11630 2565 11670 2595
rect 12030 2565 12070 2595
rect 12430 2565 12470 2595
rect -330 2555 0 2565
rect -314 2495 -56 2555
rect -4 2495 0 2555
rect -330 2295 0 2495
rect -314 2235 -56 2295
rect -4 2235 0 2295
rect -330 2225 0 2235
rect 30 2555 400 2565
rect 30 2495 34 2555
rect 86 2495 344 2555
rect 396 2495 400 2555
rect 30 2420 400 2495
rect 430 2555 800 2565
rect 430 2495 434 2555
rect 486 2495 744 2555
rect 796 2495 800 2555
rect 430 2420 800 2495
rect 830 2555 1200 2565
rect 830 2495 834 2555
rect 886 2495 1144 2555
rect 1196 2495 1200 2555
rect 830 2420 1200 2495
rect 1230 2555 1600 2565
rect 1230 2495 1234 2555
rect 1286 2495 1544 2555
rect 1596 2495 1600 2555
rect 1230 2420 1600 2495
rect 1630 2555 2000 2565
rect 1630 2495 1634 2555
rect 1686 2495 1944 2555
rect 1996 2495 2000 2555
rect 1630 2420 2000 2495
rect 2030 2555 2400 2565
rect 2030 2495 2034 2555
rect 2086 2495 2344 2555
rect 2396 2495 2400 2555
rect 2030 2420 2400 2495
rect 2430 2555 2800 2565
rect 2430 2495 2434 2555
rect 2486 2495 2744 2555
rect 2796 2495 2800 2555
rect 2430 2420 2800 2495
rect 2830 2555 3200 2565
rect 2830 2495 2834 2555
rect 2886 2495 3144 2555
rect 3196 2495 3200 2555
rect 2830 2420 3200 2495
rect 3230 2555 3600 2565
rect 3230 2495 3234 2555
rect 3286 2495 3544 2555
rect 3596 2495 3600 2555
rect 3230 2420 3600 2495
rect 3630 2555 4000 2565
rect 3630 2495 3634 2555
rect 3686 2495 3944 2555
rect 3996 2495 4000 2555
rect 3630 2420 4000 2495
rect 4030 2555 4400 2565
rect 4030 2495 4034 2555
rect 4086 2495 4344 2555
rect 4396 2495 4400 2555
rect 4030 2420 4400 2495
rect 4430 2555 4800 2565
rect 4430 2495 4434 2555
rect 4486 2495 4744 2555
rect 4796 2495 4800 2555
rect 4430 2420 4800 2495
rect 4830 2555 5200 2565
rect 4830 2495 4834 2555
rect 4886 2495 5144 2555
rect 5196 2495 5200 2555
rect 4830 2420 5200 2495
rect 5230 2555 5600 2565
rect 5230 2495 5234 2555
rect 5286 2495 5544 2555
rect 5596 2495 5600 2555
rect 5230 2420 5600 2495
rect 5630 2555 6000 2565
rect 5630 2495 5634 2555
rect 5686 2495 5944 2555
rect 5996 2495 6000 2555
rect 5630 2420 6000 2495
rect 6030 2555 6400 2565
rect 6030 2495 6034 2555
rect 6086 2495 6344 2555
rect 6396 2495 6400 2555
rect 6030 2420 6400 2495
rect 6430 2555 6800 2565
rect 6430 2495 6434 2555
rect 6486 2495 6744 2555
rect 6796 2495 6800 2555
rect 6430 2420 6800 2495
rect 6830 2555 7200 2565
rect 6830 2495 6834 2555
rect 6886 2495 7144 2555
rect 7196 2495 7200 2555
rect 6830 2420 7200 2495
rect 7230 2555 7600 2565
rect 7230 2495 7234 2555
rect 7286 2495 7544 2555
rect 7596 2495 7600 2555
rect 7230 2420 7600 2495
rect 7630 2555 8000 2565
rect 7630 2495 7634 2555
rect 7686 2495 7944 2555
rect 7996 2495 8000 2555
rect 7630 2420 8000 2495
rect 8030 2555 8400 2565
rect 8030 2495 8034 2555
rect 8086 2495 8344 2555
rect 8396 2495 8400 2555
rect 8030 2420 8400 2495
rect 8430 2555 8800 2565
rect 8430 2495 8434 2555
rect 8486 2495 8744 2555
rect 8796 2495 8800 2555
rect 8430 2420 8800 2495
rect 8830 2555 9200 2565
rect 8830 2495 8834 2555
rect 8886 2495 9144 2555
rect 9196 2495 9200 2555
rect 8830 2420 9200 2495
rect 9230 2555 9600 2565
rect 9230 2495 9234 2555
rect 9286 2495 9544 2555
rect 9596 2495 9600 2555
rect 9230 2420 9600 2495
rect 9630 2555 10000 2565
rect 9630 2495 9634 2555
rect 9686 2495 9944 2555
rect 9996 2495 10000 2555
rect 9630 2420 10000 2495
rect 10030 2555 10400 2565
rect 10030 2495 10034 2555
rect 10086 2495 10344 2555
rect 10396 2495 10400 2555
rect 10030 2420 10400 2495
rect 10430 2555 10800 2565
rect 10430 2495 10434 2555
rect 10486 2495 10744 2555
rect 10796 2495 10800 2555
rect 10430 2420 10800 2495
rect 10830 2555 11200 2565
rect 10830 2495 10834 2555
rect 10886 2495 11144 2555
rect 11196 2495 11200 2555
rect 10830 2420 11200 2495
rect 11230 2555 11600 2565
rect 11230 2495 11234 2555
rect 11286 2495 11544 2555
rect 11596 2495 11600 2555
rect 11230 2420 11600 2495
rect 11630 2555 12000 2565
rect 11630 2495 11634 2555
rect 11686 2495 11944 2555
rect 11996 2495 12000 2555
rect 11630 2420 12000 2495
rect 12030 2555 12400 2565
rect 12030 2495 12034 2555
rect 12086 2495 12344 2555
rect 12396 2495 12400 2555
rect 12030 2420 12400 2495
rect 12430 2555 12800 2565
rect 12430 2495 12434 2555
rect 12486 2495 12744 2555
rect 12796 2495 12800 2555
rect 12430 2420 12800 2495
rect 12830 2555 13200 2565
rect 12830 2495 12834 2555
rect 12886 2495 13144 2555
rect 13196 2495 13200 2555
rect 12830 2420 13200 2495
rect 30 2380 13200 2420
rect 30 2295 400 2380
rect 30 2235 34 2295
rect 86 2235 344 2295
rect 396 2235 400 2295
rect 30 2225 400 2235
rect 430 2295 800 2380
rect 430 2235 434 2295
rect 486 2235 744 2295
rect 796 2235 800 2295
rect 430 2225 800 2235
rect 830 2295 1200 2380
rect 830 2235 834 2295
rect 886 2235 1144 2295
rect 1196 2235 1200 2295
rect 830 2225 1200 2235
rect 1230 2295 1600 2380
rect 1230 2235 1234 2295
rect 1286 2235 1544 2295
rect 1596 2235 1600 2295
rect 1230 2225 1600 2235
rect 1630 2295 2000 2380
rect 1630 2235 1634 2295
rect 1686 2235 1944 2295
rect 1996 2235 2000 2295
rect 1630 2225 2000 2235
rect 2030 2295 2400 2380
rect 2030 2235 2034 2295
rect 2086 2235 2344 2295
rect 2396 2235 2400 2295
rect 2030 2225 2400 2235
rect 2430 2295 2800 2380
rect 2430 2235 2434 2295
rect 2486 2235 2744 2295
rect 2796 2235 2800 2295
rect 2430 2225 2800 2235
rect 2830 2295 3200 2380
rect 2830 2235 2834 2295
rect 2886 2235 3144 2295
rect 3196 2235 3200 2295
rect 2830 2225 3200 2235
rect 3230 2295 3600 2380
rect 3230 2235 3234 2295
rect 3286 2235 3544 2295
rect 3596 2235 3600 2295
rect 3230 2225 3600 2235
rect 3630 2295 4000 2380
rect 3630 2235 3634 2295
rect 3686 2235 3944 2295
rect 3996 2235 4000 2295
rect 3630 2225 4000 2235
rect 4030 2295 4400 2380
rect 4030 2235 4034 2295
rect 4086 2235 4344 2295
rect 4396 2235 4400 2295
rect 4030 2225 4400 2235
rect 4430 2295 4800 2380
rect 4430 2235 4434 2295
rect 4486 2235 4744 2295
rect 4796 2235 4800 2295
rect 4430 2225 4800 2235
rect 4830 2295 5200 2380
rect 4830 2235 4834 2295
rect 4886 2235 5144 2295
rect 5196 2235 5200 2295
rect 4830 2225 5200 2235
rect 5230 2295 5600 2380
rect 5230 2235 5234 2295
rect 5286 2235 5544 2295
rect 5596 2235 5600 2295
rect 5230 2225 5600 2235
rect 5630 2295 6000 2380
rect 5630 2235 5634 2295
rect 5686 2235 5944 2295
rect 5996 2235 6000 2295
rect 5630 2225 6000 2235
rect 6030 2295 6400 2380
rect 6030 2235 6034 2295
rect 6086 2235 6344 2295
rect 6396 2235 6400 2295
rect 6030 2225 6400 2235
rect 6430 2295 6800 2380
rect 6430 2235 6434 2295
rect 6486 2235 6744 2295
rect 6796 2235 6800 2295
rect 6430 2225 6800 2235
rect 6830 2295 7200 2380
rect 6830 2235 6834 2295
rect 6886 2235 7144 2295
rect 7196 2235 7200 2295
rect 6830 2225 7200 2235
rect 7230 2295 7600 2380
rect 7230 2235 7234 2295
rect 7286 2235 7544 2295
rect 7596 2235 7600 2295
rect 7230 2225 7600 2235
rect 7630 2295 8000 2380
rect 7630 2235 7634 2295
rect 7686 2235 7944 2295
rect 7996 2235 8000 2295
rect 7630 2225 8000 2235
rect 8030 2295 8400 2380
rect 8030 2235 8034 2295
rect 8086 2235 8344 2295
rect 8396 2235 8400 2295
rect 8030 2225 8400 2235
rect 8430 2295 8800 2380
rect 8430 2235 8434 2295
rect 8486 2235 8744 2295
rect 8796 2235 8800 2295
rect 8430 2225 8800 2235
rect 8830 2295 9200 2380
rect 8830 2235 8834 2295
rect 8886 2235 9144 2295
rect 9196 2235 9200 2295
rect 8830 2225 9200 2235
rect 9230 2295 9600 2380
rect 9230 2235 9234 2295
rect 9286 2235 9544 2295
rect 9596 2235 9600 2295
rect 9230 2225 9600 2235
rect 9630 2295 10000 2380
rect 9630 2235 9634 2295
rect 9686 2235 9944 2295
rect 9996 2235 10000 2295
rect 9630 2225 10000 2235
rect 10030 2295 10400 2380
rect 10030 2235 10034 2295
rect 10086 2235 10344 2295
rect 10396 2235 10400 2295
rect 10030 2225 10400 2235
rect 10430 2295 10800 2380
rect 10430 2235 10434 2295
rect 10486 2235 10744 2295
rect 10796 2235 10800 2295
rect 10430 2225 10800 2235
rect 10830 2295 11200 2380
rect 10830 2235 10834 2295
rect 10886 2235 11144 2295
rect 11196 2235 11200 2295
rect 10830 2225 11200 2235
rect 11230 2295 11600 2380
rect 11230 2235 11234 2295
rect 11286 2235 11544 2295
rect 11596 2235 11600 2295
rect 11230 2225 11600 2235
rect 11630 2295 12000 2380
rect 11630 2235 11634 2295
rect 11686 2235 11944 2295
rect 11996 2235 12000 2295
rect 11630 2225 12000 2235
rect 12030 2295 12400 2380
rect 12030 2235 12034 2295
rect 12086 2235 12344 2295
rect 12396 2235 12400 2295
rect 12030 2225 12400 2235
rect 12430 2295 12800 2380
rect 12430 2235 12434 2295
rect 12486 2235 12744 2295
rect 12796 2235 12800 2295
rect 12430 2225 12800 2235
rect 12830 2295 13200 2380
rect 12830 2235 12834 2295
rect 12886 2235 13144 2295
rect 13196 2235 13200 2295
rect 12830 2225 13200 2235
rect -330 2195 -324 2225
rect 30 2195 70 2225
rect 430 2195 470 2225
rect 830 2195 870 2225
rect 1230 2195 1270 2225
rect 1630 2195 1670 2225
rect 2030 2195 2070 2225
rect 2430 2195 2470 2225
rect 2830 2195 2870 2225
rect 3230 2195 3270 2225
rect 3630 2195 3670 2225
rect 4030 2195 4070 2225
rect 4430 2195 4470 2225
rect 4830 2195 4870 2225
rect 5230 2195 5270 2225
rect 5630 2195 5670 2225
rect 6030 2195 6070 2225
rect 6430 2195 6470 2225
rect 6830 2195 6870 2225
rect 7230 2195 7270 2225
rect 7630 2195 7670 2225
rect 8030 2195 8070 2225
rect 8430 2195 8470 2225
rect 8830 2195 8870 2225
rect 9230 2195 9270 2225
rect 9630 2195 9670 2225
rect 10030 2195 10070 2225
rect 10430 2195 10470 2225
rect 10830 2195 10870 2225
rect 11230 2195 11270 2225
rect 11630 2195 11670 2225
rect 12030 2195 12070 2225
rect 12430 2195 12470 2225
rect -330 2185 0 2195
rect -314 2125 -56 2185
rect -4 2125 0 2185
rect -330 1925 0 2125
rect -314 1865 -56 1925
rect -4 1865 0 1925
rect -330 1855 0 1865
rect 30 2185 400 2195
rect 30 2125 34 2185
rect 86 2125 344 2185
rect 396 2125 400 2185
rect 30 2050 400 2125
rect 430 2185 800 2195
rect 430 2125 434 2185
rect 486 2125 744 2185
rect 796 2125 800 2185
rect 430 2050 800 2125
rect 830 2185 1200 2195
rect 830 2125 834 2185
rect 886 2125 1144 2185
rect 1196 2125 1200 2185
rect 830 2050 1200 2125
rect 1230 2185 1600 2195
rect 1230 2125 1234 2185
rect 1286 2125 1544 2185
rect 1596 2125 1600 2185
rect 1230 2050 1600 2125
rect 1630 2185 2000 2195
rect 1630 2125 1634 2185
rect 1686 2125 1944 2185
rect 1996 2125 2000 2185
rect 1630 2050 2000 2125
rect 2030 2185 2400 2195
rect 2030 2125 2034 2185
rect 2086 2125 2344 2185
rect 2396 2125 2400 2185
rect 2030 2050 2400 2125
rect 2430 2185 2800 2195
rect 2430 2125 2434 2185
rect 2486 2125 2744 2185
rect 2796 2125 2800 2185
rect 2430 2050 2800 2125
rect 2830 2185 3200 2195
rect 2830 2125 2834 2185
rect 2886 2125 3144 2185
rect 3196 2125 3200 2185
rect 2830 2050 3200 2125
rect 3230 2185 3600 2195
rect 3230 2125 3234 2185
rect 3286 2125 3544 2185
rect 3596 2125 3600 2185
rect 3230 2050 3600 2125
rect 3630 2185 4000 2195
rect 3630 2125 3634 2185
rect 3686 2125 3944 2185
rect 3996 2125 4000 2185
rect 3630 2050 4000 2125
rect 4030 2185 4400 2195
rect 4030 2125 4034 2185
rect 4086 2125 4344 2185
rect 4396 2125 4400 2185
rect 4030 2050 4400 2125
rect 4430 2185 4800 2195
rect 4430 2125 4434 2185
rect 4486 2125 4744 2185
rect 4796 2125 4800 2185
rect 4430 2050 4800 2125
rect 4830 2185 5200 2195
rect 4830 2125 4834 2185
rect 4886 2125 5144 2185
rect 5196 2125 5200 2185
rect 4830 2050 5200 2125
rect 5230 2185 5600 2195
rect 5230 2125 5234 2185
rect 5286 2125 5544 2185
rect 5596 2125 5600 2185
rect 5230 2050 5600 2125
rect 5630 2185 6000 2195
rect 5630 2125 5634 2185
rect 5686 2125 5944 2185
rect 5996 2125 6000 2185
rect 5630 2050 6000 2125
rect 6030 2185 6400 2195
rect 6030 2125 6034 2185
rect 6086 2125 6344 2185
rect 6396 2125 6400 2185
rect 6030 2050 6400 2125
rect 6430 2185 6800 2195
rect 6430 2125 6434 2185
rect 6486 2125 6744 2185
rect 6796 2125 6800 2185
rect 6430 2050 6800 2125
rect 6830 2185 7200 2195
rect 6830 2125 6834 2185
rect 6886 2125 7144 2185
rect 7196 2125 7200 2185
rect 6830 2050 7200 2125
rect 7230 2185 7600 2195
rect 7230 2125 7234 2185
rect 7286 2125 7544 2185
rect 7596 2125 7600 2185
rect 7230 2050 7600 2125
rect 7630 2185 8000 2195
rect 7630 2125 7634 2185
rect 7686 2125 7944 2185
rect 7996 2125 8000 2185
rect 7630 2050 8000 2125
rect 8030 2185 8400 2195
rect 8030 2125 8034 2185
rect 8086 2125 8344 2185
rect 8396 2125 8400 2185
rect 8030 2050 8400 2125
rect 8430 2185 8800 2195
rect 8430 2125 8434 2185
rect 8486 2125 8744 2185
rect 8796 2125 8800 2185
rect 8430 2050 8800 2125
rect 8830 2185 9200 2195
rect 8830 2125 8834 2185
rect 8886 2125 9144 2185
rect 9196 2125 9200 2185
rect 8830 2050 9200 2125
rect 9230 2185 9600 2195
rect 9230 2125 9234 2185
rect 9286 2125 9544 2185
rect 9596 2125 9600 2185
rect 9230 2050 9600 2125
rect 9630 2185 10000 2195
rect 9630 2125 9634 2185
rect 9686 2125 9944 2185
rect 9996 2125 10000 2185
rect 9630 2050 10000 2125
rect 10030 2185 10400 2195
rect 10030 2125 10034 2185
rect 10086 2125 10344 2185
rect 10396 2125 10400 2185
rect 10030 2050 10400 2125
rect 10430 2185 10800 2195
rect 10430 2125 10434 2185
rect 10486 2125 10744 2185
rect 10796 2125 10800 2185
rect 10430 2050 10800 2125
rect 10830 2185 11200 2195
rect 10830 2125 10834 2185
rect 10886 2125 11144 2185
rect 11196 2125 11200 2185
rect 10830 2050 11200 2125
rect 11230 2185 11600 2195
rect 11230 2125 11234 2185
rect 11286 2125 11544 2185
rect 11596 2125 11600 2185
rect 11230 2050 11600 2125
rect 11630 2185 12000 2195
rect 11630 2125 11634 2185
rect 11686 2125 11944 2185
rect 11996 2125 12000 2185
rect 11630 2050 12000 2125
rect 12030 2185 12400 2195
rect 12030 2125 12034 2185
rect 12086 2125 12344 2185
rect 12396 2125 12400 2185
rect 12030 2050 12400 2125
rect 12430 2185 12800 2195
rect 12430 2125 12434 2185
rect 12486 2125 12744 2185
rect 12796 2125 12800 2185
rect 12430 2050 12800 2125
rect 12830 2185 13200 2195
rect 12830 2125 12834 2185
rect 12886 2125 13144 2185
rect 13196 2125 13200 2185
rect 12830 2050 13200 2125
rect 30 2010 13200 2050
rect 30 1925 400 2010
rect 30 1865 34 1925
rect 86 1865 344 1925
rect 396 1865 400 1925
rect 30 1855 400 1865
rect 430 1925 800 2010
rect 430 1865 434 1925
rect 486 1865 744 1925
rect 796 1865 800 1925
rect 430 1855 800 1865
rect 830 1925 1200 2010
rect 830 1865 834 1925
rect 886 1865 1144 1925
rect 1196 1865 1200 1925
rect 830 1855 1200 1865
rect 1230 1925 1600 2010
rect 1230 1865 1234 1925
rect 1286 1865 1544 1925
rect 1596 1865 1600 1925
rect 1230 1855 1600 1865
rect 1630 1925 2000 2010
rect 1630 1865 1634 1925
rect 1686 1865 1944 1925
rect 1996 1865 2000 1925
rect 1630 1855 2000 1865
rect 2030 1925 2400 2010
rect 2030 1865 2034 1925
rect 2086 1865 2344 1925
rect 2396 1865 2400 1925
rect 2030 1855 2400 1865
rect 2430 1925 2800 2010
rect 2430 1865 2434 1925
rect 2486 1865 2744 1925
rect 2796 1865 2800 1925
rect 2430 1855 2800 1865
rect 2830 1925 3200 2010
rect 2830 1865 2834 1925
rect 2886 1865 3144 1925
rect 3196 1865 3200 1925
rect 2830 1855 3200 1865
rect 3230 1925 3600 2010
rect 3230 1865 3234 1925
rect 3286 1865 3544 1925
rect 3596 1865 3600 1925
rect 3230 1855 3600 1865
rect 3630 1925 4000 2010
rect 3630 1865 3634 1925
rect 3686 1865 3944 1925
rect 3996 1865 4000 1925
rect 3630 1855 4000 1865
rect 4030 1925 4400 2010
rect 4030 1865 4034 1925
rect 4086 1865 4344 1925
rect 4396 1865 4400 1925
rect 4030 1855 4400 1865
rect 4430 1925 4800 2010
rect 4430 1865 4434 1925
rect 4486 1865 4744 1925
rect 4796 1865 4800 1925
rect 4430 1855 4800 1865
rect 4830 1925 5200 2010
rect 4830 1865 4834 1925
rect 4886 1865 5144 1925
rect 5196 1865 5200 1925
rect 4830 1855 5200 1865
rect 5230 1925 5600 2010
rect 5230 1865 5234 1925
rect 5286 1865 5544 1925
rect 5596 1865 5600 1925
rect 5230 1855 5600 1865
rect 5630 1925 6000 2010
rect 5630 1865 5634 1925
rect 5686 1865 5944 1925
rect 5996 1865 6000 1925
rect 5630 1855 6000 1865
rect 6030 1925 6400 2010
rect 6030 1865 6034 1925
rect 6086 1865 6344 1925
rect 6396 1865 6400 1925
rect 6030 1855 6400 1865
rect 6430 1925 6800 2010
rect 6430 1865 6434 1925
rect 6486 1865 6744 1925
rect 6796 1865 6800 1925
rect 6430 1855 6800 1865
rect 6830 1925 7200 2010
rect 6830 1865 6834 1925
rect 6886 1865 7144 1925
rect 7196 1865 7200 1925
rect 6830 1855 7200 1865
rect 7230 1925 7600 2010
rect 7230 1865 7234 1925
rect 7286 1865 7544 1925
rect 7596 1865 7600 1925
rect 7230 1855 7600 1865
rect 7630 1925 8000 2010
rect 7630 1865 7634 1925
rect 7686 1865 7944 1925
rect 7996 1865 8000 1925
rect 7630 1855 8000 1865
rect 8030 1925 8400 2010
rect 8030 1865 8034 1925
rect 8086 1865 8344 1925
rect 8396 1865 8400 1925
rect 8030 1855 8400 1865
rect 8430 1925 8800 2010
rect 8430 1865 8434 1925
rect 8486 1865 8744 1925
rect 8796 1865 8800 1925
rect 8430 1855 8800 1865
rect 8830 1925 9200 2010
rect 8830 1865 8834 1925
rect 8886 1865 9144 1925
rect 9196 1865 9200 1925
rect 8830 1855 9200 1865
rect 9230 1925 9600 2010
rect 9230 1865 9234 1925
rect 9286 1865 9544 1925
rect 9596 1865 9600 1925
rect 9230 1855 9600 1865
rect 9630 1925 10000 2010
rect 9630 1865 9634 1925
rect 9686 1865 9944 1925
rect 9996 1865 10000 1925
rect 9630 1855 10000 1865
rect 10030 1925 10400 2010
rect 10030 1865 10034 1925
rect 10086 1865 10344 1925
rect 10396 1865 10400 1925
rect 10030 1855 10400 1865
rect 10430 1925 10800 2010
rect 10430 1865 10434 1925
rect 10486 1865 10744 1925
rect 10796 1865 10800 1925
rect 10430 1855 10800 1865
rect 10830 1925 11200 2010
rect 10830 1865 10834 1925
rect 10886 1865 11144 1925
rect 11196 1865 11200 1925
rect 10830 1855 11200 1865
rect 11230 1925 11600 2010
rect 11230 1865 11234 1925
rect 11286 1865 11544 1925
rect 11596 1865 11600 1925
rect 11230 1855 11600 1865
rect 11630 1925 12000 2010
rect 11630 1865 11634 1925
rect 11686 1865 11944 1925
rect 11996 1865 12000 1925
rect 11630 1855 12000 1865
rect 12030 1925 12400 2010
rect 12030 1865 12034 1925
rect 12086 1865 12344 1925
rect 12396 1865 12400 1925
rect 12030 1855 12400 1865
rect 12430 1925 12800 2010
rect 12430 1865 12434 1925
rect 12486 1865 12744 1925
rect 12796 1865 12800 1925
rect 12430 1855 12800 1865
rect 12830 1925 13200 2010
rect 12830 1865 12834 1925
rect 12886 1865 13144 1925
rect 13196 1865 13200 1925
rect 12830 1855 13200 1865
rect -330 1825 -324 1855
rect 30 1825 70 1855
rect 430 1825 470 1855
rect 830 1825 870 1855
rect 1230 1825 1270 1855
rect 1630 1825 1670 1855
rect 2030 1825 2070 1855
rect 2430 1825 2470 1855
rect 2830 1825 2870 1855
rect 3230 1825 3270 1855
rect 3630 1825 3670 1855
rect 4030 1825 4070 1855
rect 4430 1825 4470 1855
rect 4830 1825 4870 1855
rect 5230 1825 5270 1855
rect 5630 1825 5670 1855
rect 6030 1825 6070 1855
rect 6430 1825 6470 1855
rect 6830 1825 6870 1855
rect 7230 1825 7270 1855
rect 7630 1825 7670 1855
rect 8030 1825 8070 1855
rect 8430 1825 8470 1855
rect 8830 1825 8870 1855
rect 9230 1825 9270 1855
rect 9630 1825 9670 1855
rect 10030 1825 10070 1855
rect 10430 1825 10470 1855
rect 10830 1825 10870 1855
rect 11230 1825 11270 1855
rect 11630 1825 11670 1855
rect 12030 1825 12070 1855
rect 12430 1825 12470 1855
rect -330 1815 0 1825
rect -314 1755 -56 1815
rect -4 1755 0 1815
rect -330 1555 0 1755
rect -314 1495 -56 1555
rect -4 1495 0 1555
rect -330 1485 0 1495
rect 30 1815 400 1825
rect 30 1755 34 1815
rect 86 1755 344 1815
rect 396 1755 400 1815
rect 30 1680 400 1755
rect 430 1815 800 1825
rect 430 1755 434 1815
rect 486 1755 744 1815
rect 796 1755 800 1815
rect 430 1680 800 1755
rect 830 1815 1200 1825
rect 830 1755 834 1815
rect 886 1755 1144 1815
rect 1196 1755 1200 1815
rect 830 1680 1200 1755
rect 1230 1815 1600 1825
rect 1230 1755 1234 1815
rect 1286 1755 1544 1815
rect 1596 1755 1600 1815
rect 1230 1680 1600 1755
rect 1630 1815 2000 1825
rect 1630 1755 1634 1815
rect 1686 1755 1944 1815
rect 1996 1755 2000 1815
rect 1630 1680 2000 1755
rect 2030 1815 2400 1825
rect 2030 1755 2034 1815
rect 2086 1755 2344 1815
rect 2396 1755 2400 1815
rect 2030 1680 2400 1755
rect 2430 1815 2800 1825
rect 2430 1755 2434 1815
rect 2486 1755 2744 1815
rect 2796 1755 2800 1815
rect 2430 1680 2800 1755
rect 2830 1815 3200 1825
rect 2830 1755 2834 1815
rect 2886 1755 3144 1815
rect 3196 1755 3200 1815
rect 2830 1680 3200 1755
rect 3230 1815 3600 1825
rect 3230 1755 3234 1815
rect 3286 1755 3544 1815
rect 3596 1755 3600 1815
rect 3230 1680 3600 1755
rect 3630 1815 4000 1825
rect 3630 1755 3634 1815
rect 3686 1755 3944 1815
rect 3996 1755 4000 1815
rect 3630 1680 4000 1755
rect 4030 1815 4400 1825
rect 4030 1755 4034 1815
rect 4086 1755 4344 1815
rect 4396 1755 4400 1815
rect 4030 1680 4400 1755
rect 4430 1815 4800 1825
rect 4430 1755 4434 1815
rect 4486 1755 4744 1815
rect 4796 1755 4800 1815
rect 4430 1680 4800 1755
rect 4830 1815 5200 1825
rect 4830 1755 4834 1815
rect 4886 1755 5144 1815
rect 5196 1755 5200 1815
rect 4830 1680 5200 1755
rect 5230 1815 5600 1825
rect 5230 1755 5234 1815
rect 5286 1755 5544 1815
rect 5596 1755 5600 1815
rect 5230 1680 5600 1755
rect 5630 1815 6000 1825
rect 5630 1755 5634 1815
rect 5686 1755 5944 1815
rect 5996 1755 6000 1815
rect 5630 1680 6000 1755
rect 6030 1815 6400 1825
rect 6030 1755 6034 1815
rect 6086 1755 6344 1815
rect 6396 1755 6400 1815
rect 6030 1680 6400 1755
rect 6430 1815 6800 1825
rect 6430 1755 6434 1815
rect 6486 1755 6744 1815
rect 6796 1755 6800 1815
rect 6430 1680 6800 1755
rect 6830 1815 7200 1825
rect 6830 1755 6834 1815
rect 6886 1755 7144 1815
rect 7196 1755 7200 1815
rect 6830 1680 7200 1755
rect 7230 1815 7600 1825
rect 7230 1755 7234 1815
rect 7286 1755 7544 1815
rect 7596 1755 7600 1815
rect 7230 1680 7600 1755
rect 7630 1815 8000 1825
rect 7630 1755 7634 1815
rect 7686 1755 7944 1815
rect 7996 1755 8000 1815
rect 7630 1680 8000 1755
rect 8030 1815 8400 1825
rect 8030 1755 8034 1815
rect 8086 1755 8344 1815
rect 8396 1755 8400 1815
rect 8030 1680 8400 1755
rect 8430 1815 8800 1825
rect 8430 1755 8434 1815
rect 8486 1755 8744 1815
rect 8796 1755 8800 1815
rect 8430 1680 8800 1755
rect 8830 1815 9200 1825
rect 8830 1755 8834 1815
rect 8886 1755 9144 1815
rect 9196 1755 9200 1815
rect 8830 1680 9200 1755
rect 9230 1815 9600 1825
rect 9230 1755 9234 1815
rect 9286 1755 9544 1815
rect 9596 1755 9600 1815
rect 9230 1680 9600 1755
rect 9630 1815 10000 1825
rect 9630 1755 9634 1815
rect 9686 1755 9944 1815
rect 9996 1755 10000 1815
rect 9630 1680 10000 1755
rect 10030 1815 10400 1825
rect 10030 1755 10034 1815
rect 10086 1755 10344 1815
rect 10396 1755 10400 1815
rect 10030 1680 10400 1755
rect 10430 1815 10800 1825
rect 10430 1755 10434 1815
rect 10486 1755 10744 1815
rect 10796 1755 10800 1815
rect 10430 1680 10800 1755
rect 10830 1815 11200 1825
rect 10830 1755 10834 1815
rect 10886 1755 11144 1815
rect 11196 1755 11200 1815
rect 10830 1680 11200 1755
rect 11230 1815 11600 1825
rect 11230 1755 11234 1815
rect 11286 1755 11544 1815
rect 11596 1755 11600 1815
rect 11230 1680 11600 1755
rect 11630 1815 12000 1825
rect 11630 1755 11634 1815
rect 11686 1755 11944 1815
rect 11996 1755 12000 1815
rect 11630 1680 12000 1755
rect 12030 1815 12400 1825
rect 12030 1755 12034 1815
rect 12086 1755 12344 1815
rect 12396 1755 12400 1815
rect 12030 1680 12400 1755
rect 12430 1815 12800 1825
rect 12430 1755 12434 1815
rect 12486 1755 12744 1815
rect 12796 1755 12800 1815
rect 12430 1680 12800 1755
rect 12830 1815 13200 1825
rect 12830 1755 12834 1815
rect 12886 1755 13144 1815
rect 13196 1755 13200 1815
rect 12830 1680 13200 1755
rect 30 1640 13200 1680
rect 30 1555 400 1640
rect 30 1495 34 1555
rect 86 1495 344 1555
rect 396 1495 400 1555
rect 30 1485 400 1495
rect 430 1555 800 1640
rect 430 1495 434 1555
rect 486 1495 744 1555
rect 796 1495 800 1555
rect 430 1485 800 1495
rect 830 1555 1200 1640
rect 830 1495 834 1555
rect 886 1495 1144 1555
rect 1196 1495 1200 1555
rect 830 1485 1200 1495
rect 1230 1555 1600 1640
rect 1230 1495 1234 1555
rect 1286 1495 1544 1555
rect 1596 1495 1600 1555
rect 1230 1485 1600 1495
rect 1630 1555 2000 1640
rect 1630 1495 1634 1555
rect 1686 1495 1944 1555
rect 1996 1495 2000 1555
rect 1630 1485 2000 1495
rect 2030 1555 2400 1640
rect 2030 1495 2034 1555
rect 2086 1495 2344 1555
rect 2396 1495 2400 1555
rect 2030 1485 2400 1495
rect 2430 1555 2800 1640
rect 2430 1495 2434 1555
rect 2486 1495 2744 1555
rect 2796 1495 2800 1555
rect 2430 1485 2800 1495
rect 2830 1555 3200 1640
rect 2830 1495 2834 1555
rect 2886 1495 3144 1555
rect 3196 1495 3200 1555
rect 2830 1485 3200 1495
rect 3230 1555 3600 1640
rect 3230 1495 3234 1555
rect 3286 1495 3544 1555
rect 3596 1495 3600 1555
rect 3230 1485 3600 1495
rect 3630 1555 4000 1640
rect 3630 1495 3634 1555
rect 3686 1495 3944 1555
rect 3996 1495 4000 1555
rect 3630 1485 4000 1495
rect 4030 1555 4400 1640
rect 4030 1495 4034 1555
rect 4086 1495 4344 1555
rect 4396 1495 4400 1555
rect 4030 1485 4400 1495
rect 4430 1555 4800 1640
rect 4430 1495 4434 1555
rect 4486 1495 4744 1555
rect 4796 1495 4800 1555
rect 4430 1485 4800 1495
rect 4830 1555 5200 1640
rect 4830 1495 4834 1555
rect 4886 1495 5144 1555
rect 5196 1495 5200 1555
rect 4830 1485 5200 1495
rect 5230 1555 5600 1640
rect 5230 1495 5234 1555
rect 5286 1495 5544 1555
rect 5596 1495 5600 1555
rect 5230 1485 5600 1495
rect 5630 1555 6000 1640
rect 5630 1495 5634 1555
rect 5686 1495 5944 1555
rect 5996 1495 6000 1555
rect 5630 1485 6000 1495
rect 6030 1555 6400 1640
rect 6030 1495 6034 1555
rect 6086 1495 6344 1555
rect 6396 1495 6400 1555
rect 6030 1485 6400 1495
rect 6430 1555 6800 1640
rect 6430 1495 6434 1555
rect 6486 1495 6744 1555
rect 6796 1495 6800 1555
rect 6430 1485 6800 1495
rect 6830 1555 7200 1640
rect 6830 1495 6834 1555
rect 6886 1495 7144 1555
rect 7196 1495 7200 1555
rect 6830 1485 7200 1495
rect 7230 1555 7600 1640
rect 7230 1495 7234 1555
rect 7286 1495 7544 1555
rect 7596 1495 7600 1555
rect 7230 1485 7600 1495
rect 7630 1555 8000 1640
rect 7630 1495 7634 1555
rect 7686 1495 7944 1555
rect 7996 1495 8000 1555
rect 7630 1485 8000 1495
rect 8030 1555 8400 1640
rect 8030 1495 8034 1555
rect 8086 1495 8344 1555
rect 8396 1495 8400 1555
rect 8030 1485 8400 1495
rect 8430 1555 8800 1640
rect 8430 1495 8434 1555
rect 8486 1495 8744 1555
rect 8796 1495 8800 1555
rect 8430 1485 8800 1495
rect 8830 1555 9200 1640
rect 8830 1495 8834 1555
rect 8886 1495 9144 1555
rect 9196 1495 9200 1555
rect 8830 1485 9200 1495
rect 9230 1555 9600 1640
rect 9230 1495 9234 1555
rect 9286 1495 9544 1555
rect 9596 1495 9600 1555
rect 9230 1485 9600 1495
rect 9630 1555 10000 1640
rect 9630 1495 9634 1555
rect 9686 1495 9944 1555
rect 9996 1495 10000 1555
rect 9630 1485 10000 1495
rect 10030 1555 10400 1640
rect 10030 1495 10034 1555
rect 10086 1495 10344 1555
rect 10396 1495 10400 1555
rect 10030 1485 10400 1495
rect 10430 1555 10800 1640
rect 10430 1495 10434 1555
rect 10486 1495 10744 1555
rect 10796 1495 10800 1555
rect 10430 1485 10800 1495
rect 10830 1555 11200 1640
rect 10830 1495 10834 1555
rect 10886 1495 11144 1555
rect 11196 1495 11200 1555
rect 10830 1485 11200 1495
rect 11230 1555 11600 1640
rect 11230 1495 11234 1555
rect 11286 1495 11544 1555
rect 11596 1495 11600 1555
rect 11230 1485 11600 1495
rect 11630 1555 12000 1640
rect 11630 1495 11634 1555
rect 11686 1495 11944 1555
rect 11996 1495 12000 1555
rect 11630 1485 12000 1495
rect 12030 1555 12400 1640
rect 12030 1495 12034 1555
rect 12086 1495 12344 1555
rect 12396 1495 12400 1555
rect 12030 1485 12400 1495
rect 12430 1555 12800 1640
rect 12430 1495 12434 1555
rect 12486 1495 12744 1555
rect 12796 1495 12800 1555
rect 12430 1485 12800 1495
rect 12830 1555 13200 1640
rect 12830 1495 12834 1555
rect 12886 1495 13144 1555
rect 13196 1495 13200 1555
rect 12830 1485 13200 1495
rect -330 1455 -324 1485
rect 30 1455 70 1485
rect 430 1455 470 1485
rect 830 1455 870 1485
rect 1230 1455 1270 1485
rect 1630 1455 1670 1485
rect 2030 1455 2070 1485
rect 2430 1455 2470 1485
rect 2830 1455 2870 1485
rect 3230 1455 3270 1485
rect 3630 1455 3670 1485
rect 4030 1455 4070 1485
rect 4430 1455 4470 1485
rect 4830 1455 4870 1485
rect 5230 1455 5270 1485
rect 5630 1455 5670 1485
rect 6030 1455 6070 1485
rect 6430 1455 6470 1485
rect 6830 1455 6870 1485
rect 7230 1455 7270 1485
rect 7630 1455 7670 1485
rect 8030 1455 8070 1485
rect 8430 1455 8470 1485
rect 8830 1455 8870 1485
rect 9230 1455 9270 1485
rect 9630 1455 9670 1485
rect 10030 1455 10070 1485
rect 10430 1455 10470 1485
rect 10830 1455 10870 1485
rect 11230 1455 11270 1485
rect 11630 1455 11670 1485
rect 12030 1455 12070 1485
rect 12430 1455 12470 1485
rect -330 1445 0 1455
rect -314 1385 -56 1445
rect -4 1385 0 1445
rect -330 1185 0 1385
rect -314 1125 -56 1185
rect -4 1125 0 1185
rect -330 1115 0 1125
rect 30 1445 400 1455
rect 30 1385 34 1445
rect 86 1385 344 1445
rect 396 1385 400 1445
rect 30 1310 400 1385
rect 430 1445 800 1455
rect 430 1385 434 1445
rect 486 1385 744 1445
rect 796 1385 800 1445
rect 430 1310 800 1385
rect 830 1445 1200 1455
rect 830 1385 834 1445
rect 886 1385 1144 1445
rect 1196 1385 1200 1445
rect 830 1310 1200 1385
rect 1230 1445 1600 1455
rect 1230 1385 1234 1445
rect 1286 1385 1544 1445
rect 1596 1385 1600 1445
rect 1230 1310 1600 1385
rect 1630 1445 2000 1455
rect 1630 1385 1634 1445
rect 1686 1385 1944 1445
rect 1996 1385 2000 1445
rect 1630 1310 2000 1385
rect 2030 1445 2400 1455
rect 2030 1385 2034 1445
rect 2086 1385 2344 1445
rect 2396 1385 2400 1445
rect 2030 1310 2400 1385
rect 2430 1445 2800 1455
rect 2430 1385 2434 1445
rect 2486 1385 2744 1445
rect 2796 1385 2800 1445
rect 2430 1310 2800 1385
rect 2830 1445 3200 1455
rect 2830 1385 2834 1445
rect 2886 1385 3144 1445
rect 3196 1385 3200 1445
rect 2830 1310 3200 1385
rect 3230 1445 3600 1455
rect 3230 1385 3234 1445
rect 3286 1385 3544 1445
rect 3596 1385 3600 1445
rect 3230 1310 3600 1385
rect 3630 1445 4000 1455
rect 3630 1385 3634 1445
rect 3686 1385 3944 1445
rect 3996 1385 4000 1445
rect 3630 1310 4000 1385
rect 4030 1445 4400 1455
rect 4030 1385 4034 1445
rect 4086 1385 4344 1445
rect 4396 1385 4400 1445
rect 4030 1310 4400 1385
rect 4430 1445 4800 1455
rect 4430 1385 4434 1445
rect 4486 1385 4744 1445
rect 4796 1385 4800 1445
rect 4430 1310 4800 1385
rect 4830 1445 5200 1455
rect 4830 1385 4834 1445
rect 4886 1385 5144 1445
rect 5196 1385 5200 1445
rect 4830 1310 5200 1385
rect 5230 1445 5600 1455
rect 5230 1385 5234 1445
rect 5286 1385 5544 1445
rect 5596 1385 5600 1445
rect 5230 1310 5600 1385
rect 5630 1445 6000 1455
rect 5630 1385 5634 1445
rect 5686 1385 5944 1445
rect 5996 1385 6000 1445
rect 5630 1310 6000 1385
rect 6030 1445 6400 1455
rect 6030 1385 6034 1445
rect 6086 1385 6344 1445
rect 6396 1385 6400 1445
rect 6030 1310 6400 1385
rect 6430 1445 6800 1455
rect 6430 1385 6434 1445
rect 6486 1385 6744 1445
rect 6796 1385 6800 1445
rect 6430 1310 6800 1385
rect 6830 1445 7200 1455
rect 6830 1385 6834 1445
rect 6886 1385 7144 1445
rect 7196 1385 7200 1445
rect 6830 1310 7200 1385
rect 7230 1445 7600 1455
rect 7230 1385 7234 1445
rect 7286 1385 7544 1445
rect 7596 1385 7600 1445
rect 7230 1310 7600 1385
rect 7630 1445 8000 1455
rect 7630 1385 7634 1445
rect 7686 1385 7944 1445
rect 7996 1385 8000 1445
rect 7630 1310 8000 1385
rect 8030 1445 8400 1455
rect 8030 1385 8034 1445
rect 8086 1385 8344 1445
rect 8396 1385 8400 1445
rect 8030 1310 8400 1385
rect 8430 1445 8800 1455
rect 8430 1385 8434 1445
rect 8486 1385 8744 1445
rect 8796 1385 8800 1445
rect 8430 1310 8800 1385
rect 8830 1445 9200 1455
rect 8830 1385 8834 1445
rect 8886 1385 9144 1445
rect 9196 1385 9200 1445
rect 8830 1310 9200 1385
rect 9230 1445 9600 1455
rect 9230 1385 9234 1445
rect 9286 1385 9544 1445
rect 9596 1385 9600 1445
rect 9230 1310 9600 1385
rect 9630 1445 10000 1455
rect 9630 1385 9634 1445
rect 9686 1385 9944 1445
rect 9996 1385 10000 1445
rect 9630 1310 10000 1385
rect 10030 1445 10400 1455
rect 10030 1385 10034 1445
rect 10086 1385 10344 1445
rect 10396 1385 10400 1445
rect 10030 1310 10400 1385
rect 10430 1445 10800 1455
rect 10430 1385 10434 1445
rect 10486 1385 10744 1445
rect 10796 1385 10800 1445
rect 10430 1310 10800 1385
rect 10830 1445 11200 1455
rect 10830 1385 10834 1445
rect 10886 1385 11144 1445
rect 11196 1385 11200 1445
rect 10830 1310 11200 1385
rect 11230 1445 11600 1455
rect 11230 1385 11234 1445
rect 11286 1385 11544 1445
rect 11596 1385 11600 1445
rect 11230 1310 11600 1385
rect 11630 1445 12000 1455
rect 11630 1385 11634 1445
rect 11686 1385 11944 1445
rect 11996 1385 12000 1445
rect 11630 1310 12000 1385
rect 12030 1445 12400 1455
rect 12030 1385 12034 1445
rect 12086 1385 12344 1445
rect 12396 1385 12400 1445
rect 12030 1310 12400 1385
rect 12430 1445 12800 1455
rect 12430 1385 12434 1445
rect 12486 1385 12744 1445
rect 12796 1385 12800 1445
rect 12430 1310 12800 1385
rect 12830 1445 13200 1455
rect 12830 1385 12834 1445
rect 12886 1385 13144 1445
rect 13196 1385 13200 1445
rect 12830 1310 13200 1385
rect 30 1270 13200 1310
rect 30 1185 400 1270
rect 30 1125 34 1185
rect 86 1125 344 1185
rect 396 1125 400 1185
rect 30 1115 400 1125
rect 430 1185 800 1270
rect 430 1125 434 1185
rect 486 1125 744 1185
rect 796 1125 800 1185
rect 430 1115 800 1125
rect 830 1185 1200 1270
rect 830 1125 834 1185
rect 886 1125 1144 1185
rect 1196 1125 1200 1185
rect 830 1115 1200 1125
rect 1230 1185 1600 1270
rect 1230 1125 1234 1185
rect 1286 1125 1544 1185
rect 1596 1125 1600 1185
rect 1230 1115 1600 1125
rect 1630 1185 2000 1270
rect 1630 1125 1634 1185
rect 1686 1125 1944 1185
rect 1996 1125 2000 1185
rect 1630 1115 2000 1125
rect 2030 1185 2400 1270
rect 2030 1125 2034 1185
rect 2086 1125 2344 1185
rect 2396 1125 2400 1185
rect 2030 1115 2400 1125
rect 2430 1185 2800 1270
rect 2430 1125 2434 1185
rect 2486 1125 2744 1185
rect 2796 1125 2800 1185
rect 2430 1115 2800 1125
rect 2830 1185 3200 1270
rect 2830 1125 2834 1185
rect 2886 1125 3144 1185
rect 3196 1125 3200 1185
rect 2830 1115 3200 1125
rect 3230 1185 3600 1270
rect 3230 1125 3234 1185
rect 3286 1125 3544 1185
rect 3596 1125 3600 1185
rect 3230 1115 3600 1125
rect 3630 1185 4000 1270
rect 3630 1125 3634 1185
rect 3686 1125 3944 1185
rect 3996 1125 4000 1185
rect 3630 1115 4000 1125
rect 4030 1185 4400 1270
rect 4030 1125 4034 1185
rect 4086 1125 4344 1185
rect 4396 1125 4400 1185
rect 4030 1115 4400 1125
rect 4430 1185 4800 1270
rect 4430 1125 4434 1185
rect 4486 1125 4744 1185
rect 4796 1125 4800 1185
rect 4430 1115 4800 1125
rect 4830 1185 5200 1270
rect 4830 1125 4834 1185
rect 4886 1125 5144 1185
rect 5196 1125 5200 1185
rect 4830 1115 5200 1125
rect 5230 1185 5600 1270
rect 5230 1125 5234 1185
rect 5286 1125 5544 1185
rect 5596 1125 5600 1185
rect 5230 1115 5600 1125
rect 5630 1185 6000 1270
rect 5630 1125 5634 1185
rect 5686 1125 5944 1185
rect 5996 1125 6000 1185
rect 5630 1115 6000 1125
rect 6030 1185 6400 1270
rect 6030 1125 6034 1185
rect 6086 1125 6344 1185
rect 6396 1125 6400 1185
rect 6030 1115 6400 1125
rect 6430 1185 6800 1270
rect 6430 1125 6434 1185
rect 6486 1125 6744 1185
rect 6796 1125 6800 1185
rect 6430 1115 6800 1125
rect 6830 1185 7200 1270
rect 6830 1125 6834 1185
rect 6886 1125 7144 1185
rect 7196 1125 7200 1185
rect 6830 1115 7200 1125
rect 7230 1185 7600 1270
rect 7230 1125 7234 1185
rect 7286 1125 7544 1185
rect 7596 1125 7600 1185
rect 7230 1115 7600 1125
rect 7630 1185 8000 1270
rect 7630 1125 7634 1185
rect 7686 1125 7944 1185
rect 7996 1125 8000 1185
rect 7630 1115 8000 1125
rect 8030 1185 8400 1270
rect 8030 1125 8034 1185
rect 8086 1125 8344 1185
rect 8396 1125 8400 1185
rect 8030 1115 8400 1125
rect 8430 1185 8800 1270
rect 8430 1125 8434 1185
rect 8486 1125 8744 1185
rect 8796 1125 8800 1185
rect 8430 1115 8800 1125
rect 8830 1185 9200 1270
rect 8830 1125 8834 1185
rect 8886 1125 9144 1185
rect 9196 1125 9200 1185
rect 8830 1115 9200 1125
rect 9230 1185 9600 1270
rect 9230 1125 9234 1185
rect 9286 1125 9544 1185
rect 9596 1125 9600 1185
rect 9230 1115 9600 1125
rect 9630 1185 10000 1270
rect 9630 1125 9634 1185
rect 9686 1125 9944 1185
rect 9996 1125 10000 1185
rect 9630 1115 10000 1125
rect 10030 1185 10400 1270
rect 10030 1125 10034 1185
rect 10086 1125 10344 1185
rect 10396 1125 10400 1185
rect 10030 1115 10400 1125
rect 10430 1185 10800 1270
rect 10430 1125 10434 1185
rect 10486 1125 10744 1185
rect 10796 1125 10800 1185
rect 10430 1115 10800 1125
rect 10830 1185 11200 1270
rect 10830 1125 10834 1185
rect 10886 1125 11144 1185
rect 11196 1125 11200 1185
rect 10830 1115 11200 1125
rect 11230 1185 11600 1270
rect 11230 1125 11234 1185
rect 11286 1125 11544 1185
rect 11596 1125 11600 1185
rect 11230 1115 11600 1125
rect 11630 1185 12000 1270
rect 11630 1125 11634 1185
rect 11686 1125 11944 1185
rect 11996 1125 12000 1185
rect 11630 1115 12000 1125
rect 12030 1185 12400 1270
rect 12030 1125 12034 1185
rect 12086 1125 12344 1185
rect 12396 1125 12400 1185
rect 12030 1115 12400 1125
rect 12430 1185 12800 1270
rect 12430 1125 12434 1185
rect 12486 1125 12744 1185
rect 12796 1125 12800 1185
rect 12430 1115 12800 1125
rect 12830 1185 13200 1270
rect 12830 1125 12834 1185
rect 12886 1125 13144 1185
rect 13196 1125 13200 1185
rect 12830 1115 13200 1125
rect -330 1085 -324 1115
rect 30 1085 70 1115
rect 430 1085 470 1115
rect 830 1085 870 1115
rect 1230 1085 1270 1115
rect 1630 1085 1670 1115
rect 2030 1085 2070 1115
rect 2430 1085 2470 1115
rect 2830 1085 2870 1115
rect 3230 1085 3270 1115
rect 3630 1085 3670 1115
rect 4030 1085 4070 1115
rect 4430 1085 4470 1115
rect 4830 1085 4870 1115
rect 5230 1085 5270 1115
rect 5630 1085 5670 1115
rect 6030 1085 6070 1115
rect 6430 1085 6470 1115
rect 6830 1085 6870 1115
rect 7230 1085 7270 1115
rect 7630 1085 7670 1115
rect 8030 1085 8070 1115
rect 8430 1085 8470 1115
rect 8830 1085 8870 1115
rect 9230 1085 9270 1115
rect 9630 1085 9670 1115
rect 10030 1085 10070 1115
rect 10430 1085 10470 1115
rect 10830 1085 10870 1115
rect 11230 1085 11270 1115
rect 11630 1085 11670 1115
rect 12030 1085 12070 1115
rect 12430 1085 12470 1115
rect -330 1075 0 1085
rect -314 1015 -56 1075
rect -4 1015 0 1075
rect -330 815 0 1015
rect -314 755 -56 815
rect -4 755 0 815
rect -330 745 0 755
rect 30 1075 400 1085
rect 30 1015 34 1075
rect 86 1015 344 1075
rect 396 1015 400 1075
rect 30 940 400 1015
rect 430 1075 800 1085
rect 430 1015 434 1075
rect 486 1015 744 1075
rect 796 1015 800 1075
rect 430 940 800 1015
rect 830 1075 1200 1085
rect 830 1015 834 1075
rect 886 1015 1144 1075
rect 1196 1015 1200 1075
rect 830 940 1200 1015
rect 1230 1075 1600 1085
rect 1230 1015 1234 1075
rect 1286 1015 1544 1075
rect 1596 1015 1600 1075
rect 1230 940 1600 1015
rect 1630 1075 2000 1085
rect 1630 1015 1634 1075
rect 1686 1015 1944 1075
rect 1996 1015 2000 1075
rect 1630 940 2000 1015
rect 2030 1075 2400 1085
rect 2030 1015 2034 1075
rect 2086 1015 2344 1075
rect 2396 1015 2400 1075
rect 2030 940 2400 1015
rect 2430 1075 2800 1085
rect 2430 1015 2434 1075
rect 2486 1015 2744 1075
rect 2796 1015 2800 1075
rect 2430 940 2800 1015
rect 2830 1075 3200 1085
rect 2830 1015 2834 1075
rect 2886 1015 3144 1075
rect 3196 1015 3200 1075
rect 2830 940 3200 1015
rect 3230 1075 3600 1085
rect 3230 1015 3234 1075
rect 3286 1015 3544 1075
rect 3596 1015 3600 1075
rect 3230 940 3600 1015
rect 3630 1075 4000 1085
rect 3630 1015 3634 1075
rect 3686 1015 3944 1075
rect 3996 1015 4000 1075
rect 3630 940 4000 1015
rect 4030 1075 4400 1085
rect 4030 1015 4034 1075
rect 4086 1015 4344 1075
rect 4396 1015 4400 1075
rect 4030 940 4400 1015
rect 4430 1075 4800 1085
rect 4430 1015 4434 1075
rect 4486 1015 4744 1075
rect 4796 1015 4800 1075
rect 4430 940 4800 1015
rect 4830 1075 5200 1085
rect 4830 1015 4834 1075
rect 4886 1015 5144 1075
rect 5196 1015 5200 1075
rect 4830 940 5200 1015
rect 5230 1075 5600 1085
rect 5230 1015 5234 1075
rect 5286 1015 5544 1075
rect 5596 1015 5600 1075
rect 5230 940 5600 1015
rect 5630 1075 6000 1085
rect 5630 1015 5634 1075
rect 5686 1015 5944 1075
rect 5996 1015 6000 1075
rect 5630 940 6000 1015
rect 6030 1075 6400 1085
rect 6030 1015 6034 1075
rect 6086 1015 6344 1075
rect 6396 1015 6400 1075
rect 6030 940 6400 1015
rect 6430 1075 6800 1085
rect 6430 1015 6434 1075
rect 6486 1015 6744 1075
rect 6796 1015 6800 1075
rect 6430 940 6800 1015
rect 6830 1075 7200 1085
rect 6830 1015 6834 1075
rect 6886 1015 7144 1075
rect 7196 1015 7200 1075
rect 6830 940 7200 1015
rect 7230 1075 7600 1085
rect 7230 1015 7234 1075
rect 7286 1015 7544 1075
rect 7596 1015 7600 1075
rect 7230 940 7600 1015
rect 7630 1075 8000 1085
rect 7630 1015 7634 1075
rect 7686 1015 7944 1075
rect 7996 1015 8000 1075
rect 7630 940 8000 1015
rect 8030 1075 8400 1085
rect 8030 1015 8034 1075
rect 8086 1015 8344 1075
rect 8396 1015 8400 1075
rect 8030 940 8400 1015
rect 8430 1075 8800 1085
rect 8430 1015 8434 1075
rect 8486 1015 8744 1075
rect 8796 1015 8800 1075
rect 8430 940 8800 1015
rect 8830 1075 9200 1085
rect 8830 1015 8834 1075
rect 8886 1015 9144 1075
rect 9196 1015 9200 1075
rect 8830 940 9200 1015
rect 9230 1075 9600 1085
rect 9230 1015 9234 1075
rect 9286 1015 9544 1075
rect 9596 1015 9600 1075
rect 9230 940 9600 1015
rect 9630 1075 10000 1085
rect 9630 1015 9634 1075
rect 9686 1015 9944 1075
rect 9996 1015 10000 1075
rect 9630 940 10000 1015
rect 10030 1075 10400 1085
rect 10030 1015 10034 1075
rect 10086 1015 10344 1075
rect 10396 1015 10400 1075
rect 10030 940 10400 1015
rect 10430 1075 10800 1085
rect 10430 1015 10434 1075
rect 10486 1015 10744 1075
rect 10796 1015 10800 1075
rect 10430 940 10800 1015
rect 10830 1075 11200 1085
rect 10830 1015 10834 1075
rect 10886 1015 11144 1075
rect 11196 1015 11200 1075
rect 10830 940 11200 1015
rect 11230 1075 11600 1085
rect 11230 1015 11234 1075
rect 11286 1015 11544 1075
rect 11596 1015 11600 1075
rect 11230 940 11600 1015
rect 11630 1075 12000 1085
rect 11630 1015 11634 1075
rect 11686 1015 11944 1075
rect 11996 1015 12000 1075
rect 11630 940 12000 1015
rect 12030 1075 12400 1085
rect 12030 1015 12034 1075
rect 12086 1015 12344 1075
rect 12396 1015 12400 1075
rect 12030 940 12400 1015
rect 12430 1075 12800 1085
rect 12430 1015 12434 1075
rect 12486 1015 12744 1075
rect 12796 1015 12800 1075
rect 12430 940 12800 1015
rect 12830 1075 13200 1085
rect 12830 1015 12834 1075
rect 12886 1015 13144 1075
rect 13196 1015 13200 1075
rect 12830 940 13200 1015
rect 30 900 13200 940
rect 30 815 400 900
rect 30 755 34 815
rect 86 755 344 815
rect 396 755 400 815
rect 30 745 400 755
rect 430 815 800 900
rect 430 755 434 815
rect 486 755 744 815
rect 796 755 800 815
rect 430 745 800 755
rect 830 815 1200 900
rect 830 755 834 815
rect 886 755 1144 815
rect 1196 755 1200 815
rect 830 745 1200 755
rect 1230 815 1600 900
rect 1230 755 1234 815
rect 1286 755 1544 815
rect 1596 755 1600 815
rect 1230 745 1600 755
rect 1630 815 2000 900
rect 1630 755 1634 815
rect 1686 755 1944 815
rect 1996 755 2000 815
rect 1630 745 2000 755
rect 2030 815 2400 900
rect 2030 755 2034 815
rect 2086 755 2344 815
rect 2396 755 2400 815
rect 2030 745 2400 755
rect 2430 815 2800 900
rect 2430 755 2434 815
rect 2486 755 2744 815
rect 2796 755 2800 815
rect 2430 745 2800 755
rect 2830 815 3200 900
rect 2830 755 2834 815
rect 2886 755 3144 815
rect 3196 755 3200 815
rect 2830 745 3200 755
rect 3230 815 3600 900
rect 3230 755 3234 815
rect 3286 755 3544 815
rect 3596 755 3600 815
rect 3230 745 3600 755
rect 3630 815 4000 900
rect 3630 755 3634 815
rect 3686 755 3944 815
rect 3996 755 4000 815
rect 3630 745 4000 755
rect 4030 815 4400 900
rect 4030 755 4034 815
rect 4086 755 4344 815
rect 4396 755 4400 815
rect 4030 745 4400 755
rect 4430 815 4800 900
rect 4430 755 4434 815
rect 4486 755 4744 815
rect 4796 755 4800 815
rect 4430 745 4800 755
rect 4830 815 5200 900
rect 4830 755 4834 815
rect 4886 755 5144 815
rect 5196 755 5200 815
rect 4830 745 5200 755
rect 5230 815 5600 900
rect 5230 755 5234 815
rect 5286 755 5544 815
rect 5596 755 5600 815
rect 5230 745 5600 755
rect 5630 815 6000 900
rect 5630 755 5634 815
rect 5686 755 5944 815
rect 5996 755 6000 815
rect 5630 745 6000 755
rect 6030 815 6400 900
rect 6030 755 6034 815
rect 6086 755 6344 815
rect 6396 755 6400 815
rect 6030 745 6400 755
rect 6430 815 6800 900
rect 6430 755 6434 815
rect 6486 755 6744 815
rect 6796 755 6800 815
rect 6430 745 6800 755
rect 6830 815 7200 900
rect 6830 755 6834 815
rect 6886 755 7144 815
rect 7196 755 7200 815
rect 6830 745 7200 755
rect 7230 815 7600 900
rect 7230 755 7234 815
rect 7286 755 7544 815
rect 7596 755 7600 815
rect 7230 745 7600 755
rect 7630 815 8000 900
rect 7630 755 7634 815
rect 7686 755 7944 815
rect 7996 755 8000 815
rect 7630 745 8000 755
rect 8030 815 8400 900
rect 8030 755 8034 815
rect 8086 755 8344 815
rect 8396 755 8400 815
rect 8030 745 8400 755
rect 8430 815 8800 900
rect 8430 755 8434 815
rect 8486 755 8744 815
rect 8796 755 8800 815
rect 8430 745 8800 755
rect 8830 815 9200 900
rect 8830 755 8834 815
rect 8886 755 9144 815
rect 9196 755 9200 815
rect 8830 745 9200 755
rect 9230 815 9600 900
rect 9230 755 9234 815
rect 9286 755 9544 815
rect 9596 755 9600 815
rect 9230 745 9600 755
rect 9630 815 10000 900
rect 9630 755 9634 815
rect 9686 755 9944 815
rect 9996 755 10000 815
rect 9630 745 10000 755
rect 10030 815 10400 900
rect 10030 755 10034 815
rect 10086 755 10344 815
rect 10396 755 10400 815
rect 10030 745 10400 755
rect 10430 815 10800 900
rect 10430 755 10434 815
rect 10486 755 10744 815
rect 10796 755 10800 815
rect 10430 745 10800 755
rect 10830 815 11200 900
rect 10830 755 10834 815
rect 10886 755 11144 815
rect 11196 755 11200 815
rect 10830 745 11200 755
rect 11230 815 11600 900
rect 11230 755 11234 815
rect 11286 755 11544 815
rect 11596 755 11600 815
rect 11230 745 11600 755
rect 11630 815 12000 900
rect 11630 755 11634 815
rect 11686 755 11944 815
rect 11996 755 12000 815
rect 11630 745 12000 755
rect 12030 815 12400 900
rect 12030 755 12034 815
rect 12086 755 12344 815
rect 12396 755 12400 815
rect 12030 745 12400 755
rect 12430 815 12800 900
rect 12430 755 12434 815
rect 12486 755 12744 815
rect 12796 755 12800 815
rect 12430 745 12800 755
rect 12830 815 13200 900
rect 12830 755 12834 815
rect 12886 755 13144 815
rect 13196 755 13200 815
rect 12830 745 13200 755
rect -330 715 -324 745
rect 30 715 70 745
rect 430 715 470 745
rect 830 715 870 745
rect 1230 715 1270 745
rect 1630 715 1670 745
rect 2030 715 2070 745
rect 2430 715 2470 745
rect 2830 715 2870 745
rect 3230 715 3270 745
rect 3630 715 3670 745
rect 4030 715 4070 745
rect 4430 715 4470 745
rect 4830 715 4870 745
rect 5230 715 5270 745
rect 5630 715 5670 745
rect 6030 715 6070 745
rect 6430 715 6470 745
rect 6830 715 6870 745
rect 7230 715 7270 745
rect 7630 715 7670 745
rect 8030 715 8070 745
rect 8430 715 8470 745
rect 8830 715 8870 745
rect 9230 715 9270 745
rect 9630 715 9670 745
rect 10030 715 10070 745
rect 10430 715 10470 745
rect 10830 715 10870 745
rect 11230 715 11270 745
rect 11630 715 11670 745
rect 12030 715 12070 745
rect 12430 715 12470 745
rect -330 705 0 715
rect -314 645 -56 705
rect -4 645 0 705
rect -330 445 0 645
rect -314 385 -56 445
rect -4 385 0 445
rect -330 375 0 385
rect 30 705 400 715
rect 30 645 34 705
rect 86 645 344 705
rect 396 645 400 705
rect 30 570 400 645
rect 430 705 800 715
rect 430 645 434 705
rect 486 645 744 705
rect 796 645 800 705
rect 430 570 800 645
rect 830 705 1200 715
rect 830 645 834 705
rect 886 645 1144 705
rect 1196 645 1200 705
rect 830 570 1200 645
rect 1230 705 1600 715
rect 1230 645 1234 705
rect 1286 645 1544 705
rect 1596 645 1600 705
rect 1230 570 1600 645
rect 1630 705 2000 715
rect 1630 645 1634 705
rect 1686 645 1944 705
rect 1996 645 2000 705
rect 1630 570 2000 645
rect 2030 705 2400 715
rect 2030 645 2034 705
rect 2086 645 2344 705
rect 2396 645 2400 705
rect 2030 570 2400 645
rect 2430 705 2800 715
rect 2430 645 2434 705
rect 2486 645 2744 705
rect 2796 645 2800 705
rect 2430 570 2800 645
rect 2830 705 3200 715
rect 2830 645 2834 705
rect 2886 645 3144 705
rect 3196 645 3200 705
rect 2830 570 3200 645
rect 3230 705 3600 715
rect 3230 645 3234 705
rect 3286 645 3544 705
rect 3596 645 3600 705
rect 3230 570 3600 645
rect 3630 705 4000 715
rect 3630 645 3634 705
rect 3686 645 3944 705
rect 3996 645 4000 705
rect 3630 570 4000 645
rect 4030 705 4400 715
rect 4030 645 4034 705
rect 4086 645 4344 705
rect 4396 645 4400 705
rect 4030 570 4400 645
rect 4430 705 4800 715
rect 4430 645 4434 705
rect 4486 645 4744 705
rect 4796 645 4800 705
rect 4430 570 4800 645
rect 4830 705 5200 715
rect 4830 645 4834 705
rect 4886 645 5144 705
rect 5196 645 5200 705
rect 4830 570 5200 645
rect 5230 705 5600 715
rect 5230 645 5234 705
rect 5286 645 5544 705
rect 5596 645 5600 705
rect 5230 570 5600 645
rect 5630 705 6000 715
rect 5630 645 5634 705
rect 5686 645 5944 705
rect 5996 645 6000 705
rect 5630 570 6000 645
rect 6030 705 6400 715
rect 6030 645 6034 705
rect 6086 645 6344 705
rect 6396 645 6400 705
rect 6030 570 6400 645
rect 6430 705 6800 715
rect 6430 645 6434 705
rect 6486 645 6744 705
rect 6796 645 6800 705
rect 6430 570 6800 645
rect 6830 705 7200 715
rect 6830 645 6834 705
rect 6886 645 7144 705
rect 7196 645 7200 705
rect 6830 570 7200 645
rect 7230 705 7600 715
rect 7230 645 7234 705
rect 7286 645 7544 705
rect 7596 645 7600 705
rect 7230 570 7600 645
rect 7630 705 8000 715
rect 7630 645 7634 705
rect 7686 645 7944 705
rect 7996 645 8000 705
rect 7630 570 8000 645
rect 8030 705 8400 715
rect 8030 645 8034 705
rect 8086 645 8344 705
rect 8396 645 8400 705
rect 8030 570 8400 645
rect 8430 705 8800 715
rect 8430 645 8434 705
rect 8486 645 8744 705
rect 8796 645 8800 705
rect 8430 570 8800 645
rect 8830 705 9200 715
rect 8830 645 8834 705
rect 8886 645 9144 705
rect 9196 645 9200 705
rect 8830 570 9200 645
rect 9230 705 9600 715
rect 9230 645 9234 705
rect 9286 645 9544 705
rect 9596 645 9600 705
rect 9230 570 9600 645
rect 9630 705 10000 715
rect 9630 645 9634 705
rect 9686 645 9944 705
rect 9996 645 10000 705
rect 9630 570 10000 645
rect 10030 705 10400 715
rect 10030 645 10034 705
rect 10086 645 10344 705
rect 10396 645 10400 705
rect 10030 570 10400 645
rect 10430 705 10800 715
rect 10430 645 10434 705
rect 10486 645 10744 705
rect 10796 645 10800 705
rect 10430 570 10800 645
rect 10830 705 11200 715
rect 10830 645 10834 705
rect 10886 645 11144 705
rect 11196 645 11200 705
rect 10830 570 11200 645
rect 11230 705 11600 715
rect 11230 645 11234 705
rect 11286 645 11544 705
rect 11596 645 11600 705
rect 11230 570 11600 645
rect 11630 705 12000 715
rect 11630 645 11634 705
rect 11686 645 11944 705
rect 11996 645 12000 705
rect 11630 570 12000 645
rect 12030 705 12400 715
rect 12030 645 12034 705
rect 12086 645 12344 705
rect 12396 645 12400 705
rect 12030 570 12400 645
rect 12430 705 12800 715
rect 12430 645 12434 705
rect 12486 645 12744 705
rect 12796 645 12800 705
rect 12430 570 12800 645
rect 12830 705 13200 715
rect 12830 645 12834 705
rect 12886 645 13144 705
rect 13196 645 13200 705
rect 12830 570 13200 645
rect 30 530 13200 570
rect 30 445 400 530
rect 30 385 34 445
rect 86 385 344 445
rect 396 385 400 445
rect 30 375 400 385
rect 430 445 800 530
rect 430 385 434 445
rect 486 385 744 445
rect 796 385 800 445
rect 430 375 800 385
rect 830 445 1200 530
rect 830 385 834 445
rect 886 385 1144 445
rect 1196 385 1200 445
rect 830 375 1200 385
rect 1230 445 1600 530
rect 1230 385 1234 445
rect 1286 385 1544 445
rect 1596 385 1600 445
rect 1230 375 1600 385
rect 1630 445 2000 530
rect 1630 385 1634 445
rect 1686 385 1944 445
rect 1996 385 2000 445
rect 1630 375 2000 385
rect 2030 445 2400 530
rect 2030 385 2034 445
rect 2086 385 2344 445
rect 2396 385 2400 445
rect 2030 375 2400 385
rect 2430 445 2800 530
rect 2430 385 2434 445
rect 2486 385 2744 445
rect 2796 385 2800 445
rect 2430 375 2800 385
rect 2830 445 3200 530
rect 2830 385 2834 445
rect 2886 385 3144 445
rect 3196 385 3200 445
rect 2830 375 3200 385
rect 3230 445 3600 530
rect 3230 385 3234 445
rect 3286 385 3544 445
rect 3596 385 3600 445
rect 3230 375 3600 385
rect 3630 445 4000 530
rect 3630 385 3634 445
rect 3686 385 3944 445
rect 3996 385 4000 445
rect 3630 375 4000 385
rect 4030 445 4400 530
rect 4030 385 4034 445
rect 4086 385 4344 445
rect 4396 385 4400 445
rect 4030 375 4400 385
rect 4430 445 4800 530
rect 4430 385 4434 445
rect 4486 385 4744 445
rect 4796 385 4800 445
rect 4430 375 4800 385
rect 4830 445 5200 530
rect 4830 385 4834 445
rect 4886 385 5144 445
rect 5196 385 5200 445
rect 4830 375 5200 385
rect 5230 445 5600 530
rect 5230 385 5234 445
rect 5286 385 5544 445
rect 5596 385 5600 445
rect 5230 375 5600 385
rect 5630 445 6000 530
rect 5630 385 5634 445
rect 5686 385 5944 445
rect 5996 385 6000 445
rect 5630 375 6000 385
rect 6030 445 6400 530
rect 6030 385 6034 445
rect 6086 385 6344 445
rect 6396 385 6400 445
rect 6030 375 6400 385
rect 6430 445 6800 530
rect 6430 385 6434 445
rect 6486 385 6744 445
rect 6796 385 6800 445
rect 6430 375 6800 385
rect 6830 445 7200 530
rect 6830 385 6834 445
rect 6886 385 7144 445
rect 7196 385 7200 445
rect 6830 375 7200 385
rect 7230 445 7600 530
rect 7230 385 7234 445
rect 7286 385 7544 445
rect 7596 385 7600 445
rect 7230 375 7600 385
rect 7630 445 8000 530
rect 7630 385 7634 445
rect 7686 385 7944 445
rect 7996 385 8000 445
rect 7630 375 8000 385
rect 8030 445 8400 530
rect 8030 385 8034 445
rect 8086 385 8344 445
rect 8396 385 8400 445
rect 8030 375 8400 385
rect 8430 445 8800 530
rect 8430 385 8434 445
rect 8486 385 8744 445
rect 8796 385 8800 445
rect 8430 375 8800 385
rect 8830 445 9200 530
rect 8830 385 8834 445
rect 8886 385 9144 445
rect 9196 385 9200 445
rect 8830 375 9200 385
rect 9230 445 9600 530
rect 9230 385 9234 445
rect 9286 385 9544 445
rect 9596 385 9600 445
rect 9230 375 9600 385
rect 9630 445 10000 530
rect 9630 385 9634 445
rect 9686 385 9944 445
rect 9996 385 10000 445
rect 9630 375 10000 385
rect 10030 445 10400 530
rect 10030 385 10034 445
rect 10086 385 10344 445
rect 10396 385 10400 445
rect 10030 375 10400 385
rect 10430 445 10800 530
rect 10430 385 10434 445
rect 10486 385 10744 445
rect 10796 385 10800 445
rect 10430 375 10800 385
rect 10830 445 11200 530
rect 10830 385 10834 445
rect 10886 385 11144 445
rect 11196 385 11200 445
rect 10830 375 11200 385
rect 11230 445 11600 530
rect 11230 385 11234 445
rect 11286 385 11544 445
rect 11596 385 11600 445
rect 11230 375 11600 385
rect 11630 445 12000 530
rect 11630 385 11634 445
rect 11686 385 11944 445
rect 11996 385 12000 445
rect 11630 375 12000 385
rect 12030 445 12400 530
rect 12030 385 12034 445
rect 12086 385 12344 445
rect 12396 385 12400 445
rect 12030 375 12400 385
rect 12430 445 12800 530
rect 12430 385 12434 445
rect 12486 385 12744 445
rect 12796 385 12800 445
rect 12430 375 12800 385
rect 12830 445 13200 530
rect 12830 385 12834 445
rect 12886 385 13144 445
rect 13196 385 13200 445
rect 12830 375 13200 385
rect -330 345 -324 375
rect 30 345 70 375
rect 430 345 470 375
rect 830 345 870 375
rect 1230 345 1270 375
rect 1630 345 1670 375
rect 2030 345 2070 375
rect 2430 345 2470 375
rect 2830 345 2870 375
rect 3230 345 3270 375
rect 3630 345 3670 375
rect 4030 345 4070 375
rect 4430 345 4470 375
rect 4830 345 4870 375
rect 5230 345 5270 375
rect 5630 345 5670 375
rect 6030 345 6070 375
rect 6430 345 6470 375
rect 6830 345 6870 375
rect 7230 345 7270 375
rect 7630 345 7670 375
rect 8030 345 8070 375
rect 8430 345 8470 375
rect 8830 345 8870 375
rect 9230 345 9270 375
rect 9630 345 9670 375
rect 10030 345 10070 375
rect 10430 345 10470 375
rect 10830 345 10870 375
rect 11230 345 11270 375
rect 11630 345 11670 375
rect 12030 345 12070 375
rect 12430 345 12470 375
rect -330 335 0 345
rect -314 275 -56 335
rect -4 275 0 335
rect -330 75 0 275
rect -314 15 -56 75
rect -4 15 0 75
rect -330 5 0 15
rect 30 335 400 345
rect 30 275 34 335
rect 86 275 344 335
rect 396 275 400 335
rect 30 200 400 275
rect 430 335 800 345
rect 430 275 434 335
rect 486 275 744 335
rect 796 275 800 335
rect 430 200 800 275
rect 830 335 1200 345
rect 830 275 834 335
rect 886 275 1144 335
rect 1196 275 1200 335
rect 830 200 1200 275
rect 1230 335 1600 345
rect 1230 275 1234 335
rect 1286 275 1544 335
rect 1596 275 1600 335
rect 1230 200 1600 275
rect 1630 335 2000 345
rect 1630 275 1634 335
rect 1686 275 1944 335
rect 1996 275 2000 335
rect 1630 200 2000 275
rect 2030 335 2400 345
rect 2030 275 2034 335
rect 2086 275 2344 335
rect 2396 275 2400 335
rect 2030 200 2400 275
rect 2430 335 2800 345
rect 2430 275 2434 335
rect 2486 275 2744 335
rect 2796 275 2800 335
rect 2430 200 2800 275
rect 2830 335 3200 345
rect 2830 275 2834 335
rect 2886 275 3144 335
rect 3196 275 3200 335
rect 2830 200 3200 275
rect 3230 335 3600 345
rect 3230 275 3234 335
rect 3286 275 3544 335
rect 3596 275 3600 335
rect 3230 200 3600 275
rect 3630 335 4000 345
rect 3630 275 3634 335
rect 3686 275 3944 335
rect 3996 275 4000 335
rect 3630 200 4000 275
rect 4030 335 4400 345
rect 4030 275 4034 335
rect 4086 275 4344 335
rect 4396 275 4400 335
rect 4030 200 4400 275
rect 4430 335 4800 345
rect 4430 275 4434 335
rect 4486 275 4744 335
rect 4796 275 4800 335
rect 4430 200 4800 275
rect 4830 335 5200 345
rect 4830 275 4834 335
rect 4886 275 5144 335
rect 5196 275 5200 335
rect 4830 200 5200 275
rect 5230 335 5600 345
rect 5230 275 5234 335
rect 5286 275 5544 335
rect 5596 275 5600 335
rect 5230 200 5600 275
rect 5630 335 6000 345
rect 5630 275 5634 335
rect 5686 275 5944 335
rect 5996 275 6000 335
rect 5630 200 6000 275
rect 6030 335 6400 345
rect 6030 275 6034 335
rect 6086 275 6344 335
rect 6396 275 6400 335
rect 6030 200 6400 275
rect 6430 335 6800 345
rect 6430 275 6434 335
rect 6486 275 6744 335
rect 6796 275 6800 335
rect 6430 200 6800 275
rect 6830 335 7200 345
rect 6830 275 6834 335
rect 6886 275 7144 335
rect 7196 275 7200 335
rect 6830 200 7200 275
rect 7230 335 7600 345
rect 7230 275 7234 335
rect 7286 275 7544 335
rect 7596 275 7600 335
rect 7230 200 7600 275
rect 7630 335 8000 345
rect 7630 275 7634 335
rect 7686 275 7944 335
rect 7996 275 8000 335
rect 7630 200 8000 275
rect 8030 335 8400 345
rect 8030 275 8034 335
rect 8086 275 8344 335
rect 8396 275 8400 335
rect 8030 200 8400 275
rect 8430 335 8800 345
rect 8430 275 8434 335
rect 8486 275 8744 335
rect 8796 275 8800 335
rect 8430 200 8800 275
rect 8830 335 9200 345
rect 8830 275 8834 335
rect 8886 275 9144 335
rect 9196 275 9200 335
rect 8830 200 9200 275
rect 9230 335 9600 345
rect 9230 275 9234 335
rect 9286 275 9544 335
rect 9596 275 9600 335
rect 9230 200 9600 275
rect 9630 335 10000 345
rect 9630 275 9634 335
rect 9686 275 9944 335
rect 9996 275 10000 335
rect 9630 200 10000 275
rect 10030 335 10400 345
rect 10030 275 10034 335
rect 10086 275 10344 335
rect 10396 275 10400 335
rect 10030 200 10400 275
rect 10430 335 10800 345
rect 10430 275 10434 335
rect 10486 275 10744 335
rect 10796 275 10800 335
rect 10430 200 10800 275
rect 10830 335 11200 345
rect 10830 275 10834 335
rect 10886 275 11144 335
rect 11196 275 11200 335
rect 10830 200 11200 275
rect 11230 335 11600 345
rect 11230 275 11234 335
rect 11286 275 11544 335
rect 11596 275 11600 335
rect 11230 200 11600 275
rect 11630 335 12000 345
rect 11630 275 11634 335
rect 11686 275 11944 335
rect 11996 275 12000 335
rect 11630 200 12000 275
rect 12030 335 12400 345
rect 12030 275 12034 335
rect 12086 275 12344 335
rect 12396 275 12400 335
rect 12030 200 12400 275
rect 12430 335 12800 345
rect 12430 275 12434 335
rect 12486 275 12744 335
rect 12796 275 12800 335
rect 12430 200 12800 275
rect 12830 335 13200 345
rect 12830 275 12834 335
rect 12886 275 13144 335
rect 13196 275 13200 335
rect 12830 200 13200 275
rect 30 160 13200 200
rect 30 75 400 160
rect 30 15 34 75
rect 86 15 344 75
rect 396 15 400 75
rect 30 5 400 15
rect 430 75 800 160
rect 430 15 434 75
rect 486 15 744 75
rect 796 15 800 75
rect 430 5 800 15
rect 830 75 1200 160
rect 830 15 834 75
rect 886 15 1144 75
rect 1196 15 1200 75
rect 830 5 1200 15
rect 1230 75 1600 160
rect 1230 15 1234 75
rect 1286 15 1544 75
rect 1596 15 1600 75
rect 1230 5 1600 15
rect 1630 75 2000 160
rect 1630 15 1634 75
rect 1686 15 1944 75
rect 1996 15 2000 75
rect 1630 5 2000 15
rect 2030 75 2400 160
rect 2030 15 2034 75
rect 2086 15 2344 75
rect 2396 15 2400 75
rect 2030 5 2400 15
rect 2430 75 2800 160
rect 2430 15 2434 75
rect 2486 15 2744 75
rect 2796 15 2800 75
rect 2430 5 2800 15
rect 2830 75 3200 160
rect 2830 15 2834 75
rect 2886 15 3144 75
rect 3196 15 3200 75
rect 2830 5 3200 15
rect 3230 75 3600 160
rect 3230 15 3234 75
rect 3286 15 3544 75
rect 3596 15 3600 75
rect 3230 5 3600 15
rect 3630 75 4000 160
rect 3630 15 3634 75
rect 3686 15 3944 75
rect 3996 15 4000 75
rect 3630 5 4000 15
rect 4030 75 4400 160
rect 4030 15 4034 75
rect 4086 15 4344 75
rect 4396 15 4400 75
rect 4030 5 4400 15
rect 4430 75 4800 160
rect 4430 15 4434 75
rect 4486 15 4744 75
rect 4796 15 4800 75
rect 4430 5 4800 15
rect 4830 75 5200 160
rect 4830 15 4834 75
rect 4886 15 5144 75
rect 5196 15 5200 75
rect 4830 5 5200 15
rect 5230 75 5600 160
rect 5230 15 5234 75
rect 5286 15 5544 75
rect 5596 15 5600 75
rect 5230 5 5600 15
rect 5630 75 6000 160
rect 5630 15 5634 75
rect 5686 15 5944 75
rect 5996 15 6000 75
rect 5630 5 6000 15
rect 6030 75 6400 160
rect 6030 15 6034 75
rect 6086 15 6344 75
rect 6396 15 6400 75
rect 6030 5 6400 15
rect 6430 75 6800 160
rect 6430 15 6434 75
rect 6486 15 6744 75
rect 6796 15 6800 75
rect 6430 5 6800 15
rect 6830 75 7200 160
rect 6830 15 6834 75
rect 6886 15 7144 75
rect 7196 15 7200 75
rect 6830 5 7200 15
rect 7230 75 7600 160
rect 7230 15 7234 75
rect 7286 15 7544 75
rect 7596 15 7600 75
rect 7230 5 7600 15
rect 7630 75 8000 160
rect 7630 15 7634 75
rect 7686 15 7944 75
rect 7996 15 8000 75
rect 7630 5 8000 15
rect 8030 75 8400 160
rect 8030 15 8034 75
rect 8086 15 8344 75
rect 8396 15 8400 75
rect 8030 5 8400 15
rect 8430 75 8800 160
rect 8430 15 8434 75
rect 8486 15 8744 75
rect 8796 15 8800 75
rect 8430 5 8800 15
rect 8830 75 9200 160
rect 8830 15 8834 75
rect 8886 15 9144 75
rect 9196 15 9200 75
rect 8830 5 9200 15
rect 9230 75 9600 160
rect 9230 15 9234 75
rect 9286 15 9544 75
rect 9596 15 9600 75
rect 9230 5 9600 15
rect 9630 75 10000 160
rect 9630 15 9634 75
rect 9686 15 9944 75
rect 9996 15 10000 75
rect 9630 5 10000 15
rect 10030 75 10400 160
rect 10030 15 10034 75
rect 10086 15 10344 75
rect 10396 15 10400 75
rect 10030 5 10400 15
rect 10430 75 10800 160
rect 10430 15 10434 75
rect 10486 15 10744 75
rect 10796 15 10800 75
rect 10430 5 10800 15
rect 10830 75 11200 160
rect 10830 15 10834 75
rect 10886 15 11144 75
rect 11196 15 11200 75
rect 10830 5 11200 15
rect 11230 75 11600 160
rect 11230 15 11234 75
rect 11286 15 11544 75
rect 11596 15 11600 75
rect 11230 5 11600 15
rect 11630 75 12000 160
rect 11630 15 11634 75
rect 11686 15 11944 75
rect 11996 15 12000 75
rect 11630 5 12000 15
rect 12030 75 12400 160
rect 12030 15 12034 75
rect 12086 15 12344 75
rect 12396 15 12400 75
rect 12030 5 12400 15
rect 12430 75 12800 160
rect 12430 15 12434 75
rect 12486 15 12744 75
rect 12796 15 12800 75
rect 12430 5 12800 15
rect 12830 75 13200 160
rect 12830 15 12834 75
rect 12886 15 13144 75
rect 13196 15 13200 75
rect 12830 5 13200 15
rect -330 -25 -324 5
rect -330 -35 0 -25
rect -376 -95 -366 -50
rect -314 -95 -56 -35
rect -4 -95 0 -35
rect -376 -103 0 -95
rect -370 -164 0 -103
rect 30 -35 400 -25
rect 30 -95 34 -35
rect 86 -95 344 -35
rect 396 -95 400 -35
rect 30 -164 400 -95
rect 430 -35 800 -25
rect 430 -95 434 -35
rect 486 -95 744 -35
rect 796 -95 800 -35
rect 430 -164 800 -95
rect 830 -35 1200 -25
rect 830 -95 834 -35
rect 886 -95 1144 -35
rect 1196 -95 1200 -35
rect 830 -164 1200 -95
rect 1230 -35 1600 -25
rect 1230 -95 1234 -35
rect 1286 -95 1544 -35
rect 1596 -95 1600 -35
rect 1230 -164 1600 -95
rect 1630 -35 2000 -25
rect 1630 -95 1634 -35
rect 1686 -95 1944 -35
rect 1996 -95 2000 -35
rect 1630 -164 2000 -95
rect 2030 -35 2400 -25
rect 2030 -95 2034 -35
rect 2086 -95 2344 -35
rect 2396 -95 2400 -35
rect 2030 -164 2400 -95
rect 2430 -35 2800 -25
rect 2430 -95 2434 -35
rect 2486 -95 2744 -35
rect 2796 -95 2800 -35
rect 2430 -164 2800 -95
rect 2830 -35 3200 -25
rect 2830 -95 2834 -35
rect 2886 -95 3144 -35
rect 3196 -95 3200 -35
rect 2830 -164 3200 -95
rect 3230 -35 3600 -25
rect 3230 -95 3234 -35
rect 3286 -95 3544 -35
rect 3596 -95 3600 -35
rect 3230 -164 3600 -95
rect 3630 -35 4000 -25
rect 3630 -95 3634 -35
rect 3686 -95 3944 -35
rect 3996 -95 4000 -35
rect 3630 -164 4000 -95
rect 4030 -35 4400 -25
rect 4030 -95 4034 -35
rect 4086 -95 4344 -35
rect 4396 -95 4400 -35
rect 4030 -164 4400 -95
rect 4430 -35 4800 -25
rect 4430 -95 4434 -35
rect 4486 -95 4744 -35
rect 4796 -95 4800 -35
rect 4430 -164 4800 -95
rect 4830 -35 5200 -25
rect 4830 -95 4834 -35
rect 4886 -95 5144 -35
rect 5196 -95 5200 -35
rect 4830 -164 5200 -95
rect 5230 -35 5600 -25
rect 5230 -95 5234 -35
rect 5286 -95 5544 -35
rect 5596 -95 5600 -35
rect 5230 -164 5600 -95
rect 5630 -35 6000 -25
rect 5630 -95 5634 -35
rect 5686 -95 5944 -35
rect 5996 -95 6000 -35
rect 5630 -164 6000 -95
rect 6030 -35 6400 -25
rect 6030 -95 6034 -35
rect 6086 -95 6344 -35
rect 6396 -95 6400 -35
rect 6030 -164 6400 -95
rect 6430 -35 6800 -25
rect 6430 -95 6434 -35
rect 6486 -95 6744 -35
rect 6796 -95 6800 -35
rect 6430 -164 6800 -95
rect 6830 -35 7200 -25
rect 6830 -95 6834 -35
rect 6886 -95 7144 -35
rect 7196 -95 7200 -35
rect 6830 -164 7200 -95
rect 7230 -35 7600 -25
rect 7230 -95 7234 -35
rect 7286 -95 7544 -35
rect 7596 -95 7600 -35
rect 7230 -164 7600 -95
rect 7630 -35 8000 -25
rect 7630 -95 7634 -35
rect 7686 -95 7944 -35
rect 7996 -95 8000 -35
rect 7630 -164 8000 -95
rect 8030 -35 8400 -25
rect 8030 -95 8034 -35
rect 8086 -95 8344 -35
rect 8396 -95 8400 -35
rect 8030 -164 8400 -95
rect 8430 -35 8800 -25
rect 8430 -95 8434 -35
rect 8486 -95 8744 -35
rect 8796 -95 8800 -35
rect 8430 -164 8800 -95
rect 8830 -35 9200 -25
rect 8830 -95 8834 -35
rect 8886 -95 9144 -35
rect 9196 -95 9200 -35
rect 8830 -164 9200 -95
rect 9230 -35 9600 -25
rect 9230 -95 9234 -35
rect 9286 -95 9544 -35
rect 9596 -95 9600 -35
rect 9230 -164 9600 -95
rect 9630 -35 10000 -25
rect 9630 -95 9634 -35
rect 9686 -95 9944 -35
rect 9996 -95 10000 -35
rect 9630 -164 10000 -95
rect 10030 -35 10400 -25
rect 10030 -95 10034 -35
rect 10086 -95 10344 -35
rect 10396 -95 10400 -35
rect 10030 -164 10400 -95
rect 10430 -35 10800 -25
rect 10430 -95 10434 -35
rect 10486 -95 10744 -35
rect 10796 -95 10800 -35
rect 10430 -164 10800 -95
rect 10830 -35 11200 -25
rect 10830 -95 10834 -35
rect 10886 -95 11144 -35
rect 11196 -95 11200 -35
rect 10830 -164 11200 -95
rect 11230 -35 11600 -25
rect 11230 -95 11234 -35
rect 11286 -95 11544 -35
rect 11596 -95 11600 -35
rect 11230 -164 11600 -95
rect 11630 -35 12000 -25
rect 11630 -95 11634 -35
rect 11686 -95 11944 -35
rect 11996 -95 12000 -35
rect 11630 -164 12000 -95
rect 12030 -35 12400 -25
rect 12030 -95 12034 -35
rect 12086 -95 12344 -35
rect 12396 -95 12400 -35
rect 12030 -164 12400 -95
rect 12430 -35 12800 -25
rect 12430 -95 12434 -35
rect 12486 -95 12744 -35
rect 12796 -95 12800 -35
rect 12430 -164 12800 -95
rect 12830 -35 13200 -25
rect 12830 -95 12834 -35
rect 12886 -95 13144 -35
rect 13196 -95 13200 -35
rect 12830 -164 13200 -95
rect -370 -170 13200 -164
rect -370 -210 -220 -170
rect 12960 -210 13200 -170
rect -370 -216 13200 -210
rect -370 -295 0 -216
rect -370 -355 -366 -295
rect -314 -355 -56 -295
rect -4 -355 0 -295
rect -370 -365 0 -355
rect 30 -295 400 -216
rect 30 -355 34 -295
rect 86 -355 344 -295
rect 396 -355 400 -295
rect 30 -365 400 -355
rect 430 -295 800 -216
rect 430 -355 434 -295
rect 486 -355 744 -295
rect 796 -355 800 -295
rect 430 -365 800 -355
rect 830 -295 1200 -216
rect 830 -355 834 -295
rect 886 -355 1144 -295
rect 1196 -355 1200 -295
rect 830 -365 1200 -355
rect 1230 -295 1600 -216
rect 1230 -355 1234 -295
rect 1286 -355 1544 -295
rect 1596 -355 1600 -295
rect 1230 -365 1600 -355
rect 1630 -295 2000 -216
rect 1630 -355 1634 -295
rect 1686 -355 1944 -295
rect 1996 -355 2000 -295
rect 1630 -365 2000 -355
rect 2030 -295 2400 -216
rect 2030 -355 2034 -295
rect 2086 -355 2344 -295
rect 2396 -355 2400 -295
rect 2030 -365 2400 -355
rect 2430 -295 2800 -216
rect 2430 -355 2434 -295
rect 2486 -355 2744 -295
rect 2796 -355 2800 -295
rect 2430 -365 2800 -355
rect 2830 -295 3200 -216
rect 2830 -355 2834 -295
rect 2886 -355 3144 -295
rect 3196 -355 3200 -295
rect 2830 -365 3200 -355
rect 3230 -295 3600 -216
rect 3230 -355 3234 -295
rect 3286 -355 3544 -295
rect 3596 -355 3600 -295
rect 3230 -365 3600 -355
rect 3630 -295 4000 -216
rect 3630 -355 3634 -295
rect 3686 -355 3944 -295
rect 3996 -355 4000 -295
rect 3630 -365 4000 -355
rect 4030 -295 4400 -216
rect 4030 -355 4034 -295
rect 4086 -355 4344 -295
rect 4396 -355 4400 -295
rect 4030 -365 4400 -355
rect 4430 -295 4800 -216
rect 4430 -355 4434 -295
rect 4486 -355 4744 -295
rect 4796 -355 4800 -295
rect 4430 -365 4800 -355
rect 4830 -295 5200 -216
rect 4830 -355 4834 -295
rect 4886 -355 5144 -295
rect 5196 -355 5200 -295
rect 4830 -365 5200 -355
rect 5230 -295 5600 -216
rect 5230 -355 5234 -295
rect 5286 -355 5544 -295
rect 5596 -355 5600 -295
rect 5230 -365 5600 -355
rect 5630 -295 6000 -216
rect 5630 -355 5634 -295
rect 5686 -355 5944 -295
rect 5996 -355 6000 -295
rect 5630 -365 6000 -355
rect 6030 -295 6400 -216
rect 6030 -355 6034 -295
rect 6086 -355 6344 -295
rect 6396 -355 6400 -295
rect 6030 -365 6400 -355
rect 6430 -295 6800 -216
rect 6430 -355 6434 -295
rect 6486 -355 6744 -295
rect 6796 -355 6800 -295
rect 6430 -365 6800 -355
rect 6830 -295 7200 -216
rect 6830 -355 6834 -295
rect 6886 -355 7144 -295
rect 7196 -355 7200 -295
rect 6830 -365 7200 -355
rect 7230 -295 7600 -216
rect 7230 -355 7234 -295
rect 7286 -355 7544 -295
rect 7596 -355 7600 -295
rect 7230 -365 7600 -355
rect 7630 -295 8000 -216
rect 7630 -355 7634 -295
rect 7686 -355 7944 -295
rect 7996 -355 8000 -295
rect 7630 -365 8000 -355
rect 8030 -295 8400 -216
rect 8030 -355 8034 -295
rect 8086 -355 8344 -295
rect 8396 -355 8400 -295
rect 8030 -365 8400 -355
rect 8430 -295 8800 -216
rect 8430 -355 8434 -295
rect 8486 -355 8744 -295
rect 8796 -355 8800 -295
rect 8430 -365 8800 -355
rect 8830 -295 9200 -216
rect 8830 -355 8834 -295
rect 8886 -355 9144 -295
rect 9196 -355 9200 -295
rect 8830 -365 9200 -355
rect 9230 -295 9600 -216
rect 9230 -355 9234 -295
rect 9286 -355 9544 -295
rect 9596 -355 9600 -295
rect 9230 -365 9600 -355
rect 9630 -295 10000 -216
rect 9630 -355 9634 -295
rect 9686 -355 9944 -295
rect 9996 -355 10000 -295
rect 9630 -365 10000 -355
rect 10030 -295 10400 -216
rect 10030 -355 10034 -295
rect 10086 -355 10344 -295
rect 10396 -355 10400 -295
rect 10030 -365 10400 -355
rect 10430 -295 10800 -216
rect 10430 -355 10434 -295
rect 10486 -355 10744 -295
rect 10796 -355 10800 -295
rect 10430 -365 10800 -355
rect 10830 -295 11200 -216
rect 10830 -355 10834 -295
rect 10886 -355 11144 -295
rect 11196 -355 11200 -295
rect 10830 -365 11200 -355
rect 11230 -295 11600 -216
rect 11230 -355 11234 -295
rect 11286 -355 11544 -295
rect 11596 -355 11600 -295
rect 11230 -365 11600 -355
rect 11630 -295 12000 -216
rect 11630 -355 11634 -295
rect 11686 -355 11944 -295
rect 11996 -355 12000 -295
rect 11630 -365 12000 -355
rect 12030 -295 12400 -216
rect 12030 -355 12034 -295
rect 12086 -355 12344 -295
rect 12396 -355 12400 -295
rect 12030 -365 12400 -355
rect 12430 -295 12800 -216
rect 12430 -355 12434 -295
rect 12486 -355 12744 -295
rect 12796 -355 12800 -295
rect 12430 -365 12800 -355
rect 12830 -295 13200 -216
rect 12830 -355 12834 -295
rect 12886 -355 13144 -295
rect 13196 -355 13200 -295
rect 12830 -365 13200 -355
<< via1 >>
rect -265 24170 -205 24180
rect -265 24130 -255 24170
rect -255 24130 -215 24170
rect -215 24130 -205 24170
rect -265 24120 -205 24130
rect -165 24170 -105 24180
rect -165 24130 -155 24170
rect -155 24130 -115 24170
rect -115 24130 -105 24170
rect -165 24120 -105 24130
rect 12930 24115 12990 24125
rect 12930 24075 12940 24115
rect 12940 24075 12980 24115
rect 12980 24075 12990 24115
rect 12930 24065 12990 24075
rect 13030 24115 13090 24125
rect 13030 24075 13040 24115
rect 13040 24075 13080 24115
rect 13080 24075 13090 24115
rect 13030 24065 13090 24075
rect -366 23955 -314 24015
rect -56 23955 -4 24015
rect 34 23955 86 24015
rect 344 23955 396 24015
rect 434 23955 486 24015
rect 744 23955 796 24015
rect 834 23955 886 24015
rect 1144 23955 1196 24015
rect 1234 23955 1286 24015
rect 1544 23955 1596 24015
rect 1634 23955 1686 24015
rect 1944 23955 1996 24015
rect 2034 23955 2086 24015
rect 2344 23955 2396 24015
rect 2434 23955 2486 24015
rect 2744 23955 2796 24015
rect 2834 23955 2886 24015
rect 3144 23955 3196 24015
rect 3234 23955 3286 24015
rect 3544 23955 3596 24015
rect 3634 23955 3686 24015
rect 3944 23955 3996 24015
rect 4034 23955 4086 24015
rect 4344 23955 4396 24015
rect 4434 23955 4486 24015
rect 4744 23955 4796 24015
rect 4834 23955 4886 24015
rect 5144 23955 5196 24015
rect 5234 23955 5286 24015
rect 5544 23955 5596 24015
rect 5634 23955 5686 24015
rect 5944 23955 5996 24015
rect 6034 23955 6086 24015
rect 6344 23955 6396 24015
rect 6434 23955 6486 24015
rect 6744 23955 6796 24015
rect 6834 23955 6886 24015
rect 7144 23955 7196 24015
rect 7234 23955 7286 24015
rect 7544 23955 7596 24015
rect 7634 23955 7686 24015
rect 7944 23955 7996 24015
rect 8034 23955 8086 24015
rect 8344 23955 8396 24015
rect 8434 23955 8486 24015
rect 8744 23955 8796 24015
rect 8834 23955 8886 24015
rect 9144 23955 9196 24015
rect 9234 23955 9286 24015
rect 9544 23955 9596 24015
rect 9634 23955 9686 24015
rect 9944 23955 9996 24015
rect 10034 23955 10086 24015
rect 10344 23955 10396 24015
rect 10434 23955 10486 24015
rect 10744 23955 10796 24015
rect 10834 23955 10886 24015
rect 11144 23955 11196 24015
rect 11234 23955 11286 24015
rect 11544 23955 11596 24015
rect 11634 23955 11686 24015
rect 11944 23955 11996 24015
rect 12034 23955 12086 24015
rect 12344 23955 12396 24015
rect 12434 23955 12486 24015
rect 12744 23955 12796 24015
rect 12834 23955 12886 24015
rect 13144 23955 13196 24015
rect -366 23740 -314 23755
rect -366 23695 -330 23740
rect -330 23695 -314 23740
rect -56 23695 -4 23755
rect 34 23695 86 23755
rect 344 23695 396 23755
rect 434 23695 486 23755
rect 744 23695 796 23755
rect 834 23695 886 23755
rect 1144 23695 1196 23755
rect 1234 23695 1286 23755
rect 1544 23695 1596 23755
rect 1634 23695 1686 23755
rect 1944 23695 1996 23755
rect 2034 23695 2086 23755
rect 2344 23695 2396 23755
rect 2434 23695 2486 23755
rect 2744 23695 2796 23755
rect 2834 23695 2886 23755
rect 3144 23695 3196 23755
rect 3234 23695 3286 23755
rect 3544 23695 3596 23755
rect 3634 23695 3686 23755
rect 3944 23695 3996 23755
rect 4034 23695 4086 23755
rect 4344 23695 4396 23755
rect 4434 23695 4486 23755
rect 4744 23695 4796 23755
rect 4834 23695 4886 23755
rect 5144 23695 5196 23755
rect 5234 23695 5286 23755
rect 5544 23695 5596 23755
rect 5634 23695 5686 23755
rect 5944 23695 5996 23755
rect 6034 23695 6086 23755
rect 6344 23695 6396 23755
rect 6434 23695 6486 23755
rect 6744 23695 6796 23755
rect 6834 23695 6886 23755
rect 7144 23695 7196 23755
rect 7234 23695 7286 23755
rect 7544 23695 7596 23755
rect 7634 23695 7686 23755
rect 7944 23695 7996 23755
rect 8034 23695 8086 23755
rect 8344 23695 8396 23755
rect 8434 23695 8486 23755
rect 8744 23695 8796 23755
rect 8834 23695 8886 23755
rect 9144 23695 9196 23755
rect 9234 23695 9286 23755
rect 9544 23695 9596 23755
rect 9634 23695 9686 23755
rect 9944 23695 9996 23755
rect 10034 23695 10086 23755
rect 10344 23695 10396 23755
rect 10434 23695 10486 23755
rect 10744 23695 10796 23755
rect 10834 23695 10886 23755
rect 11144 23695 11196 23755
rect 11234 23695 11286 23755
rect 11544 23695 11596 23755
rect 11634 23695 11686 23755
rect 11944 23695 11996 23755
rect 12034 23695 12086 23755
rect 12344 23695 12396 23755
rect 12434 23695 12486 23755
rect 12744 23695 12796 23755
rect 12834 23695 12886 23755
rect 13144 23695 13196 23755
rect -366 23585 -330 23645
rect -330 23585 -314 23645
rect -56 23585 -4 23645
rect -366 23325 -330 23385
rect -330 23325 -314 23385
rect -56 23325 -4 23385
rect 34 23585 86 23645
rect 344 23585 396 23645
rect 434 23585 486 23645
rect 744 23585 796 23645
rect 834 23585 886 23645
rect 1144 23585 1196 23645
rect 1234 23585 1286 23645
rect 1544 23585 1596 23645
rect 1634 23585 1686 23645
rect 1944 23585 1996 23645
rect 2034 23585 2086 23645
rect 2344 23585 2396 23645
rect 2434 23585 2486 23645
rect 2744 23585 2796 23645
rect 2834 23585 2886 23645
rect 3144 23585 3196 23645
rect 3234 23585 3286 23645
rect 3544 23585 3596 23645
rect 3634 23585 3686 23645
rect 3944 23585 3996 23645
rect 4034 23585 4086 23645
rect 4344 23585 4396 23645
rect 4434 23585 4486 23645
rect 4744 23585 4796 23645
rect 4834 23585 4886 23645
rect 5144 23585 5196 23645
rect 5234 23585 5286 23645
rect 5544 23585 5596 23645
rect 5634 23585 5686 23645
rect 5944 23585 5996 23645
rect 6034 23585 6086 23645
rect 6344 23585 6396 23645
rect 6434 23585 6486 23645
rect 6744 23585 6796 23645
rect 6834 23585 6886 23645
rect 7144 23585 7196 23645
rect 7234 23585 7286 23645
rect 7544 23585 7596 23645
rect 7634 23585 7686 23645
rect 7944 23585 7996 23645
rect 8034 23585 8086 23645
rect 8344 23585 8396 23645
rect 8434 23585 8486 23645
rect 8744 23585 8796 23645
rect 8834 23585 8886 23645
rect 9144 23585 9196 23645
rect 9234 23585 9286 23645
rect 9544 23585 9596 23645
rect 9634 23585 9686 23645
rect 9944 23585 9996 23645
rect 10034 23585 10086 23645
rect 10344 23585 10396 23645
rect 10434 23585 10486 23645
rect 10744 23585 10796 23645
rect 10834 23585 10886 23645
rect 11144 23585 11196 23645
rect 11234 23585 11286 23645
rect 11544 23585 11596 23645
rect 11634 23585 11686 23645
rect 11944 23585 11996 23645
rect 12034 23585 12086 23645
rect 12344 23585 12396 23645
rect 12434 23585 12486 23645
rect 12744 23585 12796 23645
rect 12834 23585 12886 23645
rect 13144 23585 13196 23645
rect 34 23325 86 23385
rect 344 23325 396 23385
rect 434 23325 486 23385
rect 744 23325 796 23385
rect 834 23325 886 23385
rect 1144 23325 1196 23385
rect 1234 23325 1286 23385
rect 1544 23325 1596 23385
rect 1634 23325 1686 23385
rect 1944 23325 1996 23385
rect 2034 23325 2086 23385
rect 2344 23325 2396 23385
rect 2434 23325 2486 23385
rect 2744 23325 2796 23385
rect 2834 23325 2886 23385
rect 3144 23325 3196 23385
rect 3234 23325 3286 23385
rect 3544 23325 3596 23385
rect 3634 23325 3686 23385
rect 3944 23325 3996 23385
rect 4034 23325 4086 23385
rect 4344 23325 4396 23385
rect 4434 23325 4486 23385
rect 4744 23325 4796 23385
rect 4834 23325 4886 23385
rect 5144 23325 5196 23385
rect 5234 23325 5286 23385
rect 5544 23325 5596 23385
rect 5634 23325 5686 23385
rect 5944 23325 5996 23385
rect 6034 23325 6086 23385
rect 6344 23325 6396 23385
rect 6434 23325 6486 23385
rect 6744 23325 6796 23385
rect 6834 23325 6886 23385
rect 7144 23325 7196 23385
rect 7234 23325 7286 23385
rect 7544 23325 7596 23385
rect 7634 23325 7686 23385
rect 7944 23325 7996 23385
rect 8034 23325 8086 23385
rect 8344 23325 8396 23385
rect 8434 23325 8486 23385
rect 8744 23325 8796 23385
rect 8834 23325 8886 23385
rect 9144 23325 9196 23385
rect 9234 23325 9286 23385
rect 9544 23325 9596 23385
rect 9634 23325 9686 23385
rect 9944 23325 9996 23385
rect 10034 23325 10086 23385
rect 10344 23325 10396 23385
rect 10434 23325 10486 23385
rect 10744 23325 10796 23385
rect 10834 23325 10886 23385
rect 11144 23325 11196 23385
rect 11234 23325 11286 23385
rect 11544 23325 11596 23385
rect 11634 23325 11686 23385
rect 11944 23325 11996 23385
rect 12034 23325 12086 23385
rect 12344 23325 12396 23385
rect 12434 23325 12486 23385
rect 12744 23325 12796 23385
rect 12834 23325 12886 23385
rect 13144 23325 13196 23385
rect -366 23215 -330 23275
rect -330 23215 -314 23275
rect -56 23215 -4 23275
rect -366 22955 -330 23015
rect -330 22955 -314 23015
rect -56 22955 -4 23015
rect 34 23215 86 23275
rect 344 23215 396 23275
rect 434 23215 486 23275
rect 744 23215 796 23275
rect 834 23215 886 23275
rect 1144 23215 1196 23275
rect 1234 23215 1286 23275
rect 1544 23215 1596 23275
rect 1634 23215 1686 23275
rect 1944 23215 1996 23275
rect 2034 23215 2086 23275
rect 2344 23215 2396 23275
rect 2434 23215 2486 23275
rect 2744 23215 2796 23275
rect 2834 23215 2886 23275
rect 3144 23215 3196 23275
rect 3234 23215 3286 23275
rect 3544 23215 3596 23275
rect 3634 23215 3686 23275
rect 3944 23215 3996 23275
rect 4034 23215 4086 23275
rect 4344 23215 4396 23275
rect 4434 23215 4486 23275
rect 4744 23215 4796 23275
rect 4834 23215 4886 23275
rect 5144 23215 5196 23275
rect 5234 23215 5286 23275
rect 5544 23215 5596 23275
rect 5634 23215 5686 23275
rect 5944 23215 5996 23275
rect 6034 23215 6086 23275
rect 6344 23215 6396 23275
rect 6434 23215 6486 23275
rect 6744 23215 6796 23275
rect 6834 23215 6886 23275
rect 7144 23215 7196 23275
rect 7234 23215 7286 23275
rect 7544 23215 7596 23275
rect 7634 23215 7686 23275
rect 7944 23215 7996 23275
rect 8034 23215 8086 23275
rect 8344 23215 8396 23275
rect 8434 23215 8486 23275
rect 8744 23215 8796 23275
rect 8834 23215 8886 23275
rect 9144 23215 9196 23275
rect 9234 23215 9286 23275
rect 9544 23215 9596 23275
rect 9634 23215 9686 23275
rect 9944 23215 9996 23275
rect 10034 23215 10086 23275
rect 10344 23215 10396 23275
rect 10434 23215 10486 23275
rect 10744 23215 10796 23275
rect 10834 23215 10886 23275
rect 11144 23215 11196 23275
rect 11234 23215 11286 23275
rect 11544 23215 11596 23275
rect 11634 23215 11686 23275
rect 11944 23215 11996 23275
rect 12034 23215 12086 23275
rect 12344 23215 12396 23275
rect 12434 23215 12486 23275
rect 12744 23215 12796 23275
rect 12834 23215 12886 23275
rect 13144 23215 13196 23275
rect 34 22955 86 23015
rect 344 22955 396 23015
rect 434 22955 486 23015
rect 744 22955 796 23015
rect 834 22955 886 23015
rect 1144 22955 1196 23015
rect 1234 22955 1286 23015
rect 1544 22955 1596 23015
rect 1634 22955 1686 23015
rect 1944 22955 1996 23015
rect 2034 22955 2086 23015
rect 2344 22955 2396 23015
rect 2434 22955 2486 23015
rect 2744 22955 2796 23015
rect 2834 22955 2886 23015
rect 3144 22955 3196 23015
rect 3234 22955 3286 23015
rect 3544 22955 3596 23015
rect 3634 22955 3686 23015
rect 3944 22955 3996 23015
rect 4034 22955 4086 23015
rect 4344 22955 4396 23015
rect 4434 22955 4486 23015
rect 4744 22955 4796 23015
rect 4834 22955 4886 23015
rect 5144 22955 5196 23015
rect 5234 22955 5286 23015
rect 5544 22955 5596 23015
rect 5634 22955 5686 23015
rect 5944 22955 5996 23015
rect 6034 22955 6086 23015
rect 6344 22955 6396 23015
rect 6434 22955 6486 23015
rect 6744 22955 6796 23015
rect 6834 22955 6886 23015
rect 7144 22955 7196 23015
rect 7234 22955 7286 23015
rect 7544 22955 7596 23015
rect 7634 22955 7686 23015
rect 7944 22955 7996 23015
rect 8034 22955 8086 23015
rect 8344 22955 8396 23015
rect 8434 22955 8486 23015
rect 8744 22955 8796 23015
rect 8834 22955 8886 23015
rect 9144 22955 9196 23015
rect 9234 22955 9286 23015
rect 9544 22955 9596 23015
rect 9634 22955 9686 23015
rect 9944 22955 9996 23015
rect 10034 22955 10086 23015
rect 10344 22955 10396 23015
rect 10434 22955 10486 23015
rect 10744 22955 10796 23015
rect 10834 22955 10886 23015
rect 11144 22955 11196 23015
rect 11234 22955 11286 23015
rect 11544 22955 11596 23015
rect 11634 22955 11686 23015
rect 11944 22955 11996 23015
rect 12034 22955 12086 23015
rect 12344 22955 12396 23015
rect 12434 22955 12486 23015
rect 12744 22955 12796 23015
rect 12834 22955 12886 23015
rect 13144 22955 13196 23015
rect -366 22845 -330 22905
rect -330 22845 -314 22905
rect -56 22845 -4 22905
rect -366 22585 -330 22645
rect -330 22585 -314 22645
rect -56 22585 -4 22645
rect 34 22845 86 22905
rect 344 22845 396 22905
rect 434 22845 486 22905
rect 744 22845 796 22905
rect 834 22845 886 22905
rect 1144 22845 1196 22905
rect 1234 22845 1286 22905
rect 1544 22845 1596 22905
rect 1634 22845 1686 22905
rect 1944 22845 1996 22905
rect 2034 22845 2086 22905
rect 2344 22845 2396 22905
rect 2434 22845 2486 22905
rect 2744 22845 2796 22905
rect 2834 22845 2886 22905
rect 3144 22845 3196 22905
rect 3234 22845 3286 22905
rect 3544 22845 3596 22905
rect 3634 22845 3686 22905
rect 3944 22845 3996 22905
rect 4034 22845 4086 22905
rect 4344 22845 4396 22905
rect 4434 22845 4486 22905
rect 4744 22845 4796 22905
rect 4834 22845 4886 22905
rect 5144 22845 5196 22905
rect 5234 22845 5286 22905
rect 5544 22845 5596 22905
rect 5634 22845 5686 22905
rect 5944 22845 5996 22905
rect 6034 22845 6086 22905
rect 6344 22845 6396 22905
rect 6434 22845 6486 22905
rect 6744 22845 6796 22905
rect 6834 22845 6886 22905
rect 7144 22845 7196 22905
rect 7234 22845 7286 22905
rect 7544 22845 7596 22905
rect 7634 22845 7686 22905
rect 7944 22845 7996 22905
rect 8034 22845 8086 22905
rect 8344 22845 8396 22905
rect 8434 22845 8486 22905
rect 8744 22845 8796 22905
rect 8834 22845 8886 22905
rect 9144 22845 9196 22905
rect 9234 22845 9286 22905
rect 9544 22845 9596 22905
rect 9634 22845 9686 22905
rect 9944 22845 9996 22905
rect 10034 22845 10086 22905
rect 10344 22845 10396 22905
rect 10434 22845 10486 22905
rect 10744 22845 10796 22905
rect 10834 22845 10886 22905
rect 11144 22845 11196 22905
rect 11234 22845 11286 22905
rect 11544 22845 11596 22905
rect 11634 22845 11686 22905
rect 11944 22845 11996 22905
rect 12034 22845 12086 22905
rect 12344 22845 12396 22905
rect 12434 22845 12486 22905
rect 12744 22845 12796 22905
rect 12834 22845 12886 22905
rect 13144 22845 13196 22905
rect 34 22585 86 22645
rect 344 22585 396 22645
rect 434 22585 486 22645
rect 744 22585 796 22645
rect 834 22585 886 22645
rect 1144 22585 1196 22645
rect 1234 22585 1286 22645
rect 1544 22585 1596 22645
rect 1634 22585 1686 22645
rect 1944 22585 1996 22645
rect 2034 22585 2086 22645
rect 2344 22585 2396 22645
rect 2434 22585 2486 22645
rect 2744 22585 2796 22645
rect 2834 22585 2886 22645
rect 3144 22585 3196 22645
rect 3234 22585 3286 22645
rect 3544 22585 3596 22645
rect 3634 22585 3686 22645
rect 3944 22585 3996 22645
rect 4034 22585 4086 22645
rect 4344 22585 4396 22645
rect 4434 22585 4486 22645
rect 4744 22585 4796 22645
rect 4834 22585 4886 22645
rect 5144 22585 5196 22645
rect 5234 22585 5286 22645
rect 5544 22585 5596 22645
rect 5634 22585 5686 22645
rect 5944 22585 5996 22645
rect 6034 22585 6086 22645
rect 6344 22585 6396 22645
rect 6434 22585 6486 22645
rect 6744 22585 6796 22645
rect 6834 22585 6886 22645
rect 7144 22585 7196 22645
rect 7234 22585 7286 22645
rect 7544 22585 7596 22645
rect 7634 22585 7686 22645
rect 7944 22585 7996 22645
rect 8034 22585 8086 22645
rect 8344 22585 8396 22645
rect 8434 22585 8486 22645
rect 8744 22585 8796 22645
rect 8834 22585 8886 22645
rect 9144 22585 9196 22645
rect 9234 22585 9286 22645
rect 9544 22585 9596 22645
rect 9634 22585 9686 22645
rect 9944 22585 9996 22645
rect 10034 22585 10086 22645
rect 10344 22585 10396 22645
rect 10434 22585 10486 22645
rect 10744 22585 10796 22645
rect 10834 22585 10886 22645
rect 11144 22585 11196 22645
rect 11234 22585 11286 22645
rect 11544 22585 11596 22645
rect 11634 22585 11686 22645
rect 11944 22585 11996 22645
rect 12034 22585 12086 22645
rect 12344 22585 12396 22645
rect 12434 22585 12486 22645
rect 12744 22585 12796 22645
rect 12834 22585 12886 22645
rect 13144 22585 13196 22645
rect -366 22475 -330 22535
rect -330 22475 -314 22535
rect -56 22475 -4 22535
rect -366 22215 -330 22275
rect -330 22215 -314 22275
rect -56 22215 -4 22275
rect 34 22475 86 22535
rect 344 22475 396 22535
rect 434 22475 486 22535
rect 744 22475 796 22535
rect 834 22475 886 22535
rect 1144 22475 1196 22535
rect 1234 22475 1286 22535
rect 1544 22475 1596 22535
rect 1634 22475 1686 22535
rect 1944 22475 1996 22535
rect 2034 22475 2086 22535
rect 2344 22475 2396 22535
rect 2434 22475 2486 22535
rect 2744 22475 2796 22535
rect 2834 22475 2886 22535
rect 3144 22475 3196 22535
rect 3234 22475 3286 22535
rect 3544 22475 3596 22535
rect 3634 22475 3686 22535
rect 3944 22475 3996 22535
rect 4034 22475 4086 22535
rect 4344 22475 4396 22535
rect 4434 22475 4486 22535
rect 4744 22475 4796 22535
rect 4834 22475 4886 22535
rect 5144 22475 5196 22535
rect 5234 22475 5286 22535
rect 5544 22475 5596 22535
rect 5634 22475 5686 22535
rect 5944 22475 5996 22535
rect 6034 22475 6086 22535
rect 6344 22475 6396 22535
rect 6434 22475 6486 22535
rect 6744 22475 6796 22535
rect 6834 22475 6886 22535
rect 7144 22475 7196 22535
rect 7234 22475 7286 22535
rect 7544 22475 7596 22535
rect 7634 22475 7686 22535
rect 7944 22475 7996 22535
rect 8034 22475 8086 22535
rect 8344 22475 8396 22535
rect 8434 22475 8486 22535
rect 8744 22475 8796 22535
rect 8834 22475 8886 22535
rect 9144 22475 9196 22535
rect 9234 22475 9286 22535
rect 9544 22475 9596 22535
rect 9634 22475 9686 22535
rect 9944 22475 9996 22535
rect 10034 22475 10086 22535
rect 10344 22475 10396 22535
rect 10434 22475 10486 22535
rect 10744 22475 10796 22535
rect 10834 22475 10886 22535
rect 11144 22475 11196 22535
rect 11234 22475 11286 22535
rect 11544 22475 11596 22535
rect 11634 22475 11686 22535
rect 11944 22475 11996 22535
rect 12034 22475 12086 22535
rect 12344 22475 12396 22535
rect 12434 22475 12486 22535
rect 12744 22475 12796 22535
rect 12834 22475 12886 22535
rect 13144 22475 13196 22535
rect 34 22215 86 22275
rect 344 22215 396 22275
rect 434 22215 486 22275
rect 744 22215 796 22275
rect 834 22215 886 22275
rect 1144 22215 1196 22275
rect 1234 22215 1286 22275
rect 1544 22215 1596 22275
rect 1634 22215 1686 22275
rect 1944 22215 1996 22275
rect 2034 22215 2086 22275
rect 2344 22215 2396 22275
rect 2434 22215 2486 22275
rect 2744 22215 2796 22275
rect 2834 22215 2886 22275
rect 3144 22215 3196 22275
rect 3234 22215 3286 22275
rect 3544 22215 3596 22275
rect 3634 22215 3686 22275
rect 3944 22215 3996 22275
rect 4034 22215 4086 22275
rect 4344 22215 4396 22275
rect 4434 22215 4486 22275
rect 4744 22215 4796 22275
rect 4834 22215 4886 22275
rect 5144 22215 5196 22275
rect 5234 22215 5286 22275
rect 5544 22215 5596 22275
rect 5634 22215 5686 22275
rect 5944 22215 5996 22275
rect 6034 22215 6086 22275
rect 6344 22215 6396 22275
rect 6434 22215 6486 22275
rect 6744 22215 6796 22275
rect 6834 22215 6886 22275
rect 7144 22215 7196 22275
rect 7234 22215 7286 22275
rect 7544 22215 7596 22275
rect 7634 22215 7686 22275
rect 7944 22215 7996 22275
rect 8034 22215 8086 22275
rect 8344 22215 8396 22275
rect 8434 22215 8486 22275
rect 8744 22215 8796 22275
rect 8834 22215 8886 22275
rect 9144 22215 9196 22275
rect 9234 22215 9286 22275
rect 9544 22215 9596 22275
rect 9634 22215 9686 22275
rect 9944 22215 9996 22275
rect 10034 22215 10086 22275
rect 10344 22215 10396 22275
rect 10434 22215 10486 22275
rect 10744 22215 10796 22275
rect 10834 22215 10886 22275
rect 11144 22215 11196 22275
rect 11234 22215 11286 22275
rect 11544 22215 11596 22275
rect 11634 22215 11686 22275
rect 11944 22215 11996 22275
rect 12034 22215 12086 22275
rect 12344 22215 12396 22275
rect 12434 22215 12486 22275
rect 12744 22215 12796 22275
rect 12834 22215 12886 22275
rect 13144 22215 13196 22275
rect -366 22105 -330 22165
rect -330 22105 -314 22165
rect -56 22105 -4 22165
rect -366 21845 -330 21905
rect -330 21845 -314 21905
rect -56 21845 -4 21905
rect 34 22105 86 22165
rect 344 22105 396 22165
rect 434 22105 486 22165
rect 744 22105 796 22165
rect 834 22105 886 22165
rect 1144 22105 1196 22165
rect 1234 22105 1286 22165
rect 1544 22105 1596 22165
rect 1634 22105 1686 22165
rect 1944 22105 1996 22165
rect 2034 22105 2086 22165
rect 2344 22105 2396 22165
rect 2434 22105 2486 22165
rect 2744 22105 2796 22165
rect 2834 22105 2886 22165
rect 3144 22105 3196 22165
rect 3234 22105 3286 22165
rect 3544 22105 3596 22165
rect 3634 22105 3686 22165
rect 3944 22105 3996 22165
rect 4034 22105 4086 22165
rect 4344 22105 4396 22165
rect 4434 22105 4486 22165
rect 4744 22105 4796 22165
rect 4834 22105 4886 22165
rect 5144 22105 5196 22165
rect 5234 22105 5286 22165
rect 5544 22105 5596 22165
rect 5634 22105 5686 22165
rect 5944 22105 5996 22165
rect 6034 22105 6086 22165
rect 6344 22105 6396 22165
rect 6434 22105 6486 22165
rect 6744 22105 6796 22165
rect 6834 22105 6886 22165
rect 7144 22105 7196 22165
rect 7234 22105 7286 22165
rect 7544 22105 7596 22165
rect 7634 22105 7686 22165
rect 7944 22105 7996 22165
rect 8034 22105 8086 22165
rect 8344 22105 8396 22165
rect 8434 22105 8486 22165
rect 8744 22105 8796 22165
rect 8834 22105 8886 22165
rect 9144 22105 9196 22165
rect 9234 22105 9286 22165
rect 9544 22105 9596 22165
rect 9634 22105 9686 22165
rect 9944 22105 9996 22165
rect 10034 22105 10086 22165
rect 10344 22105 10396 22165
rect 10434 22105 10486 22165
rect 10744 22105 10796 22165
rect 10834 22105 10886 22165
rect 11144 22105 11196 22165
rect 11234 22105 11286 22165
rect 11544 22105 11596 22165
rect 11634 22105 11686 22165
rect 11944 22105 11996 22165
rect 12034 22105 12086 22165
rect 12344 22105 12396 22165
rect 12434 22105 12486 22165
rect 12744 22105 12796 22165
rect 12834 22105 12886 22165
rect 13144 22105 13196 22165
rect 34 21845 86 21905
rect 344 21845 396 21905
rect 434 21845 486 21905
rect 744 21845 796 21905
rect 834 21845 886 21905
rect 1144 21845 1196 21905
rect 1234 21845 1286 21905
rect 1544 21845 1596 21905
rect 1634 21845 1686 21905
rect 1944 21845 1996 21905
rect 2034 21845 2086 21905
rect 2344 21845 2396 21905
rect 2434 21845 2486 21905
rect 2744 21845 2796 21905
rect 2834 21845 2886 21905
rect 3144 21845 3196 21905
rect 3234 21845 3286 21905
rect 3544 21845 3596 21905
rect 3634 21845 3686 21905
rect 3944 21845 3996 21905
rect 4034 21845 4086 21905
rect 4344 21845 4396 21905
rect 4434 21845 4486 21905
rect 4744 21845 4796 21905
rect 4834 21845 4886 21905
rect 5144 21845 5196 21905
rect 5234 21845 5286 21905
rect 5544 21845 5596 21905
rect 5634 21845 5686 21905
rect 5944 21845 5996 21905
rect 6034 21845 6086 21905
rect 6344 21845 6396 21905
rect 6434 21845 6486 21905
rect 6744 21845 6796 21905
rect 6834 21845 6886 21905
rect 7144 21845 7196 21905
rect 7234 21845 7286 21905
rect 7544 21845 7596 21905
rect 7634 21845 7686 21905
rect 7944 21845 7996 21905
rect 8034 21845 8086 21905
rect 8344 21845 8396 21905
rect 8434 21845 8486 21905
rect 8744 21845 8796 21905
rect 8834 21845 8886 21905
rect 9144 21845 9196 21905
rect 9234 21845 9286 21905
rect 9544 21845 9596 21905
rect 9634 21845 9686 21905
rect 9944 21845 9996 21905
rect 10034 21845 10086 21905
rect 10344 21845 10396 21905
rect 10434 21845 10486 21905
rect 10744 21845 10796 21905
rect 10834 21845 10886 21905
rect 11144 21845 11196 21905
rect 11234 21845 11286 21905
rect 11544 21845 11596 21905
rect 11634 21845 11686 21905
rect 11944 21845 11996 21905
rect 12034 21845 12086 21905
rect 12344 21845 12396 21905
rect 12434 21845 12486 21905
rect 12744 21845 12796 21905
rect 12834 21845 12886 21905
rect 13144 21845 13196 21905
rect -366 21735 -330 21795
rect -330 21735 -314 21795
rect -56 21735 -4 21795
rect -366 21475 -330 21535
rect -330 21475 -314 21535
rect -56 21475 -4 21535
rect 34 21735 86 21795
rect 344 21735 396 21795
rect 434 21735 486 21795
rect 744 21735 796 21795
rect 834 21735 886 21795
rect 1144 21735 1196 21795
rect 1234 21735 1286 21795
rect 1544 21735 1596 21795
rect 1634 21735 1686 21795
rect 1944 21735 1996 21795
rect 2034 21735 2086 21795
rect 2344 21735 2396 21795
rect 2434 21735 2486 21795
rect 2744 21735 2796 21795
rect 2834 21735 2886 21795
rect 3144 21735 3196 21795
rect 3234 21735 3286 21795
rect 3544 21735 3596 21795
rect 3634 21735 3686 21795
rect 3944 21735 3996 21795
rect 4034 21735 4086 21795
rect 4344 21735 4396 21795
rect 4434 21735 4486 21795
rect 4744 21735 4796 21795
rect 4834 21735 4886 21795
rect 5144 21735 5196 21795
rect 5234 21735 5286 21795
rect 5544 21735 5596 21795
rect 5634 21735 5686 21795
rect 5944 21735 5996 21795
rect 6034 21735 6086 21795
rect 6344 21735 6396 21795
rect 6434 21735 6486 21795
rect 6744 21735 6796 21795
rect 6834 21735 6886 21795
rect 7144 21735 7196 21795
rect 7234 21735 7286 21795
rect 7544 21735 7596 21795
rect 7634 21735 7686 21795
rect 7944 21735 7996 21795
rect 8034 21735 8086 21795
rect 8344 21735 8396 21795
rect 8434 21735 8486 21795
rect 8744 21735 8796 21795
rect 8834 21735 8886 21795
rect 9144 21735 9196 21795
rect 9234 21735 9286 21795
rect 9544 21735 9596 21795
rect 9634 21735 9686 21795
rect 9944 21735 9996 21795
rect 10034 21735 10086 21795
rect 10344 21735 10396 21795
rect 10434 21735 10486 21795
rect 10744 21735 10796 21795
rect 10834 21735 10886 21795
rect 11144 21735 11196 21795
rect 11234 21735 11286 21795
rect 11544 21735 11596 21795
rect 11634 21735 11686 21795
rect 11944 21735 11996 21795
rect 12034 21735 12086 21795
rect 12344 21735 12396 21795
rect 12434 21735 12486 21795
rect 12744 21735 12796 21795
rect 12834 21735 12886 21795
rect 13144 21735 13196 21795
rect 34 21475 86 21535
rect 344 21475 396 21535
rect 434 21475 486 21535
rect 744 21475 796 21535
rect 834 21475 886 21535
rect 1144 21475 1196 21535
rect 1234 21475 1286 21535
rect 1544 21475 1596 21535
rect 1634 21475 1686 21535
rect 1944 21475 1996 21535
rect 2034 21475 2086 21535
rect 2344 21475 2396 21535
rect 2434 21475 2486 21535
rect 2744 21475 2796 21535
rect 2834 21475 2886 21535
rect 3144 21475 3196 21535
rect 3234 21475 3286 21535
rect 3544 21475 3596 21535
rect 3634 21475 3686 21535
rect 3944 21475 3996 21535
rect 4034 21475 4086 21535
rect 4344 21475 4396 21535
rect 4434 21475 4486 21535
rect 4744 21475 4796 21535
rect 4834 21475 4886 21535
rect 5144 21475 5196 21535
rect 5234 21475 5286 21535
rect 5544 21475 5596 21535
rect 5634 21475 5686 21535
rect 5944 21475 5996 21535
rect 6034 21475 6086 21535
rect 6344 21475 6396 21535
rect 6434 21475 6486 21535
rect 6744 21475 6796 21535
rect 6834 21475 6886 21535
rect 7144 21475 7196 21535
rect 7234 21475 7286 21535
rect 7544 21475 7596 21535
rect 7634 21475 7686 21535
rect 7944 21475 7996 21535
rect 8034 21475 8086 21535
rect 8344 21475 8396 21535
rect 8434 21475 8486 21535
rect 8744 21475 8796 21535
rect 8834 21475 8886 21535
rect 9144 21475 9196 21535
rect 9234 21475 9286 21535
rect 9544 21475 9596 21535
rect 9634 21475 9686 21535
rect 9944 21475 9996 21535
rect 10034 21475 10086 21535
rect 10344 21475 10396 21535
rect 10434 21475 10486 21535
rect 10744 21475 10796 21535
rect 10834 21475 10886 21535
rect 11144 21475 11196 21535
rect 11234 21475 11286 21535
rect 11544 21475 11596 21535
rect 11634 21475 11686 21535
rect 11944 21475 11996 21535
rect 12034 21475 12086 21535
rect 12344 21475 12396 21535
rect 12434 21475 12486 21535
rect 12744 21475 12796 21535
rect 12834 21475 12886 21535
rect 13144 21475 13196 21535
rect -366 21365 -330 21425
rect -330 21365 -314 21425
rect -56 21365 -4 21425
rect -366 21105 -330 21165
rect -330 21105 -314 21165
rect -56 21105 -4 21165
rect 34 21365 86 21425
rect 344 21365 396 21425
rect 434 21365 486 21425
rect 744 21365 796 21425
rect 834 21365 886 21425
rect 1144 21365 1196 21425
rect 1234 21365 1286 21425
rect 1544 21365 1596 21425
rect 1634 21365 1686 21425
rect 1944 21365 1996 21425
rect 2034 21365 2086 21425
rect 2344 21365 2396 21425
rect 2434 21365 2486 21425
rect 2744 21365 2796 21425
rect 2834 21365 2886 21425
rect 3144 21365 3196 21425
rect 3234 21365 3286 21425
rect 3544 21365 3596 21425
rect 3634 21365 3686 21425
rect 3944 21365 3996 21425
rect 4034 21365 4086 21425
rect 4344 21365 4396 21425
rect 4434 21365 4486 21425
rect 4744 21365 4796 21425
rect 4834 21365 4886 21425
rect 5144 21365 5196 21425
rect 5234 21365 5286 21425
rect 5544 21365 5596 21425
rect 5634 21365 5686 21425
rect 5944 21365 5996 21425
rect 6034 21365 6086 21425
rect 6344 21365 6396 21425
rect 6434 21365 6486 21425
rect 6744 21365 6796 21425
rect 6834 21365 6886 21425
rect 7144 21365 7196 21425
rect 7234 21365 7286 21425
rect 7544 21365 7596 21425
rect 7634 21365 7686 21425
rect 7944 21365 7996 21425
rect 8034 21365 8086 21425
rect 8344 21365 8396 21425
rect 8434 21365 8486 21425
rect 8744 21365 8796 21425
rect 8834 21365 8886 21425
rect 9144 21365 9196 21425
rect 9234 21365 9286 21425
rect 9544 21365 9596 21425
rect 9634 21365 9686 21425
rect 9944 21365 9996 21425
rect 10034 21365 10086 21425
rect 10344 21365 10396 21425
rect 10434 21365 10486 21425
rect 10744 21365 10796 21425
rect 10834 21365 10886 21425
rect 11144 21365 11196 21425
rect 11234 21365 11286 21425
rect 11544 21365 11596 21425
rect 11634 21365 11686 21425
rect 11944 21365 11996 21425
rect 12034 21365 12086 21425
rect 12344 21365 12396 21425
rect 12434 21365 12486 21425
rect 12744 21365 12796 21425
rect 12834 21365 12886 21425
rect 13144 21365 13196 21425
rect 34 21105 86 21165
rect 344 21105 396 21165
rect 434 21105 486 21165
rect 744 21105 796 21165
rect 834 21105 886 21165
rect 1144 21105 1196 21165
rect 1234 21105 1286 21165
rect 1544 21105 1596 21165
rect 1634 21105 1686 21165
rect 1944 21105 1996 21165
rect 2034 21105 2086 21165
rect 2344 21105 2396 21165
rect 2434 21105 2486 21165
rect 2744 21105 2796 21165
rect 2834 21105 2886 21165
rect 3144 21105 3196 21165
rect 3234 21105 3286 21165
rect 3544 21105 3596 21165
rect 3634 21105 3686 21165
rect 3944 21105 3996 21165
rect 4034 21105 4086 21165
rect 4344 21105 4396 21165
rect 4434 21105 4486 21165
rect 4744 21105 4796 21165
rect 4834 21105 4886 21165
rect 5144 21105 5196 21165
rect 5234 21105 5286 21165
rect 5544 21105 5596 21165
rect 5634 21105 5686 21165
rect 5944 21105 5996 21165
rect 6034 21105 6086 21165
rect 6344 21105 6396 21165
rect 6434 21105 6486 21165
rect 6744 21105 6796 21165
rect 6834 21105 6886 21165
rect 7144 21105 7196 21165
rect 7234 21105 7286 21165
rect 7544 21105 7596 21165
rect 7634 21105 7686 21165
rect 7944 21105 7996 21165
rect 8034 21105 8086 21165
rect 8344 21105 8396 21165
rect 8434 21105 8486 21165
rect 8744 21105 8796 21165
rect 8834 21105 8886 21165
rect 9144 21105 9196 21165
rect 9234 21105 9286 21165
rect 9544 21105 9596 21165
rect 9634 21105 9686 21165
rect 9944 21105 9996 21165
rect 10034 21105 10086 21165
rect 10344 21105 10396 21165
rect 10434 21105 10486 21165
rect 10744 21105 10796 21165
rect 10834 21105 10886 21165
rect 11144 21105 11196 21165
rect 11234 21105 11286 21165
rect 11544 21105 11596 21165
rect 11634 21105 11686 21165
rect 11944 21105 11996 21165
rect 12034 21105 12086 21165
rect 12344 21105 12396 21165
rect 12434 21105 12486 21165
rect 12744 21105 12796 21165
rect 12834 21105 12886 21165
rect 13144 21105 13196 21165
rect -366 20995 -330 21055
rect -330 20995 -314 21055
rect -56 20995 -4 21055
rect -366 20735 -330 20795
rect -330 20735 -314 20795
rect -56 20735 -4 20795
rect 34 20995 86 21055
rect 344 20995 396 21055
rect 434 20995 486 21055
rect 744 20995 796 21055
rect 834 20995 886 21055
rect 1144 20995 1196 21055
rect 1234 20995 1286 21055
rect 1544 20995 1596 21055
rect 1634 20995 1686 21055
rect 1944 20995 1996 21055
rect 2034 20995 2086 21055
rect 2344 20995 2396 21055
rect 2434 20995 2486 21055
rect 2744 20995 2796 21055
rect 2834 20995 2886 21055
rect 3144 20995 3196 21055
rect 3234 20995 3286 21055
rect 3544 20995 3596 21055
rect 3634 20995 3686 21055
rect 3944 20995 3996 21055
rect 4034 20995 4086 21055
rect 4344 20995 4396 21055
rect 4434 20995 4486 21055
rect 4744 20995 4796 21055
rect 4834 20995 4886 21055
rect 5144 20995 5196 21055
rect 5234 20995 5286 21055
rect 5544 20995 5596 21055
rect 5634 20995 5686 21055
rect 5944 20995 5996 21055
rect 6034 20995 6086 21055
rect 6344 20995 6396 21055
rect 6434 20995 6486 21055
rect 6744 20995 6796 21055
rect 6834 20995 6886 21055
rect 7144 20995 7196 21055
rect 7234 20995 7286 21055
rect 7544 20995 7596 21055
rect 7634 20995 7686 21055
rect 7944 20995 7996 21055
rect 8034 20995 8086 21055
rect 8344 20995 8396 21055
rect 8434 20995 8486 21055
rect 8744 20995 8796 21055
rect 8834 20995 8886 21055
rect 9144 20995 9196 21055
rect 9234 20995 9286 21055
rect 9544 20995 9596 21055
rect 9634 20995 9686 21055
rect 9944 20995 9996 21055
rect 10034 20995 10086 21055
rect 10344 20995 10396 21055
rect 10434 20995 10486 21055
rect 10744 20995 10796 21055
rect 10834 20995 10886 21055
rect 11144 20995 11196 21055
rect 11234 20995 11286 21055
rect 11544 20995 11596 21055
rect 11634 20995 11686 21055
rect 11944 20995 11996 21055
rect 12034 20995 12086 21055
rect 12344 20995 12396 21055
rect 12434 20995 12486 21055
rect 12744 20995 12796 21055
rect 12834 20995 12886 21055
rect 13144 20995 13196 21055
rect 34 20735 86 20795
rect 344 20735 396 20795
rect 434 20735 486 20795
rect 744 20735 796 20795
rect 834 20735 886 20795
rect 1144 20735 1196 20795
rect 1234 20735 1286 20795
rect 1544 20735 1596 20795
rect 1634 20735 1686 20795
rect 1944 20735 1996 20795
rect 2034 20735 2086 20795
rect 2344 20735 2396 20795
rect 2434 20735 2486 20795
rect 2744 20735 2796 20795
rect 2834 20735 2886 20795
rect 3144 20735 3196 20795
rect 3234 20735 3286 20795
rect 3544 20735 3596 20795
rect 3634 20735 3686 20795
rect 3944 20735 3996 20795
rect 4034 20735 4086 20795
rect 4344 20735 4396 20795
rect 4434 20735 4486 20795
rect 4744 20735 4796 20795
rect 4834 20735 4886 20795
rect 5144 20735 5196 20795
rect 5234 20735 5286 20795
rect 5544 20735 5596 20795
rect 5634 20735 5686 20795
rect 5944 20735 5996 20795
rect 6034 20735 6086 20795
rect 6344 20735 6396 20795
rect 6434 20735 6486 20795
rect 6744 20735 6796 20795
rect 6834 20735 6886 20795
rect 7144 20735 7196 20795
rect 7234 20735 7286 20795
rect 7544 20735 7596 20795
rect 7634 20735 7686 20795
rect 7944 20735 7996 20795
rect 8034 20735 8086 20795
rect 8344 20735 8396 20795
rect 8434 20735 8486 20795
rect 8744 20735 8796 20795
rect 8834 20735 8886 20795
rect 9144 20735 9196 20795
rect 9234 20735 9286 20795
rect 9544 20735 9596 20795
rect 9634 20735 9686 20795
rect 9944 20735 9996 20795
rect 10034 20735 10086 20795
rect 10344 20735 10396 20795
rect 10434 20735 10486 20795
rect 10744 20735 10796 20795
rect 10834 20735 10886 20795
rect 11144 20735 11196 20795
rect 11234 20735 11286 20795
rect 11544 20735 11596 20795
rect 11634 20735 11686 20795
rect 11944 20735 11996 20795
rect 12034 20735 12086 20795
rect 12344 20735 12396 20795
rect 12434 20735 12486 20795
rect 12744 20735 12796 20795
rect 12834 20735 12886 20795
rect 13144 20735 13196 20795
rect -366 20625 -330 20685
rect -330 20625 -314 20685
rect -56 20625 -4 20685
rect -366 20365 -330 20425
rect -330 20365 -314 20425
rect -56 20365 -4 20425
rect 34 20625 86 20685
rect 344 20625 396 20685
rect 434 20625 486 20685
rect 744 20625 796 20685
rect 834 20625 886 20685
rect 1144 20625 1196 20685
rect 1234 20625 1286 20685
rect 1544 20625 1596 20685
rect 1634 20625 1686 20685
rect 1944 20625 1996 20685
rect 2034 20625 2086 20685
rect 2344 20625 2396 20685
rect 2434 20625 2486 20685
rect 2744 20625 2796 20685
rect 2834 20625 2886 20685
rect 3144 20625 3196 20685
rect 3234 20625 3286 20685
rect 3544 20625 3596 20685
rect 3634 20625 3686 20685
rect 3944 20625 3996 20685
rect 4034 20625 4086 20685
rect 4344 20625 4396 20685
rect 4434 20625 4486 20685
rect 4744 20625 4796 20685
rect 4834 20625 4886 20685
rect 5144 20625 5196 20685
rect 5234 20625 5286 20685
rect 5544 20625 5596 20685
rect 5634 20625 5686 20685
rect 5944 20625 5996 20685
rect 6034 20625 6086 20685
rect 6344 20625 6396 20685
rect 6434 20625 6486 20685
rect 6744 20625 6796 20685
rect 6834 20625 6886 20685
rect 7144 20625 7196 20685
rect 7234 20625 7286 20685
rect 7544 20625 7596 20685
rect 7634 20625 7686 20685
rect 7944 20625 7996 20685
rect 8034 20625 8086 20685
rect 8344 20625 8396 20685
rect 8434 20625 8486 20685
rect 8744 20625 8796 20685
rect 8834 20625 8886 20685
rect 9144 20625 9196 20685
rect 9234 20625 9286 20685
rect 9544 20625 9596 20685
rect 9634 20625 9686 20685
rect 9944 20625 9996 20685
rect 10034 20625 10086 20685
rect 10344 20625 10396 20685
rect 10434 20625 10486 20685
rect 10744 20625 10796 20685
rect 10834 20625 10886 20685
rect 11144 20625 11196 20685
rect 11234 20625 11286 20685
rect 11544 20625 11596 20685
rect 11634 20625 11686 20685
rect 11944 20625 11996 20685
rect 12034 20625 12086 20685
rect 12344 20625 12396 20685
rect 12434 20625 12486 20685
rect 12744 20625 12796 20685
rect 12834 20625 12886 20685
rect 13144 20625 13196 20685
rect 34 20365 86 20425
rect 344 20365 396 20425
rect 434 20365 486 20425
rect 744 20365 796 20425
rect 834 20365 886 20425
rect 1144 20365 1196 20425
rect 1234 20365 1286 20425
rect 1544 20365 1596 20425
rect 1634 20365 1686 20425
rect 1944 20365 1996 20425
rect 2034 20365 2086 20425
rect 2344 20365 2396 20425
rect 2434 20365 2486 20425
rect 2744 20365 2796 20425
rect 2834 20365 2886 20425
rect 3144 20365 3196 20425
rect 3234 20365 3286 20425
rect 3544 20365 3596 20425
rect 3634 20365 3686 20425
rect 3944 20365 3996 20425
rect 4034 20365 4086 20425
rect 4344 20365 4396 20425
rect 4434 20365 4486 20425
rect 4744 20365 4796 20425
rect 4834 20365 4886 20425
rect 5144 20365 5196 20425
rect 5234 20365 5286 20425
rect 5544 20365 5596 20425
rect 5634 20365 5686 20425
rect 5944 20365 5996 20425
rect 6034 20365 6086 20425
rect 6344 20365 6396 20425
rect 6434 20365 6486 20425
rect 6744 20365 6796 20425
rect 6834 20365 6886 20425
rect 7144 20365 7196 20425
rect 7234 20365 7286 20425
rect 7544 20365 7596 20425
rect 7634 20365 7686 20425
rect 7944 20365 7996 20425
rect 8034 20365 8086 20425
rect 8344 20365 8396 20425
rect 8434 20365 8486 20425
rect 8744 20365 8796 20425
rect 8834 20365 8886 20425
rect 9144 20365 9196 20425
rect 9234 20365 9286 20425
rect 9544 20365 9596 20425
rect 9634 20365 9686 20425
rect 9944 20365 9996 20425
rect 10034 20365 10086 20425
rect 10344 20365 10396 20425
rect 10434 20365 10486 20425
rect 10744 20365 10796 20425
rect 10834 20365 10886 20425
rect 11144 20365 11196 20425
rect 11234 20365 11286 20425
rect 11544 20365 11596 20425
rect 11634 20365 11686 20425
rect 11944 20365 11996 20425
rect 12034 20365 12086 20425
rect 12344 20365 12396 20425
rect 12434 20365 12486 20425
rect 12744 20365 12796 20425
rect 12834 20365 12886 20425
rect 13144 20365 13196 20425
rect -366 20255 -330 20315
rect -330 20255 -314 20315
rect -56 20255 -4 20315
rect -366 19995 -330 20055
rect -330 19995 -314 20055
rect -56 19995 -4 20055
rect 34 20255 86 20315
rect 344 20255 396 20315
rect 434 20255 486 20315
rect 744 20255 796 20315
rect 834 20255 886 20315
rect 1144 20255 1196 20315
rect 1234 20255 1286 20315
rect 1544 20255 1596 20315
rect 1634 20255 1686 20315
rect 1944 20255 1996 20315
rect 2034 20255 2086 20315
rect 2344 20255 2396 20315
rect 2434 20255 2486 20315
rect 2744 20255 2796 20315
rect 2834 20255 2886 20315
rect 3144 20255 3196 20315
rect 3234 20255 3286 20315
rect 3544 20255 3596 20315
rect 3634 20255 3686 20315
rect 3944 20255 3996 20315
rect 4034 20255 4086 20315
rect 4344 20255 4396 20315
rect 4434 20255 4486 20315
rect 4744 20255 4796 20315
rect 4834 20255 4886 20315
rect 5144 20255 5196 20315
rect 5234 20255 5286 20315
rect 5544 20255 5596 20315
rect 5634 20255 5686 20315
rect 5944 20255 5996 20315
rect 6034 20255 6086 20315
rect 6344 20255 6396 20315
rect 6434 20255 6486 20315
rect 6744 20255 6796 20315
rect 6834 20255 6886 20315
rect 7144 20255 7196 20315
rect 7234 20255 7286 20315
rect 7544 20255 7596 20315
rect 7634 20255 7686 20315
rect 7944 20255 7996 20315
rect 8034 20255 8086 20315
rect 8344 20255 8396 20315
rect 8434 20255 8486 20315
rect 8744 20255 8796 20315
rect 8834 20255 8886 20315
rect 9144 20255 9196 20315
rect 9234 20255 9286 20315
rect 9544 20255 9596 20315
rect 9634 20255 9686 20315
rect 9944 20255 9996 20315
rect 10034 20255 10086 20315
rect 10344 20255 10396 20315
rect 10434 20255 10486 20315
rect 10744 20255 10796 20315
rect 10834 20255 10886 20315
rect 11144 20255 11196 20315
rect 11234 20255 11286 20315
rect 11544 20255 11596 20315
rect 11634 20255 11686 20315
rect 11944 20255 11996 20315
rect 12034 20255 12086 20315
rect 12344 20255 12396 20315
rect 12434 20255 12486 20315
rect 12744 20255 12796 20315
rect 12834 20255 12886 20315
rect 13144 20255 13196 20315
rect 34 19995 86 20055
rect 344 19995 396 20055
rect 434 19995 486 20055
rect 744 19995 796 20055
rect 834 19995 886 20055
rect 1144 19995 1196 20055
rect 1234 19995 1286 20055
rect 1544 19995 1596 20055
rect 1634 19995 1686 20055
rect 1944 19995 1996 20055
rect 2034 19995 2086 20055
rect 2344 19995 2396 20055
rect 2434 19995 2486 20055
rect 2744 19995 2796 20055
rect 2834 19995 2886 20055
rect 3144 19995 3196 20055
rect 3234 19995 3286 20055
rect 3544 19995 3596 20055
rect 3634 19995 3686 20055
rect 3944 19995 3996 20055
rect 4034 19995 4086 20055
rect 4344 19995 4396 20055
rect 4434 19995 4486 20055
rect 4744 19995 4796 20055
rect 4834 19995 4886 20055
rect 5144 19995 5196 20055
rect 5234 19995 5286 20055
rect 5544 19995 5596 20055
rect 5634 19995 5686 20055
rect 5944 19995 5996 20055
rect 6034 19995 6086 20055
rect 6344 19995 6396 20055
rect 6434 19995 6486 20055
rect 6744 19995 6796 20055
rect 6834 19995 6886 20055
rect 7144 19995 7196 20055
rect 7234 19995 7286 20055
rect 7544 19995 7596 20055
rect 7634 19995 7686 20055
rect 7944 19995 7996 20055
rect 8034 19995 8086 20055
rect 8344 19995 8396 20055
rect 8434 19995 8486 20055
rect 8744 19995 8796 20055
rect 8834 19995 8886 20055
rect 9144 19995 9196 20055
rect 9234 19995 9286 20055
rect 9544 19995 9596 20055
rect 9634 19995 9686 20055
rect 9944 19995 9996 20055
rect 10034 19995 10086 20055
rect 10344 19995 10396 20055
rect 10434 19995 10486 20055
rect 10744 19995 10796 20055
rect 10834 19995 10886 20055
rect 11144 19995 11196 20055
rect 11234 19995 11286 20055
rect 11544 19995 11596 20055
rect 11634 19995 11686 20055
rect 11944 19995 11996 20055
rect 12034 19995 12086 20055
rect 12344 19995 12396 20055
rect 12434 19995 12486 20055
rect 12744 19995 12796 20055
rect 12834 19995 12886 20055
rect 13144 19995 13196 20055
rect -366 19885 -330 19945
rect -330 19885 -314 19945
rect -56 19885 -4 19945
rect -366 19625 -330 19685
rect -330 19625 -314 19685
rect -56 19625 -4 19685
rect 34 19885 86 19945
rect 344 19885 396 19945
rect 434 19885 486 19945
rect 744 19885 796 19945
rect 834 19885 886 19945
rect 1144 19885 1196 19945
rect 1234 19885 1286 19945
rect 1544 19885 1596 19945
rect 1634 19885 1686 19945
rect 1944 19885 1996 19945
rect 2034 19885 2086 19945
rect 2344 19885 2396 19945
rect 2434 19885 2486 19945
rect 2744 19885 2796 19945
rect 2834 19885 2886 19945
rect 3144 19885 3196 19945
rect 3234 19885 3286 19945
rect 3544 19885 3596 19945
rect 3634 19885 3686 19945
rect 3944 19885 3996 19945
rect 4034 19885 4086 19945
rect 4344 19885 4396 19945
rect 4434 19885 4486 19945
rect 4744 19885 4796 19945
rect 4834 19885 4886 19945
rect 5144 19885 5196 19945
rect 5234 19885 5286 19945
rect 5544 19885 5596 19945
rect 5634 19885 5686 19945
rect 5944 19885 5996 19945
rect 6034 19885 6086 19945
rect 6344 19885 6396 19945
rect 6434 19885 6486 19945
rect 6744 19885 6796 19945
rect 6834 19885 6886 19945
rect 7144 19885 7196 19945
rect 7234 19885 7286 19945
rect 7544 19885 7596 19945
rect 7634 19885 7686 19945
rect 7944 19885 7996 19945
rect 8034 19885 8086 19945
rect 8344 19885 8396 19945
rect 8434 19885 8486 19945
rect 8744 19885 8796 19945
rect 8834 19885 8886 19945
rect 9144 19885 9196 19945
rect 9234 19885 9286 19945
rect 9544 19885 9596 19945
rect 9634 19885 9686 19945
rect 9944 19885 9996 19945
rect 10034 19885 10086 19945
rect 10344 19885 10396 19945
rect 10434 19885 10486 19945
rect 10744 19885 10796 19945
rect 10834 19885 10886 19945
rect 11144 19885 11196 19945
rect 11234 19885 11286 19945
rect 11544 19885 11596 19945
rect 11634 19885 11686 19945
rect 11944 19885 11996 19945
rect 12034 19885 12086 19945
rect 12344 19885 12396 19945
rect 12434 19885 12486 19945
rect 12744 19885 12796 19945
rect 12834 19885 12886 19945
rect 13144 19885 13196 19945
rect 34 19625 86 19685
rect 344 19625 396 19685
rect 434 19625 486 19685
rect 744 19625 796 19685
rect 834 19625 886 19685
rect 1144 19625 1196 19685
rect 1234 19625 1286 19685
rect 1544 19625 1596 19685
rect 1634 19625 1686 19685
rect 1944 19625 1996 19685
rect 2034 19625 2086 19685
rect 2344 19625 2396 19685
rect 2434 19625 2486 19685
rect 2744 19625 2796 19685
rect 2834 19625 2886 19685
rect 3144 19625 3196 19685
rect 3234 19625 3286 19685
rect 3544 19625 3596 19685
rect 3634 19625 3686 19685
rect 3944 19625 3996 19685
rect 4034 19625 4086 19685
rect 4344 19625 4396 19685
rect 4434 19625 4486 19685
rect 4744 19625 4796 19685
rect 4834 19625 4886 19685
rect 5144 19625 5196 19685
rect 5234 19625 5286 19685
rect 5544 19625 5596 19685
rect 5634 19625 5686 19685
rect 5944 19625 5996 19685
rect 6034 19625 6086 19685
rect 6344 19625 6396 19685
rect 6434 19625 6486 19685
rect 6744 19625 6796 19685
rect 6834 19625 6886 19685
rect 7144 19625 7196 19685
rect 7234 19625 7286 19685
rect 7544 19625 7596 19685
rect 7634 19625 7686 19685
rect 7944 19625 7996 19685
rect 8034 19625 8086 19685
rect 8344 19625 8396 19685
rect 8434 19625 8486 19685
rect 8744 19625 8796 19685
rect 8834 19625 8886 19685
rect 9144 19625 9196 19685
rect 9234 19625 9286 19685
rect 9544 19625 9596 19685
rect 9634 19625 9686 19685
rect 9944 19625 9996 19685
rect 10034 19625 10086 19685
rect 10344 19625 10396 19685
rect 10434 19625 10486 19685
rect 10744 19625 10796 19685
rect 10834 19625 10886 19685
rect 11144 19625 11196 19685
rect 11234 19625 11286 19685
rect 11544 19625 11596 19685
rect 11634 19625 11686 19685
rect 11944 19625 11996 19685
rect 12034 19625 12086 19685
rect 12344 19625 12396 19685
rect 12434 19625 12486 19685
rect 12744 19625 12796 19685
rect 12834 19625 12886 19685
rect 13144 19625 13196 19685
rect -366 19515 -330 19575
rect -330 19515 -314 19575
rect -56 19515 -4 19575
rect -366 19255 -330 19315
rect -330 19255 -314 19315
rect -56 19255 -4 19315
rect 34 19515 86 19575
rect 344 19515 396 19575
rect 434 19515 486 19575
rect 744 19515 796 19575
rect 834 19515 886 19575
rect 1144 19515 1196 19575
rect 1234 19515 1286 19575
rect 1544 19515 1596 19575
rect 1634 19515 1686 19575
rect 1944 19515 1996 19575
rect 2034 19515 2086 19575
rect 2344 19515 2396 19575
rect 2434 19515 2486 19575
rect 2744 19515 2796 19575
rect 2834 19515 2886 19575
rect 3144 19515 3196 19575
rect 34 19255 86 19315
rect 344 19255 396 19315
rect 434 19255 486 19315
rect 744 19255 796 19315
rect 834 19255 886 19315
rect 1144 19255 1196 19315
rect 1234 19255 1286 19315
rect 1544 19255 1596 19315
rect 1634 19255 1686 19315
rect 1944 19255 1996 19315
rect 2034 19255 2086 19315
rect 2344 19255 2396 19315
rect 2434 19255 2486 19315
rect 2744 19255 2796 19315
rect 2834 19255 2886 19315
rect 3144 19255 3196 19315
rect 3234 19515 3286 19575
rect 3544 19515 3596 19575
rect 3634 19515 3686 19575
rect 3944 19515 3996 19575
rect 4034 19515 4086 19575
rect 4344 19515 4396 19575
rect 4434 19515 4486 19575
rect 4744 19515 4796 19575
rect 4834 19515 4886 19575
rect 5144 19515 5196 19575
rect 5234 19515 5286 19575
rect 5544 19515 5596 19575
rect 5634 19515 5686 19575
rect 5944 19515 5996 19575
rect 6034 19515 6086 19575
rect 6344 19515 6396 19575
rect 6434 19515 6486 19575
rect 6744 19515 6796 19575
rect 6834 19515 6886 19575
rect 7144 19515 7196 19575
rect 7234 19515 7286 19575
rect 7544 19515 7596 19575
rect 7634 19515 7686 19575
rect 7944 19515 7996 19575
rect 8034 19515 8086 19575
rect 8344 19515 8396 19575
rect 8434 19515 8486 19575
rect 8744 19515 8796 19575
rect 8834 19515 8886 19575
rect 9144 19515 9196 19575
rect 9234 19515 9286 19575
rect 9544 19515 9596 19575
rect 9634 19515 9686 19575
rect 9944 19515 9996 19575
rect 10034 19515 10086 19575
rect 10344 19515 10396 19575
rect 10434 19515 10486 19575
rect 10744 19515 10796 19575
rect 10834 19515 10886 19575
rect 11144 19515 11196 19575
rect 11234 19515 11286 19575
rect 11544 19515 11596 19575
rect 11634 19515 11686 19575
rect 11944 19515 11996 19575
rect 12034 19515 12086 19575
rect 12344 19515 12396 19575
rect 12434 19515 12486 19575
rect 12744 19515 12796 19575
rect 12834 19515 12886 19575
rect 13144 19515 13196 19575
rect 3234 19255 3286 19315
rect 3544 19255 3596 19315
rect 3634 19255 3686 19315
rect 3944 19255 3996 19315
rect 4034 19255 4086 19315
rect 4344 19255 4396 19315
rect 4434 19255 4486 19315
rect 4744 19255 4796 19315
rect 4834 19255 4886 19315
rect 5144 19255 5196 19315
rect 5234 19255 5286 19315
rect 5544 19255 5596 19315
rect 5634 19255 5686 19315
rect 5944 19255 5996 19315
rect 6034 19255 6086 19315
rect 6344 19255 6396 19315
rect 6434 19255 6486 19315
rect 6744 19255 6796 19315
rect 6834 19255 6886 19315
rect 7144 19255 7196 19315
rect 7234 19255 7286 19315
rect 7544 19255 7596 19315
rect 7634 19255 7686 19315
rect 7944 19255 7996 19315
rect 8034 19255 8086 19315
rect 8344 19255 8396 19315
rect 8434 19255 8486 19315
rect 8744 19255 8796 19315
rect 8834 19255 8886 19315
rect 9144 19255 9196 19315
rect 9234 19255 9286 19315
rect 9544 19255 9596 19315
rect 9634 19255 9686 19315
rect 9944 19255 9996 19315
rect 10034 19255 10086 19315
rect 10344 19255 10396 19315
rect 10434 19255 10486 19315
rect 10744 19255 10796 19315
rect 10834 19255 10886 19315
rect 11144 19255 11196 19315
rect 11234 19255 11286 19315
rect 11544 19255 11596 19315
rect 11634 19255 11686 19315
rect 11944 19255 11996 19315
rect 12034 19255 12086 19315
rect 12344 19255 12396 19315
rect 12434 19255 12486 19315
rect 12744 19255 12796 19315
rect 12834 19255 12886 19315
rect 13144 19255 13196 19315
rect -366 19145 -330 19205
rect -330 19145 -314 19205
rect -56 19145 -4 19205
rect -366 18885 -330 18945
rect -330 18885 -314 18945
rect -56 18885 -4 18945
rect 34 19145 86 19205
rect 344 19145 396 19205
rect 434 19145 486 19205
rect 744 19145 796 19205
rect 834 19145 886 19205
rect 1144 19145 1196 19205
rect 1234 19145 1286 19205
rect 1544 19145 1596 19205
rect 1634 19145 1686 19205
rect 1944 19145 1996 19205
rect 2034 19145 2086 19205
rect 2344 19145 2396 19205
rect 2434 19145 2486 19205
rect 2744 19145 2796 19205
rect 2834 19145 2886 19205
rect 3144 19145 3196 19205
rect 34 18885 86 18945
rect 344 18885 396 18945
rect 434 18885 486 18945
rect 744 18885 796 18945
rect 834 18885 886 18945
rect 1144 18885 1196 18945
rect 1234 18885 1286 18945
rect 1544 18885 1596 18945
rect 1634 18885 1686 18945
rect 1944 18885 1996 18945
rect 2034 18885 2086 18945
rect 2344 18885 2396 18945
rect 2434 18885 2486 18945
rect 2744 18885 2796 18945
rect 2834 18885 2886 18945
rect 3144 18885 3196 18945
rect 3234 19145 3286 19205
rect 3544 19145 3596 19205
rect 3634 19145 3686 19205
rect 3944 19145 3996 19205
rect 4034 19145 4086 19205
rect 4344 19145 4396 19205
rect 4434 19145 4486 19205
rect 4744 19145 4796 19205
rect 4834 19145 4886 19205
rect 5144 19145 5196 19205
rect 5234 19145 5286 19205
rect 5544 19145 5596 19205
rect 5634 19145 5686 19205
rect 5944 19145 5996 19205
rect 6034 19145 6086 19205
rect 6344 19145 6396 19205
rect 6434 19145 6486 19205
rect 6744 19145 6796 19205
rect 6834 19145 6886 19205
rect 7144 19145 7196 19205
rect 7234 19145 7286 19205
rect 7544 19145 7596 19205
rect 7634 19145 7686 19205
rect 7944 19145 7996 19205
rect 8034 19145 8086 19205
rect 8344 19145 8396 19205
rect 8434 19145 8486 19205
rect 8744 19145 8796 19205
rect 8834 19145 8886 19205
rect 9144 19145 9196 19205
rect 9234 19145 9286 19205
rect 9544 19145 9596 19205
rect 9634 19145 9686 19205
rect 9944 19145 9996 19205
rect 10034 19145 10086 19205
rect 10344 19145 10396 19205
rect 10434 19145 10486 19205
rect 10744 19145 10796 19205
rect 10834 19145 10886 19205
rect 11144 19145 11196 19205
rect 11234 19145 11286 19205
rect 11544 19145 11596 19205
rect 11634 19145 11686 19205
rect 11944 19145 11996 19205
rect 12034 19145 12086 19205
rect 12344 19145 12396 19205
rect 12434 19145 12486 19205
rect 12744 19145 12796 19205
rect 12834 19145 12886 19205
rect 13144 19145 13196 19205
rect 3234 18885 3286 18945
rect 3544 18885 3596 18945
rect 3634 18885 3686 18945
rect 3944 18885 3996 18945
rect 4034 18885 4086 18945
rect 4344 18885 4396 18945
rect 4434 18885 4486 18945
rect 4744 18885 4796 18945
rect 4834 18885 4886 18945
rect 5144 18885 5196 18945
rect 5234 18885 5286 18945
rect 5544 18885 5596 18945
rect 5634 18885 5686 18945
rect 5944 18885 5996 18945
rect 6034 18885 6086 18945
rect 6344 18885 6396 18945
rect 6434 18885 6486 18945
rect 6744 18885 6796 18945
rect 6834 18885 6886 18945
rect 7144 18885 7196 18945
rect 7234 18885 7286 18945
rect 7544 18885 7596 18945
rect 7634 18885 7686 18945
rect 7944 18885 7996 18945
rect 8034 18885 8086 18945
rect 8344 18885 8396 18945
rect 8434 18885 8486 18945
rect 8744 18885 8796 18945
rect 8834 18885 8886 18945
rect 9144 18885 9196 18945
rect 9234 18885 9286 18945
rect 9544 18885 9596 18945
rect 9634 18885 9686 18945
rect 9944 18885 9996 18945
rect 10034 18885 10086 18945
rect 10344 18885 10396 18945
rect 10434 18885 10486 18945
rect 10744 18885 10796 18945
rect 10834 18885 10886 18945
rect 11144 18885 11196 18945
rect 11234 18885 11286 18945
rect 11544 18885 11596 18945
rect 11634 18885 11686 18945
rect 11944 18885 11996 18945
rect 12034 18885 12086 18945
rect 12344 18885 12396 18945
rect 12434 18885 12486 18945
rect 12744 18885 12796 18945
rect 12834 18885 12886 18945
rect 13144 18885 13196 18945
rect -366 18775 -330 18835
rect -330 18775 -314 18835
rect -56 18775 -4 18835
rect -366 18515 -330 18575
rect -330 18515 -314 18575
rect -56 18515 -4 18575
rect 34 18775 86 18835
rect 344 18775 396 18835
rect 434 18775 486 18835
rect 744 18775 796 18835
rect 834 18775 886 18835
rect 1144 18775 1196 18835
rect 1234 18775 1286 18835
rect 1544 18775 1596 18835
rect 1634 18775 1686 18835
rect 1944 18775 1996 18835
rect 2034 18775 2086 18835
rect 2344 18775 2396 18835
rect 2434 18775 2486 18835
rect 2744 18775 2796 18835
rect 2834 18775 2886 18835
rect 3144 18775 3196 18835
rect 34 18515 86 18575
rect 344 18515 396 18575
rect 434 18515 486 18575
rect 744 18515 796 18575
rect 834 18515 886 18575
rect 1144 18515 1196 18575
rect 1234 18515 1286 18575
rect 1544 18515 1596 18575
rect 1634 18515 1686 18575
rect 1944 18515 1996 18575
rect 2034 18515 2086 18575
rect 2344 18515 2396 18575
rect 2434 18515 2486 18575
rect 2744 18515 2796 18575
rect 2834 18515 2886 18575
rect 3144 18515 3196 18575
rect 3234 18775 3286 18835
rect 3544 18775 3596 18835
rect 3634 18775 3686 18835
rect 3944 18775 3996 18835
rect 4034 18775 4086 18835
rect 4344 18775 4396 18835
rect 4434 18775 4486 18835
rect 4744 18775 4796 18835
rect 4834 18775 4886 18835
rect 5144 18775 5196 18835
rect 5234 18775 5286 18835
rect 5544 18775 5596 18835
rect 5634 18775 5686 18835
rect 5944 18775 5996 18835
rect 6034 18775 6086 18835
rect 6344 18775 6396 18835
rect 6434 18775 6486 18835
rect 6744 18775 6796 18835
rect 6834 18775 6886 18835
rect 7144 18775 7196 18835
rect 7234 18775 7286 18835
rect 7544 18775 7596 18835
rect 7634 18775 7686 18835
rect 7944 18775 7996 18835
rect 8034 18775 8086 18835
rect 8344 18775 8396 18835
rect 8434 18775 8486 18835
rect 8744 18775 8796 18835
rect 8834 18775 8886 18835
rect 9144 18775 9196 18835
rect 9234 18775 9286 18835
rect 9544 18775 9596 18835
rect 9634 18775 9686 18835
rect 9944 18775 9996 18835
rect 10034 18775 10086 18835
rect 10344 18775 10396 18835
rect 10434 18775 10486 18835
rect 10744 18775 10796 18835
rect 10834 18775 10886 18835
rect 11144 18775 11196 18835
rect 11234 18775 11286 18835
rect 11544 18775 11596 18835
rect 11634 18775 11686 18835
rect 11944 18775 11996 18835
rect 12034 18775 12086 18835
rect 12344 18775 12396 18835
rect 12434 18775 12486 18835
rect 12744 18775 12796 18835
rect 12834 18775 12886 18835
rect 13144 18775 13196 18835
rect 3234 18515 3286 18575
rect 3544 18515 3596 18575
rect 3634 18515 3686 18575
rect 3944 18515 3996 18575
rect 4034 18515 4086 18575
rect 4344 18515 4396 18575
rect 4434 18515 4486 18575
rect 4744 18515 4796 18575
rect 4834 18515 4886 18575
rect 5144 18515 5196 18575
rect 5234 18515 5286 18575
rect 5544 18515 5596 18575
rect 5634 18515 5686 18575
rect 5944 18515 5996 18575
rect 6034 18515 6086 18575
rect 6344 18515 6396 18575
rect 6434 18515 6486 18575
rect 6744 18515 6796 18575
rect 6834 18515 6886 18575
rect 7144 18515 7196 18575
rect 7234 18515 7286 18575
rect 7544 18515 7596 18575
rect 7634 18515 7686 18575
rect 7944 18515 7996 18575
rect 8034 18515 8086 18575
rect 8344 18515 8396 18575
rect 8434 18515 8486 18575
rect 8744 18515 8796 18575
rect 8834 18515 8886 18575
rect 9144 18515 9196 18575
rect 9234 18515 9286 18575
rect 9544 18515 9596 18575
rect 9634 18515 9686 18575
rect 9944 18515 9996 18575
rect 10034 18515 10086 18575
rect 10344 18515 10396 18575
rect 10434 18515 10486 18575
rect 10744 18515 10796 18575
rect 10834 18515 10886 18575
rect 11144 18515 11196 18575
rect 11234 18515 11286 18575
rect 11544 18515 11596 18575
rect 11634 18515 11686 18575
rect 11944 18515 11996 18575
rect 12034 18515 12086 18575
rect 12344 18515 12396 18575
rect 12434 18515 12486 18575
rect 12744 18515 12796 18575
rect 12834 18515 12886 18575
rect 13144 18515 13196 18575
rect -366 18405 -330 18465
rect -330 18405 -314 18465
rect -56 18405 -4 18465
rect -366 18145 -330 18205
rect -330 18145 -314 18205
rect -56 18145 -4 18205
rect 34 18405 86 18465
rect 344 18405 396 18465
rect 434 18405 486 18465
rect 744 18405 796 18465
rect 834 18405 886 18465
rect 1144 18405 1196 18465
rect 1234 18405 1286 18465
rect 1544 18405 1596 18465
rect 1634 18405 1686 18465
rect 1944 18405 1996 18465
rect 2034 18405 2086 18465
rect 2344 18405 2396 18465
rect 2434 18405 2486 18465
rect 2744 18405 2796 18465
rect 2834 18405 2886 18465
rect 3144 18405 3196 18465
rect 34 18145 86 18205
rect 344 18145 396 18205
rect 434 18145 486 18205
rect 744 18145 796 18205
rect 834 18145 886 18205
rect 1144 18145 1196 18205
rect 1234 18145 1286 18205
rect 1544 18145 1596 18205
rect 1634 18145 1686 18205
rect 1944 18145 1996 18205
rect 2034 18145 2086 18205
rect 2344 18145 2396 18205
rect 2434 18145 2486 18205
rect 2744 18145 2796 18205
rect 2834 18145 2886 18205
rect 3144 18145 3196 18205
rect 3234 18405 3286 18465
rect 3544 18405 3596 18465
rect 3634 18405 3686 18465
rect 3944 18405 3996 18465
rect 4034 18405 4086 18465
rect 4344 18405 4396 18465
rect 4434 18405 4486 18465
rect 4744 18405 4796 18465
rect 4834 18405 4886 18465
rect 5144 18405 5196 18465
rect 5234 18405 5286 18465
rect 5544 18405 5596 18465
rect 5634 18405 5686 18465
rect 5944 18405 5996 18465
rect 6034 18405 6086 18465
rect 6344 18405 6396 18465
rect 6434 18405 6486 18465
rect 6744 18405 6796 18465
rect 6834 18405 6886 18465
rect 7144 18405 7196 18465
rect 7234 18405 7286 18465
rect 7544 18405 7596 18465
rect 7634 18405 7686 18465
rect 7944 18405 7996 18465
rect 8034 18405 8086 18465
rect 8344 18405 8396 18465
rect 8434 18405 8486 18465
rect 8744 18405 8796 18465
rect 8834 18405 8886 18465
rect 9144 18405 9196 18465
rect 9234 18405 9286 18465
rect 9544 18405 9596 18465
rect 9634 18405 9686 18465
rect 9944 18405 9996 18465
rect 10034 18405 10086 18465
rect 10344 18405 10396 18465
rect 10434 18405 10486 18465
rect 10744 18405 10796 18465
rect 10834 18405 10886 18465
rect 11144 18405 11196 18465
rect 11234 18405 11286 18465
rect 11544 18405 11596 18465
rect 11634 18405 11686 18465
rect 11944 18405 11996 18465
rect 12034 18405 12086 18465
rect 12344 18405 12396 18465
rect 12434 18405 12486 18465
rect 12744 18405 12796 18465
rect 12834 18405 12886 18465
rect 13144 18405 13196 18465
rect 3234 18145 3286 18205
rect 3544 18145 3596 18205
rect 3634 18145 3686 18205
rect 3944 18145 3996 18205
rect 4034 18145 4086 18205
rect 4344 18145 4396 18205
rect 4434 18145 4486 18205
rect 4744 18145 4796 18205
rect 4834 18145 4886 18205
rect 5144 18145 5196 18205
rect 5234 18145 5286 18205
rect 5544 18145 5596 18205
rect 5634 18145 5686 18205
rect 5944 18145 5996 18205
rect 6034 18145 6086 18205
rect 6344 18145 6396 18205
rect 6434 18145 6486 18205
rect 6744 18145 6796 18205
rect 6834 18145 6886 18205
rect 7144 18145 7196 18205
rect 7234 18145 7286 18205
rect 7544 18145 7596 18205
rect 7634 18145 7686 18205
rect 7944 18145 7996 18205
rect 8034 18145 8086 18205
rect 8344 18145 8396 18205
rect 8434 18145 8486 18205
rect 8744 18145 8796 18205
rect 8834 18145 8886 18205
rect 9144 18145 9196 18205
rect 9234 18145 9286 18205
rect 9544 18145 9596 18205
rect 9634 18145 9686 18205
rect 9944 18145 9996 18205
rect 10034 18145 10086 18205
rect 10344 18145 10396 18205
rect 10434 18145 10486 18205
rect 10744 18145 10796 18205
rect 10834 18145 10886 18205
rect 11144 18145 11196 18205
rect 11234 18145 11286 18205
rect 11544 18145 11596 18205
rect 11634 18145 11686 18205
rect 11944 18145 11996 18205
rect 12034 18145 12086 18205
rect 12344 18145 12396 18205
rect 12434 18145 12486 18205
rect 12744 18145 12796 18205
rect 12834 18145 12886 18205
rect 13144 18145 13196 18205
rect -366 18035 -330 18095
rect -330 18035 -314 18095
rect -56 18035 -4 18095
rect -366 17775 -330 17835
rect -330 17775 -314 17835
rect -56 17775 -4 17835
rect 34 18035 86 18095
rect 344 18035 396 18095
rect 434 18035 486 18095
rect 744 18035 796 18095
rect 834 18035 886 18095
rect 1144 18035 1196 18095
rect 1234 18035 1286 18095
rect 1544 18035 1596 18095
rect 1634 18035 1686 18095
rect 1944 18035 1996 18095
rect 2034 18035 2086 18095
rect 2344 18035 2396 18095
rect 2434 18035 2486 18095
rect 2744 18035 2796 18095
rect 2834 18035 2886 18095
rect 3144 18035 3196 18095
rect 34 17775 86 17835
rect 344 17775 396 17835
rect 434 17775 486 17835
rect 744 17775 796 17835
rect 834 17775 886 17835
rect 1144 17775 1196 17835
rect 1234 17775 1286 17835
rect 1544 17775 1596 17835
rect 1634 17775 1686 17835
rect 1944 17775 1996 17835
rect 2034 17775 2086 17835
rect 2344 17775 2396 17835
rect 2434 17775 2486 17835
rect 2744 17775 2796 17835
rect 2834 17775 2886 17835
rect 3144 17775 3196 17835
rect 3234 18035 3286 18095
rect 3544 18035 3596 18095
rect 3634 18035 3686 18095
rect 3944 18035 3996 18095
rect 4034 18035 4086 18095
rect 4344 18035 4396 18095
rect 4434 18035 4486 18095
rect 4744 18035 4796 18095
rect 4834 18035 4886 18095
rect 5144 18035 5196 18095
rect 5234 18035 5286 18095
rect 5544 18035 5596 18095
rect 5634 18035 5686 18095
rect 5944 18035 5996 18095
rect 6034 18035 6086 18095
rect 6344 18035 6396 18095
rect 6434 18035 6486 18095
rect 6744 18035 6796 18095
rect 6834 18035 6886 18095
rect 7144 18035 7196 18095
rect 7234 18035 7286 18095
rect 7544 18035 7596 18095
rect 7634 18035 7686 18095
rect 7944 18035 7996 18095
rect 8034 18035 8086 18095
rect 8344 18035 8396 18095
rect 8434 18035 8486 18095
rect 8744 18035 8796 18095
rect 8834 18035 8886 18095
rect 9144 18035 9196 18095
rect 9234 18035 9286 18095
rect 9544 18035 9596 18095
rect 9634 18035 9686 18095
rect 9944 18035 9996 18095
rect 10034 18035 10086 18095
rect 10344 18035 10396 18095
rect 10434 18035 10486 18095
rect 10744 18035 10796 18095
rect 10834 18035 10886 18095
rect 11144 18035 11196 18095
rect 11234 18035 11286 18095
rect 11544 18035 11596 18095
rect 11634 18035 11686 18095
rect 11944 18035 11996 18095
rect 12034 18035 12086 18095
rect 12344 18035 12396 18095
rect 12434 18035 12486 18095
rect 12744 18035 12796 18095
rect 12834 18035 12886 18095
rect 13144 18035 13196 18095
rect 3234 17775 3286 17835
rect 3544 17775 3596 17835
rect 3634 17775 3686 17835
rect 3944 17775 3996 17835
rect 4034 17775 4086 17835
rect 4344 17775 4396 17835
rect 4434 17775 4486 17835
rect 4744 17775 4796 17835
rect 4834 17775 4886 17835
rect 5144 17775 5196 17835
rect 5234 17775 5286 17835
rect 5544 17775 5596 17835
rect 5634 17775 5686 17835
rect 5944 17775 5996 17835
rect 6034 17775 6086 17835
rect 6344 17775 6396 17835
rect 6434 17775 6486 17835
rect 6744 17775 6796 17835
rect 6834 17775 6886 17835
rect 7144 17775 7196 17835
rect 7234 17775 7286 17835
rect 7544 17775 7596 17835
rect 7634 17775 7686 17835
rect 7944 17775 7996 17835
rect 8034 17775 8086 17835
rect 8344 17775 8396 17835
rect 8434 17775 8486 17835
rect 8744 17775 8796 17835
rect 8834 17775 8886 17835
rect 9144 17775 9196 17835
rect 9234 17775 9286 17835
rect 9544 17775 9596 17835
rect 9634 17775 9686 17835
rect 9944 17775 9996 17835
rect 10034 17775 10086 17835
rect 10344 17775 10396 17835
rect 10434 17775 10486 17835
rect 10744 17775 10796 17835
rect 10834 17775 10886 17835
rect 11144 17775 11196 17835
rect 11234 17775 11286 17835
rect 11544 17775 11596 17835
rect 11634 17775 11686 17835
rect 11944 17775 11996 17835
rect 12034 17775 12086 17835
rect 12344 17775 12396 17835
rect 12434 17775 12486 17835
rect 12744 17775 12796 17835
rect 12834 17775 12886 17835
rect 13144 17775 13196 17835
rect -366 17665 -330 17725
rect -330 17665 -314 17725
rect -56 17665 -4 17725
rect -366 17405 -330 17465
rect -330 17405 -314 17465
rect -56 17405 -4 17465
rect 34 17665 86 17725
rect 344 17665 396 17725
rect 434 17665 486 17725
rect 744 17665 796 17725
rect 834 17665 886 17725
rect 1144 17665 1196 17725
rect 1234 17665 1286 17725
rect 1544 17665 1596 17725
rect 1634 17665 1686 17725
rect 1944 17665 1996 17725
rect 2034 17665 2086 17725
rect 2344 17665 2396 17725
rect 2434 17665 2486 17725
rect 2744 17665 2796 17725
rect 2834 17665 2886 17725
rect 3144 17665 3196 17725
rect 34 17405 86 17465
rect 344 17405 396 17465
rect 434 17405 486 17465
rect 744 17405 796 17465
rect 834 17405 886 17465
rect 1144 17405 1196 17465
rect 1234 17405 1286 17465
rect 1544 17405 1596 17465
rect 1634 17405 1686 17465
rect 1944 17405 1996 17465
rect 2034 17405 2086 17465
rect 2344 17405 2396 17465
rect 2434 17405 2486 17465
rect 2744 17405 2796 17465
rect 2834 17405 2886 17465
rect 3144 17405 3196 17465
rect 3234 17665 3286 17725
rect 3544 17665 3596 17725
rect 3634 17665 3686 17725
rect 3944 17665 3996 17725
rect 4034 17665 4086 17725
rect 4344 17665 4396 17725
rect 4434 17665 4486 17725
rect 4744 17665 4796 17725
rect 4834 17665 4886 17725
rect 5144 17665 5196 17725
rect 5234 17665 5286 17725
rect 5544 17665 5596 17725
rect 5634 17665 5686 17725
rect 5944 17665 5996 17725
rect 6034 17665 6086 17725
rect 6344 17665 6396 17725
rect 6434 17665 6486 17725
rect 6744 17665 6796 17725
rect 6834 17665 6886 17725
rect 7144 17665 7196 17725
rect 7234 17665 7286 17725
rect 7544 17665 7596 17725
rect 7634 17665 7686 17725
rect 7944 17665 7996 17725
rect 8034 17665 8086 17725
rect 8344 17665 8396 17725
rect 8434 17665 8486 17725
rect 8744 17665 8796 17725
rect 8834 17665 8886 17725
rect 9144 17665 9196 17725
rect 9234 17665 9286 17725
rect 9544 17665 9596 17725
rect 9634 17665 9686 17725
rect 9944 17665 9996 17725
rect 10034 17665 10086 17725
rect 10344 17665 10396 17725
rect 10434 17665 10486 17725
rect 10744 17665 10796 17725
rect 10834 17665 10886 17725
rect 11144 17665 11196 17725
rect 11234 17665 11286 17725
rect 11544 17665 11596 17725
rect 11634 17665 11686 17725
rect 11944 17665 11996 17725
rect 12034 17665 12086 17725
rect 12344 17665 12396 17725
rect 12434 17665 12486 17725
rect 12744 17665 12796 17725
rect 12834 17665 12886 17725
rect 13144 17665 13196 17725
rect 3234 17405 3286 17465
rect 3544 17405 3596 17465
rect 3634 17405 3686 17465
rect 3944 17405 3996 17465
rect 4034 17405 4086 17465
rect 4344 17405 4396 17465
rect 4434 17405 4486 17465
rect 4744 17405 4796 17465
rect 4834 17405 4886 17465
rect 5144 17405 5196 17465
rect 5234 17405 5286 17465
rect 5544 17405 5596 17465
rect 5634 17405 5686 17465
rect 5944 17405 5996 17465
rect 6034 17405 6086 17465
rect 6344 17405 6396 17465
rect 6434 17405 6486 17465
rect 6744 17405 6796 17465
rect 6834 17405 6886 17465
rect 7144 17405 7196 17465
rect 7234 17405 7286 17465
rect 7544 17405 7596 17465
rect 7634 17405 7686 17465
rect 7944 17405 7996 17465
rect 8034 17405 8086 17465
rect 8344 17405 8396 17465
rect 8434 17405 8486 17465
rect 8744 17405 8796 17465
rect 8834 17405 8886 17465
rect 9144 17405 9196 17465
rect 9234 17405 9286 17465
rect 9544 17405 9596 17465
rect 9634 17405 9686 17465
rect 9944 17405 9996 17465
rect 10034 17405 10086 17465
rect 10344 17405 10396 17465
rect 10434 17405 10486 17465
rect 10744 17405 10796 17465
rect 10834 17405 10886 17465
rect 11144 17405 11196 17465
rect 11234 17405 11286 17465
rect 11544 17405 11596 17465
rect 11634 17405 11686 17465
rect 11944 17405 11996 17465
rect 12034 17405 12086 17465
rect 12344 17405 12396 17465
rect 12434 17405 12486 17465
rect 12744 17405 12796 17465
rect 12834 17405 12886 17465
rect 13144 17405 13196 17465
rect -366 17295 -330 17355
rect -330 17295 -314 17355
rect -56 17295 -4 17355
rect -366 17035 -330 17095
rect -330 17035 -314 17095
rect -56 17035 -4 17095
rect 34 17295 86 17355
rect 344 17295 396 17355
rect 434 17295 486 17355
rect 744 17295 796 17355
rect 834 17295 886 17355
rect 1144 17295 1196 17355
rect 1234 17295 1286 17355
rect 1544 17295 1596 17355
rect 1634 17295 1686 17355
rect 1944 17295 1996 17355
rect 2034 17295 2086 17355
rect 2344 17295 2396 17355
rect 2434 17295 2486 17355
rect 2744 17295 2796 17355
rect 2834 17295 2886 17355
rect 3144 17295 3196 17355
rect 34 17035 86 17095
rect 344 17035 396 17095
rect 434 17035 486 17095
rect 744 17035 796 17095
rect 834 17035 886 17095
rect 1144 17035 1196 17095
rect 1234 17035 1286 17095
rect 1544 17035 1596 17095
rect 1634 17035 1686 17095
rect 1944 17035 1996 17095
rect 2034 17035 2086 17095
rect 2344 17035 2396 17095
rect 2434 17035 2486 17095
rect 2744 17035 2796 17095
rect 2834 17035 2886 17095
rect 3144 17035 3196 17095
rect 3234 17295 3286 17355
rect 3544 17295 3596 17355
rect 3634 17295 3686 17355
rect 3944 17295 3996 17355
rect 4034 17295 4086 17355
rect 4344 17295 4396 17355
rect 4434 17295 4486 17355
rect 4744 17295 4796 17355
rect 4834 17295 4886 17355
rect 5144 17295 5196 17355
rect 5234 17295 5286 17355
rect 5544 17295 5596 17355
rect 5634 17295 5686 17355
rect 5944 17295 5996 17355
rect 3234 17035 3286 17095
rect 3544 17035 3596 17095
rect 3634 17035 3686 17095
rect 3944 17035 3996 17095
rect 4034 17035 4086 17095
rect 4344 17035 4396 17095
rect 4434 17035 4486 17095
rect 4744 17035 4796 17095
rect 4834 17035 4886 17095
rect 5144 17035 5196 17095
rect 5234 17035 5286 17095
rect 5544 17035 5596 17095
rect 5634 17035 5686 17095
rect 5944 17035 5996 17095
rect 6034 17295 6086 17355
rect 6344 17295 6396 17355
rect 6434 17295 6486 17355
rect 6744 17295 6796 17355
rect 6834 17295 6886 17355
rect 7144 17295 7196 17355
rect 7234 17295 7286 17355
rect 7544 17295 7596 17355
rect 7634 17295 7686 17355
rect 7944 17295 7996 17355
rect 8034 17295 8086 17355
rect 8344 17295 8396 17355
rect 8434 17295 8486 17355
rect 8744 17295 8796 17355
rect 8834 17295 8886 17355
rect 9144 17295 9196 17355
rect 9234 17295 9286 17355
rect 9544 17295 9596 17355
rect 9634 17295 9686 17355
rect 9944 17295 9996 17355
rect 10034 17295 10086 17355
rect 10344 17295 10396 17355
rect 10434 17295 10486 17355
rect 10744 17295 10796 17355
rect 10834 17295 10886 17355
rect 11144 17295 11196 17355
rect 11234 17295 11286 17355
rect 11544 17295 11596 17355
rect 11634 17295 11686 17355
rect 11944 17295 11996 17355
rect 12034 17295 12086 17355
rect 12344 17295 12396 17355
rect 12434 17295 12486 17355
rect 12744 17295 12796 17355
rect 12834 17295 12886 17355
rect 13144 17295 13196 17355
rect 6034 17035 6086 17095
rect 6344 17035 6396 17095
rect 6434 17035 6486 17095
rect 6744 17035 6796 17095
rect 6834 17035 6886 17095
rect 7144 17035 7196 17095
rect 7234 17035 7286 17095
rect 7544 17035 7596 17095
rect 7634 17035 7686 17095
rect 7944 17035 7996 17095
rect 8034 17035 8086 17095
rect 8344 17035 8396 17095
rect 8434 17035 8486 17095
rect 8744 17035 8796 17095
rect 8834 17035 8886 17095
rect 9144 17035 9196 17095
rect 9234 17035 9286 17095
rect 9544 17035 9596 17095
rect 9634 17035 9686 17095
rect 9944 17035 9996 17095
rect 10034 17035 10086 17095
rect 10344 17035 10396 17095
rect 10434 17035 10486 17095
rect 10744 17035 10796 17095
rect 10834 17035 10886 17095
rect 11144 17035 11196 17095
rect 11234 17035 11286 17095
rect 11544 17035 11596 17095
rect 11634 17035 11686 17095
rect 11944 17035 11996 17095
rect 12034 17035 12086 17095
rect 12344 17035 12396 17095
rect 12434 17035 12486 17095
rect 12744 17035 12796 17095
rect 12834 17035 12886 17095
rect 13144 17035 13196 17095
rect -366 16925 -330 16985
rect -330 16925 -314 16985
rect -56 16925 -4 16985
rect -366 16665 -330 16725
rect -330 16665 -314 16725
rect -56 16665 -4 16725
rect 34 16925 86 16985
rect 344 16925 396 16985
rect 434 16925 486 16985
rect 744 16925 796 16985
rect 834 16925 886 16985
rect 1144 16925 1196 16985
rect 1234 16925 1286 16985
rect 1544 16925 1596 16985
rect 1634 16925 1686 16985
rect 1944 16925 1996 16985
rect 2034 16925 2086 16985
rect 2344 16925 2396 16985
rect 2434 16925 2486 16985
rect 2744 16925 2796 16985
rect 2834 16925 2886 16985
rect 3144 16925 3196 16985
rect 34 16665 86 16725
rect 344 16665 396 16725
rect 434 16665 486 16725
rect 744 16665 796 16725
rect 834 16665 886 16725
rect 1144 16665 1196 16725
rect 1234 16665 1286 16725
rect 1544 16665 1596 16725
rect 1634 16665 1686 16725
rect 1944 16665 1996 16725
rect 2034 16665 2086 16725
rect 2344 16665 2396 16725
rect 2434 16665 2486 16725
rect 2744 16665 2796 16725
rect 2834 16665 2886 16725
rect 3144 16665 3196 16725
rect 3234 16925 3286 16985
rect 3544 16925 3596 16985
rect 3634 16925 3686 16985
rect 3944 16925 3996 16985
rect 4034 16925 4086 16985
rect 4344 16925 4396 16985
rect 4434 16925 4486 16985
rect 4744 16925 4796 16985
rect 4834 16925 4886 16985
rect 5144 16925 5196 16985
rect 5234 16925 5286 16985
rect 5544 16925 5596 16985
rect 5634 16925 5686 16985
rect 5944 16925 5996 16985
rect 3234 16665 3286 16725
rect 3544 16665 3596 16725
rect 3634 16665 3686 16725
rect 3944 16665 3996 16725
rect 4034 16665 4086 16725
rect 4344 16665 4396 16725
rect 4434 16665 4486 16725
rect 4744 16665 4796 16725
rect 4834 16665 4886 16725
rect 5144 16665 5196 16725
rect 5234 16665 5286 16725
rect 5544 16665 5596 16725
rect 5634 16665 5686 16725
rect 5944 16665 5996 16725
rect 6034 16925 6086 16985
rect 6344 16925 6396 16985
rect 6434 16925 6486 16985
rect 6744 16925 6796 16985
rect 6834 16925 6886 16985
rect 7144 16925 7196 16985
rect 7234 16925 7286 16985
rect 7544 16925 7596 16985
rect 7634 16925 7686 16985
rect 7944 16925 7996 16985
rect 8034 16925 8086 16985
rect 8344 16925 8396 16985
rect 8434 16925 8486 16985
rect 8744 16925 8796 16985
rect 8834 16925 8886 16985
rect 9144 16925 9196 16985
rect 9234 16925 9286 16985
rect 9544 16925 9596 16985
rect 9634 16925 9686 16985
rect 9944 16925 9996 16985
rect 10034 16925 10086 16985
rect 10344 16925 10396 16985
rect 10434 16925 10486 16985
rect 10744 16925 10796 16985
rect 10834 16925 10886 16985
rect 11144 16925 11196 16985
rect 11234 16925 11286 16985
rect 11544 16925 11596 16985
rect 11634 16925 11686 16985
rect 11944 16925 11996 16985
rect 12034 16925 12086 16985
rect 12344 16925 12396 16985
rect 12434 16925 12486 16985
rect 12744 16925 12796 16985
rect 12834 16925 12886 16985
rect 13144 16925 13196 16985
rect 6034 16665 6086 16725
rect 6344 16665 6396 16725
rect 6434 16665 6486 16725
rect 6744 16665 6796 16725
rect 6834 16665 6886 16725
rect 7144 16665 7196 16725
rect 7234 16665 7286 16725
rect 7544 16665 7596 16725
rect 7634 16665 7686 16725
rect 7944 16665 7996 16725
rect 8034 16665 8086 16725
rect 8344 16665 8396 16725
rect 8434 16665 8486 16725
rect 8744 16665 8796 16725
rect 8834 16665 8886 16725
rect 9144 16665 9196 16725
rect 9234 16665 9286 16725
rect 9544 16665 9596 16725
rect 9634 16665 9686 16725
rect 9944 16665 9996 16725
rect 10034 16665 10086 16725
rect 10344 16665 10396 16725
rect 10434 16665 10486 16725
rect 10744 16665 10796 16725
rect 10834 16665 10886 16725
rect 11144 16665 11196 16725
rect 11234 16665 11286 16725
rect 11544 16665 11596 16725
rect 11634 16665 11686 16725
rect 11944 16665 11996 16725
rect 12034 16665 12086 16725
rect 12344 16665 12396 16725
rect 12434 16665 12486 16725
rect 12744 16665 12796 16725
rect 12834 16665 12886 16725
rect 13144 16665 13196 16725
rect -366 16555 -330 16615
rect -330 16555 -314 16615
rect -56 16555 -4 16615
rect -366 16295 -330 16355
rect -330 16295 -314 16355
rect -56 16295 -4 16355
rect 34 16555 86 16615
rect 344 16555 396 16615
rect 434 16555 486 16615
rect 744 16555 796 16615
rect 834 16555 886 16615
rect 1144 16555 1196 16615
rect 1234 16555 1286 16615
rect 1544 16555 1596 16615
rect 1634 16555 1686 16615
rect 1944 16555 1996 16615
rect 2034 16555 2086 16615
rect 2344 16555 2396 16615
rect 2434 16555 2486 16615
rect 2744 16555 2796 16615
rect 2834 16555 2886 16615
rect 3144 16555 3196 16615
rect 34 16295 86 16355
rect 344 16295 396 16355
rect 434 16295 486 16355
rect 744 16295 796 16355
rect 834 16295 886 16355
rect 1144 16295 1196 16355
rect 1234 16295 1286 16355
rect 1544 16295 1596 16355
rect 1634 16295 1686 16355
rect 1944 16295 1996 16355
rect 2034 16295 2086 16355
rect 2344 16295 2396 16355
rect 2434 16295 2486 16355
rect 2744 16295 2796 16355
rect 2834 16295 2886 16355
rect 3144 16295 3196 16355
rect 3234 16555 3286 16615
rect 3544 16555 3596 16615
rect 3634 16555 3686 16615
rect 3944 16555 3996 16615
rect 4034 16555 4086 16615
rect 4344 16555 4396 16615
rect 4434 16555 4486 16615
rect 4744 16555 4796 16615
rect 4834 16555 4886 16615
rect 5144 16555 5196 16615
rect 5234 16555 5286 16615
rect 5544 16555 5596 16615
rect 5634 16555 5686 16615
rect 5944 16555 5996 16615
rect 3234 16295 3286 16355
rect 3544 16295 3596 16355
rect 3634 16295 3686 16355
rect 3944 16295 3996 16355
rect 4034 16295 4086 16355
rect 4344 16295 4396 16355
rect 4434 16295 4486 16355
rect 4744 16295 4796 16355
rect 4834 16295 4886 16355
rect 5144 16295 5196 16355
rect 5234 16295 5286 16355
rect 5544 16295 5596 16355
rect 5634 16295 5686 16355
rect 5944 16295 5996 16355
rect 6034 16555 6086 16615
rect 6344 16555 6396 16615
rect 6434 16555 6486 16615
rect 6744 16555 6796 16615
rect 6834 16555 6886 16615
rect 7144 16555 7196 16615
rect 7234 16555 7286 16615
rect 7544 16555 7596 16615
rect 7634 16555 7686 16615
rect 7944 16555 7996 16615
rect 8034 16555 8086 16615
rect 8344 16555 8396 16615
rect 8434 16555 8486 16615
rect 8744 16555 8796 16615
rect 8834 16555 8886 16615
rect 9144 16555 9196 16615
rect 9234 16555 9286 16615
rect 9544 16555 9596 16615
rect 9634 16555 9686 16615
rect 9944 16555 9996 16615
rect 10034 16555 10086 16615
rect 10344 16555 10396 16615
rect 10434 16555 10486 16615
rect 10744 16555 10796 16615
rect 10834 16555 10886 16615
rect 11144 16555 11196 16615
rect 11234 16555 11286 16615
rect 11544 16555 11596 16615
rect 11634 16555 11686 16615
rect 11944 16555 11996 16615
rect 12034 16555 12086 16615
rect 12344 16555 12396 16615
rect 12434 16555 12486 16615
rect 12744 16555 12796 16615
rect 12834 16555 12886 16615
rect 13144 16555 13196 16615
rect 6034 16295 6086 16355
rect 6344 16295 6396 16355
rect 6434 16295 6486 16355
rect 6744 16295 6796 16355
rect 6834 16295 6886 16355
rect 7144 16295 7196 16355
rect 7234 16295 7286 16355
rect 7544 16295 7596 16355
rect 7634 16295 7686 16355
rect 7944 16295 7996 16355
rect 8034 16295 8086 16355
rect 8344 16295 8396 16355
rect 8434 16295 8486 16355
rect 8744 16295 8796 16355
rect 8834 16295 8886 16355
rect 9144 16295 9196 16355
rect 9234 16295 9286 16355
rect 9544 16295 9596 16355
rect 9634 16295 9686 16355
rect 9944 16295 9996 16355
rect 10034 16295 10086 16355
rect 10344 16295 10396 16355
rect 10434 16295 10486 16355
rect 10744 16295 10796 16355
rect 10834 16295 10886 16355
rect 11144 16295 11196 16355
rect 11234 16295 11286 16355
rect 11544 16295 11596 16355
rect 11634 16295 11686 16355
rect 11944 16295 11996 16355
rect 12034 16295 12086 16355
rect 12344 16295 12396 16355
rect 12434 16295 12486 16355
rect 12744 16295 12796 16355
rect 12834 16295 12886 16355
rect 13144 16295 13196 16355
rect -366 16185 -330 16245
rect -330 16185 -314 16245
rect -56 16185 -4 16245
rect -366 15925 -330 15985
rect -330 15925 -314 15985
rect -56 15925 -4 15985
rect 34 16185 86 16245
rect 344 16185 396 16245
rect 434 16185 486 16245
rect 744 16185 796 16245
rect 834 16185 886 16245
rect 1144 16185 1196 16245
rect 1234 16185 1286 16245
rect 1544 16185 1596 16245
rect 1634 16185 1686 16245
rect 1944 16185 1996 16245
rect 2034 16185 2086 16245
rect 2344 16185 2396 16245
rect 2434 16185 2486 16245
rect 2744 16185 2796 16245
rect 2834 16185 2886 16245
rect 3144 16185 3196 16245
rect 34 15925 86 15985
rect 344 15925 396 15985
rect 434 15925 486 15985
rect 744 15925 796 15985
rect 834 15925 886 15985
rect 1144 15925 1196 15985
rect 1234 15925 1286 15985
rect 1544 15925 1596 15985
rect 1634 15925 1686 15985
rect 1944 15925 1996 15985
rect 2034 15925 2086 15985
rect 2344 15925 2396 15985
rect 2434 15925 2486 15985
rect 2744 15925 2796 15985
rect 2834 15925 2886 15985
rect 3144 15925 3196 15985
rect 3234 16185 3286 16245
rect 3544 16185 3596 16245
rect 3634 16185 3686 16245
rect 3944 16185 3996 16245
rect 4034 16185 4086 16245
rect 4344 16185 4396 16245
rect 4434 16185 4486 16245
rect 4744 16185 4796 16245
rect 4834 16185 4886 16245
rect 5144 16185 5196 16245
rect 5234 16185 5286 16245
rect 5544 16185 5596 16245
rect 5634 16185 5686 16245
rect 5944 16185 5996 16245
rect 3234 15925 3286 15985
rect 3544 15925 3596 15985
rect 3634 15925 3686 15985
rect 3944 15925 3996 15985
rect 4034 15925 4086 15985
rect 4344 15925 4396 15985
rect 4434 15925 4486 15985
rect 4744 15925 4796 15985
rect 4834 15925 4886 15985
rect 5144 15925 5196 15985
rect 5234 15925 5286 15985
rect 5544 15925 5596 15985
rect 5634 15925 5686 15985
rect 5944 15925 5996 15985
rect 6034 16185 6086 16245
rect 6344 16185 6396 16245
rect 6434 16185 6486 16245
rect 6744 16185 6796 16245
rect 6834 16185 6886 16245
rect 7144 16185 7196 16245
rect 7234 16185 7286 16245
rect 7544 16185 7596 16245
rect 7634 16185 7686 16245
rect 7944 16185 7996 16245
rect 8034 16185 8086 16245
rect 8344 16185 8396 16245
rect 8434 16185 8486 16245
rect 8744 16185 8796 16245
rect 8834 16185 8886 16245
rect 9144 16185 9196 16245
rect 9234 16185 9286 16245
rect 9544 16185 9596 16245
rect 9634 16185 9686 16245
rect 9944 16185 9996 16245
rect 10034 16185 10086 16245
rect 10344 16185 10396 16245
rect 10434 16185 10486 16245
rect 10744 16185 10796 16245
rect 10834 16185 10886 16245
rect 11144 16185 11196 16245
rect 11234 16185 11286 16245
rect 11544 16185 11596 16245
rect 11634 16185 11686 16245
rect 11944 16185 11996 16245
rect 12034 16185 12086 16245
rect 12344 16185 12396 16245
rect 12434 16185 12486 16245
rect 12744 16185 12796 16245
rect 12834 16185 12886 16245
rect 13144 16185 13196 16245
rect 6034 15925 6086 15985
rect 6344 15925 6396 15985
rect 6434 15925 6486 15985
rect 6744 15925 6796 15985
rect 6834 15925 6886 15985
rect 7144 15925 7196 15985
rect 7234 15925 7286 15985
rect 7544 15925 7596 15985
rect 7634 15925 7686 15985
rect 7944 15925 7996 15985
rect 8034 15925 8086 15985
rect 8344 15925 8396 15985
rect 8434 15925 8486 15985
rect 8744 15925 8796 15985
rect 8834 15925 8886 15985
rect 9144 15925 9196 15985
rect 9234 15925 9286 15985
rect 9544 15925 9596 15985
rect 9634 15925 9686 15985
rect 9944 15925 9996 15985
rect 10034 15925 10086 15985
rect 10344 15925 10396 15985
rect 10434 15925 10486 15985
rect 10744 15925 10796 15985
rect 10834 15925 10886 15985
rect 11144 15925 11196 15985
rect 11234 15925 11286 15985
rect 11544 15925 11596 15985
rect 11634 15925 11686 15985
rect 11944 15925 11996 15985
rect 12034 15925 12086 15985
rect 12344 15925 12396 15985
rect 12434 15925 12486 15985
rect 12744 15925 12796 15985
rect 12834 15925 12886 15985
rect 13144 15925 13196 15985
rect -366 15815 -330 15875
rect -330 15815 -314 15875
rect -56 15815 -4 15875
rect -366 15555 -330 15615
rect -330 15555 -314 15615
rect -56 15555 -4 15615
rect 34 15815 86 15875
rect 344 15815 396 15875
rect 434 15815 486 15875
rect 744 15815 796 15875
rect 834 15815 886 15875
rect 1144 15815 1196 15875
rect 1234 15815 1286 15875
rect 1544 15815 1596 15875
rect 1634 15815 1686 15875
rect 1944 15815 1996 15875
rect 2034 15815 2086 15875
rect 2344 15815 2396 15875
rect 2434 15815 2486 15875
rect 2744 15815 2796 15875
rect 2834 15815 2886 15875
rect 3144 15815 3196 15875
rect 34 15555 86 15615
rect 344 15555 396 15615
rect 434 15555 486 15615
rect 744 15555 796 15615
rect 834 15555 886 15615
rect 1144 15555 1196 15615
rect 1234 15555 1286 15615
rect 1544 15555 1596 15615
rect 1634 15555 1686 15615
rect 1944 15555 1996 15615
rect 2034 15555 2086 15615
rect 2344 15555 2396 15615
rect 2434 15555 2486 15615
rect 2744 15555 2796 15615
rect 2834 15555 2886 15615
rect 3144 15555 3196 15615
rect 3234 15815 3286 15875
rect 3544 15815 3596 15875
rect 3634 15815 3686 15875
rect 3944 15815 3996 15875
rect 4034 15815 4086 15875
rect 4344 15815 4396 15875
rect 4434 15815 4486 15875
rect 4744 15815 4796 15875
rect 4834 15815 4886 15875
rect 5144 15815 5196 15875
rect 5234 15815 5286 15875
rect 5544 15815 5596 15875
rect 5634 15815 5686 15875
rect 5944 15815 5996 15875
rect 3234 15555 3286 15615
rect 3544 15555 3596 15615
rect 3634 15555 3686 15615
rect 3944 15555 3996 15615
rect 4034 15555 4086 15615
rect 4344 15555 4396 15615
rect 4434 15555 4486 15615
rect 4744 15555 4796 15615
rect 4834 15555 4886 15615
rect 5144 15555 5196 15615
rect 5234 15555 5286 15615
rect 5544 15555 5596 15615
rect 5634 15555 5686 15615
rect 5944 15555 5996 15615
rect 6034 15815 6086 15875
rect 6344 15815 6396 15875
rect 6434 15815 6486 15875
rect 6744 15815 6796 15875
rect 6834 15815 6886 15875
rect 7144 15815 7196 15875
rect 7234 15815 7286 15875
rect 7544 15815 7596 15875
rect 7634 15815 7686 15875
rect 7944 15815 7996 15875
rect 8034 15815 8086 15875
rect 8344 15815 8396 15875
rect 8434 15815 8486 15875
rect 8744 15815 8796 15875
rect 8834 15815 8886 15875
rect 9144 15815 9196 15875
rect 9234 15815 9286 15875
rect 9544 15815 9596 15875
rect 9634 15815 9686 15875
rect 9944 15815 9996 15875
rect 10034 15815 10086 15875
rect 10344 15815 10396 15875
rect 10434 15815 10486 15875
rect 10744 15815 10796 15875
rect 10834 15815 10886 15875
rect 11144 15815 11196 15875
rect 11234 15815 11286 15875
rect 11544 15815 11596 15875
rect 11634 15815 11686 15875
rect 11944 15815 11996 15875
rect 12034 15815 12086 15875
rect 12344 15815 12396 15875
rect 12434 15815 12486 15875
rect 12744 15815 12796 15875
rect 12834 15815 12886 15875
rect 13144 15815 13196 15875
rect 6034 15555 6086 15615
rect 6344 15555 6396 15615
rect 6434 15555 6486 15615
rect 6744 15555 6796 15615
rect 6834 15555 6886 15615
rect 7144 15555 7196 15615
rect 7234 15555 7286 15615
rect 7544 15555 7596 15615
rect 7634 15555 7686 15615
rect 7944 15555 7996 15615
rect 8034 15555 8086 15615
rect 8344 15555 8396 15615
rect 8434 15555 8486 15615
rect 8744 15555 8796 15615
rect 8834 15555 8886 15615
rect 9144 15555 9196 15615
rect 9234 15555 9286 15615
rect 9544 15555 9596 15615
rect 9634 15555 9686 15615
rect 9944 15555 9996 15615
rect 10034 15555 10086 15615
rect 10344 15555 10396 15615
rect 10434 15555 10486 15615
rect 10744 15555 10796 15615
rect 10834 15555 10886 15615
rect 11144 15555 11196 15615
rect 11234 15555 11286 15615
rect 11544 15555 11596 15615
rect 11634 15555 11686 15615
rect 11944 15555 11996 15615
rect 12034 15555 12086 15615
rect 12344 15555 12396 15615
rect 12434 15555 12486 15615
rect 12744 15555 12796 15615
rect 12834 15555 12886 15615
rect 13144 15555 13196 15615
rect -366 15445 -330 15505
rect -330 15445 -314 15505
rect -56 15445 -4 15505
rect -366 15185 -330 15245
rect -330 15185 -314 15245
rect -56 15185 -4 15245
rect 34 15445 86 15505
rect 344 15445 396 15505
rect 434 15445 486 15505
rect 744 15445 796 15505
rect 834 15445 886 15505
rect 1144 15445 1196 15505
rect 1234 15445 1286 15505
rect 1544 15445 1596 15505
rect 1634 15445 1686 15505
rect 1944 15445 1996 15505
rect 2034 15445 2086 15505
rect 2344 15445 2396 15505
rect 2434 15445 2486 15505
rect 2744 15445 2796 15505
rect 2834 15445 2886 15505
rect 3144 15445 3196 15505
rect 34 15185 86 15245
rect 344 15185 396 15245
rect 434 15185 486 15245
rect 744 15185 796 15245
rect 834 15185 886 15245
rect 1144 15185 1196 15245
rect 1234 15185 1286 15245
rect 1544 15185 1596 15245
rect 1634 15185 1686 15245
rect 1944 15185 1996 15245
rect 2034 15185 2086 15245
rect 2344 15185 2396 15245
rect 2434 15185 2486 15245
rect 2744 15185 2796 15245
rect 2834 15185 2886 15245
rect 3144 15185 3196 15245
rect 3234 15445 3286 15505
rect 3544 15445 3596 15505
rect 3634 15445 3686 15505
rect 3944 15445 3996 15505
rect 4034 15445 4086 15505
rect 4344 15445 4396 15505
rect 4434 15445 4486 15505
rect 4744 15445 4796 15505
rect 4834 15445 4886 15505
rect 5144 15445 5196 15505
rect 5234 15445 5286 15505
rect 5544 15445 5596 15505
rect 5634 15445 5686 15505
rect 5944 15445 5996 15505
rect 3234 15185 3286 15245
rect 3544 15185 3596 15245
rect 3634 15185 3686 15245
rect 3944 15185 3996 15245
rect 4034 15185 4086 15245
rect 4344 15185 4396 15245
rect 4434 15185 4486 15245
rect 4744 15185 4796 15245
rect 4834 15185 4886 15245
rect 5144 15185 5196 15245
rect 5234 15185 5286 15245
rect 5544 15185 5596 15245
rect 5634 15185 5686 15245
rect 5944 15185 5996 15245
rect 6034 15445 6086 15505
rect 6344 15445 6396 15505
rect 6434 15445 6486 15505
rect 6744 15445 6796 15505
rect 6834 15445 6886 15505
rect 7144 15445 7196 15505
rect 7234 15445 7286 15505
rect 7544 15445 7596 15505
rect 7634 15445 7686 15505
rect 7944 15445 7996 15505
rect 6034 15185 6086 15245
rect 6344 15185 6396 15245
rect 6434 15185 6486 15245
rect 6744 15185 6796 15245
rect 6834 15185 6886 15245
rect 7144 15185 7196 15245
rect 7234 15185 7286 15245
rect 7544 15185 7596 15245
rect 7634 15185 7686 15245
rect 7944 15185 7996 15245
rect 8034 15445 8086 15505
rect 8344 15445 8396 15505
rect 8434 15445 8486 15505
rect 8744 15445 8796 15505
rect 8834 15445 8886 15505
rect 9144 15445 9196 15505
rect 9234 15445 9286 15505
rect 9544 15445 9596 15505
rect 9634 15445 9686 15505
rect 9944 15445 9996 15505
rect 10034 15445 10086 15505
rect 10344 15445 10396 15505
rect 10434 15445 10486 15505
rect 10744 15445 10796 15505
rect 10834 15445 10886 15505
rect 11144 15445 11196 15505
rect 11234 15445 11286 15505
rect 11544 15445 11596 15505
rect 11634 15445 11686 15505
rect 11944 15445 11996 15505
rect 12034 15445 12086 15505
rect 12344 15445 12396 15505
rect 12434 15445 12486 15505
rect 12744 15445 12796 15505
rect 12834 15445 12886 15505
rect 13144 15445 13196 15505
rect 8034 15185 8086 15245
rect 8344 15185 8396 15245
rect 8434 15185 8486 15245
rect 8744 15185 8796 15245
rect 8834 15185 8886 15245
rect 9144 15185 9196 15245
rect 9234 15185 9286 15245
rect 9544 15185 9596 15245
rect 9634 15185 9686 15245
rect 9944 15185 9996 15245
rect 10034 15185 10086 15245
rect 10344 15185 10396 15245
rect 10434 15185 10486 15245
rect 10744 15185 10796 15245
rect 10834 15185 10886 15245
rect 11144 15185 11196 15245
rect 11234 15185 11286 15245
rect 11544 15185 11596 15245
rect 11634 15185 11686 15245
rect 11944 15185 11996 15245
rect 12034 15185 12086 15245
rect 12344 15185 12396 15245
rect 12434 15185 12486 15245
rect 12744 15185 12796 15245
rect 12834 15185 12886 15245
rect 13144 15185 13196 15245
rect -366 15075 -330 15135
rect -330 15075 -314 15135
rect -56 15075 -4 15135
rect -366 14815 -330 14875
rect -330 14815 -314 14875
rect -56 14815 -4 14875
rect 34 15075 86 15135
rect 344 15075 396 15135
rect 434 15075 486 15135
rect 744 15075 796 15135
rect 834 15075 886 15135
rect 1144 15075 1196 15135
rect 1234 15075 1286 15135
rect 1544 15075 1596 15135
rect 1634 15075 1686 15135
rect 1944 15075 1996 15135
rect 2034 15075 2086 15135
rect 2344 15075 2396 15135
rect 2434 15075 2486 15135
rect 2744 15075 2796 15135
rect 2834 15075 2886 15135
rect 3144 15075 3196 15135
rect 34 14815 86 14875
rect 344 14815 396 14875
rect 434 14815 486 14875
rect 744 14815 796 14875
rect 834 14815 886 14875
rect 1144 14815 1196 14875
rect 1234 14815 1286 14875
rect 1544 14815 1596 14875
rect 1634 14815 1686 14875
rect 1944 14815 1996 14875
rect 2034 14815 2086 14875
rect 2344 14815 2396 14875
rect 2434 14815 2486 14875
rect 2744 14815 2796 14875
rect 2834 14815 2886 14875
rect 3144 14815 3196 14875
rect 3234 15075 3286 15135
rect 3544 15075 3596 15135
rect 3634 15075 3686 15135
rect 3944 15075 3996 15135
rect 4034 15075 4086 15135
rect 4344 15075 4396 15135
rect 4434 15075 4486 15135
rect 4744 15075 4796 15135
rect 4834 15075 4886 15135
rect 5144 15075 5196 15135
rect 5234 15075 5286 15135
rect 5544 15075 5596 15135
rect 5634 15075 5686 15135
rect 5944 15075 5996 15135
rect 3234 14815 3286 14875
rect 3544 14815 3596 14875
rect 3634 14815 3686 14875
rect 3944 14815 3996 14875
rect 4034 14815 4086 14875
rect 4344 14815 4396 14875
rect 4434 14815 4486 14875
rect 4744 14815 4796 14875
rect 4834 14815 4886 14875
rect 5144 14815 5196 14875
rect 5234 14815 5286 14875
rect 5544 14815 5596 14875
rect 5634 14815 5686 14875
rect 5944 14815 5996 14875
rect 6034 15075 6086 15135
rect 6344 15075 6396 15135
rect 6434 15075 6486 15135
rect 6744 15075 6796 15135
rect 6834 15075 6886 15135
rect 7144 15075 7196 15135
rect 7234 15075 7286 15135
rect 7544 15075 7596 15135
rect 7634 15075 7686 15135
rect 7944 15075 7996 15135
rect 6034 14815 6086 14875
rect 6344 14815 6396 14875
rect 6434 14815 6486 14875
rect 6744 14815 6796 14875
rect 6834 14815 6886 14875
rect 7144 14815 7196 14875
rect 7234 14815 7286 14875
rect 7544 14815 7596 14875
rect 7634 14815 7686 14875
rect 7944 14815 7996 14875
rect 8034 15075 8086 15135
rect 8344 15075 8396 15135
rect 8434 15075 8486 15135
rect 8744 15075 8796 15135
rect 8834 15075 8886 15135
rect 9144 15075 9196 15135
rect 9234 15075 9286 15135
rect 9544 15075 9596 15135
rect 9634 15075 9686 15135
rect 9944 15075 9996 15135
rect 10034 15075 10086 15135
rect 10344 15075 10396 15135
rect 10434 15075 10486 15135
rect 10744 15075 10796 15135
rect 10834 15075 10886 15135
rect 11144 15075 11196 15135
rect 11234 15075 11286 15135
rect 11544 15075 11596 15135
rect 11634 15075 11686 15135
rect 11944 15075 11996 15135
rect 12034 15075 12086 15135
rect 12344 15075 12396 15135
rect 12434 15075 12486 15135
rect 12744 15075 12796 15135
rect 12834 15075 12886 15135
rect 13144 15075 13196 15135
rect 8034 14815 8086 14875
rect 8344 14815 8396 14875
rect 8434 14815 8486 14875
rect 8744 14815 8796 14875
rect 8834 14815 8886 14875
rect 9144 14815 9196 14875
rect 9234 14815 9286 14875
rect 9544 14815 9596 14875
rect 9634 14815 9686 14875
rect 9944 14815 9996 14875
rect 10034 14815 10086 14875
rect 10344 14815 10396 14875
rect 10434 14815 10486 14875
rect 10744 14815 10796 14875
rect 10834 14815 10886 14875
rect 11144 14815 11196 14875
rect 11234 14815 11286 14875
rect 11544 14815 11596 14875
rect 11634 14815 11686 14875
rect 11944 14815 11996 14875
rect 12034 14815 12086 14875
rect 12344 14815 12396 14875
rect 12434 14815 12486 14875
rect 12744 14815 12796 14875
rect 12834 14815 12886 14875
rect 13144 14815 13196 14875
rect -366 14705 -330 14765
rect -330 14705 -314 14765
rect -56 14705 -4 14765
rect -366 14445 -330 14505
rect -330 14445 -314 14505
rect -56 14445 -4 14505
rect 34 14705 86 14765
rect 344 14705 396 14765
rect 434 14705 486 14765
rect 744 14705 796 14765
rect 834 14705 886 14765
rect 1144 14705 1196 14765
rect 1234 14705 1286 14765
rect 1544 14705 1596 14765
rect 1634 14705 1686 14765
rect 1944 14705 1996 14765
rect 2034 14705 2086 14765
rect 2344 14705 2396 14765
rect 2434 14705 2486 14765
rect 2744 14705 2796 14765
rect 34 14445 86 14505
rect 344 14445 396 14505
rect 434 14445 486 14505
rect 744 14445 796 14505
rect 834 14445 886 14505
rect 1144 14445 1196 14505
rect 1234 14445 1286 14505
rect 1544 14445 1596 14505
rect 1634 14445 1686 14505
rect 1944 14445 1996 14505
rect 2034 14445 2086 14505
rect 2344 14445 2396 14505
rect 2434 14445 2486 14505
rect 2744 14445 2796 14505
rect 2834 14705 2886 14765
rect 3144 14705 3196 14765
rect 3234 14705 3286 14765
rect 3544 14705 3596 14765
rect 3634 14705 3686 14765
rect 3944 14705 3996 14765
rect 4034 14705 4086 14765
rect 4344 14705 4396 14765
rect 4434 14705 4486 14765
rect 4744 14705 4796 14765
rect 4834 14705 4886 14765
rect 5144 14705 5196 14765
rect 5234 14705 5286 14765
rect 5544 14705 5596 14765
rect 5634 14705 5686 14765
rect 5944 14705 5996 14765
rect 2834 14445 2886 14505
rect 3144 14445 3196 14505
rect 3234 14445 3286 14505
rect 3544 14445 3596 14505
rect 3634 14445 3686 14505
rect 3944 14445 3996 14505
rect 4034 14445 4086 14505
rect 4344 14445 4396 14505
rect 4434 14445 4486 14505
rect 4744 14445 4796 14505
rect 4834 14445 4886 14505
rect 5144 14445 5196 14505
rect 5234 14445 5286 14505
rect 5544 14445 5596 14505
rect 5634 14445 5686 14505
rect 5944 14445 5996 14505
rect 6034 14705 6086 14765
rect 6344 14705 6396 14765
rect 6434 14705 6486 14765
rect 6744 14705 6796 14765
rect 6834 14705 6886 14765
rect 7144 14705 7196 14765
rect 7234 14705 7286 14765
rect 7544 14705 7596 14765
rect 6034 14445 6086 14505
rect 6344 14445 6396 14505
rect 6434 14445 6486 14505
rect 6744 14445 6796 14505
rect 6834 14445 6886 14505
rect 7144 14445 7196 14505
rect 7234 14445 7286 14505
rect 7544 14445 7596 14505
rect 7634 14705 7686 14765
rect 7944 14705 7996 14765
rect 8034 14705 8086 14765
rect 8344 14705 8396 14765
rect 8434 14705 8486 14765
rect 8744 14705 8796 14765
rect 8834 14705 8886 14765
rect 9144 14705 9196 14765
rect 9234 14705 9286 14765
rect 9544 14705 9596 14765
rect 9634 14705 9686 14765
rect 9944 14705 9996 14765
rect 10034 14705 10086 14765
rect 10344 14705 10396 14765
rect 10434 14705 10486 14765
rect 10744 14705 10796 14765
rect 10834 14705 10886 14765
rect 11144 14705 11196 14765
rect 11234 14705 11286 14765
rect 11544 14705 11596 14765
rect 11634 14705 11686 14765
rect 11944 14705 11996 14765
rect 12034 14705 12086 14765
rect 12344 14705 12396 14765
rect 12434 14705 12486 14765
rect 12744 14705 12796 14765
rect 12834 14705 12886 14765
rect 13144 14705 13196 14765
rect 7634 14445 7686 14505
rect 7944 14445 7996 14505
rect 8034 14445 8086 14505
rect 8344 14445 8396 14505
rect 8434 14445 8486 14505
rect 8744 14445 8796 14505
rect 8834 14445 8886 14505
rect 9144 14445 9196 14505
rect 9234 14445 9286 14505
rect 9544 14445 9596 14505
rect 9634 14445 9686 14505
rect 9944 14445 9996 14505
rect 10034 14445 10086 14505
rect 10344 14445 10396 14505
rect 10434 14445 10486 14505
rect 10744 14445 10796 14505
rect 10834 14445 10886 14505
rect 11144 14445 11196 14505
rect 11234 14445 11286 14505
rect 11544 14445 11596 14505
rect 11634 14445 11686 14505
rect 11944 14445 11996 14505
rect 12034 14445 12086 14505
rect 12344 14445 12396 14505
rect 12434 14445 12486 14505
rect 12744 14445 12796 14505
rect 12834 14445 12886 14505
rect 13144 14445 13196 14505
rect -366 14335 -330 14395
rect -330 14335 -314 14395
rect -56 14335 -4 14395
rect -366 14075 -330 14135
rect -330 14075 -314 14135
rect -56 14075 -4 14135
rect 34 14335 86 14395
rect 344 14335 396 14395
rect 434 14335 486 14395
rect 744 14335 796 14395
rect 834 14335 886 14395
rect 1144 14335 1196 14395
rect 1234 14335 1286 14395
rect 1544 14335 1596 14395
rect 1634 14335 1686 14395
rect 1944 14335 1996 14395
rect 2034 14335 2086 14395
rect 2344 14335 2396 14395
rect 2434 14335 2486 14395
rect 2744 14335 2796 14395
rect 34 14075 86 14135
rect 344 14075 396 14135
rect 434 14075 486 14135
rect 744 14075 796 14135
rect 834 14075 886 14135
rect 1144 14075 1196 14135
rect 1234 14075 1286 14135
rect 1544 14075 1596 14135
rect 1634 14075 1686 14135
rect 1944 14075 1996 14135
rect 2034 14075 2086 14135
rect 2344 14075 2396 14135
rect 2434 14075 2486 14135
rect 2744 14075 2796 14135
rect 2834 14335 2886 14395
rect 3144 14335 3196 14395
rect 3234 14335 3286 14395
rect 3544 14335 3596 14395
rect 3634 14335 3686 14395
rect 3944 14335 3996 14395
rect 4034 14335 4086 14395
rect 4344 14335 4396 14395
rect 4434 14335 4486 14395
rect 4744 14335 4796 14395
rect 4834 14335 4886 14395
rect 5144 14335 5196 14395
rect 5234 14335 5286 14395
rect 5544 14335 5596 14395
rect 5634 14335 5686 14395
rect 5944 14335 5996 14395
rect 2834 14075 2886 14135
rect 3144 14075 3196 14135
rect 3234 14075 3286 14135
rect 3544 14075 3596 14135
rect 3634 14075 3686 14135
rect 3944 14075 3996 14135
rect 4034 14075 4086 14135
rect 4344 14075 4396 14135
rect 4434 14075 4486 14135
rect 4744 14075 4796 14135
rect 4834 14075 4886 14135
rect 5144 14075 5196 14135
rect 5234 14075 5286 14135
rect 5544 14075 5596 14135
rect 5634 14075 5686 14135
rect 5944 14075 5996 14135
rect 6034 14335 6086 14395
rect 6344 14335 6396 14395
rect 6434 14335 6486 14395
rect 6744 14335 6796 14395
rect 6834 14335 6886 14395
rect 7144 14335 7196 14395
rect 7234 14335 7286 14395
rect 7544 14335 7596 14395
rect 6034 14075 6086 14135
rect 6344 14075 6396 14135
rect 6434 14075 6486 14135
rect 6744 14075 6796 14135
rect 6834 14075 6886 14135
rect 7144 14075 7196 14135
rect 7234 14075 7286 14135
rect 7544 14075 7596 14135
rect 7634 14335 7686 14395
rect 7944 14335 7996 14395
rect 8034 14335 8086 14395
rect 8344 14335 8396 14395
rect 7634 14075 7686 14135
rect 7944 14075 7996 14135
rect 8034 14075 8086 14135
rect 8344 14075 8396 14135
rect 8434 14335 8486 14395
rect 8744 14335 8796 14395
rect 8434 14075 8486 14135
rect 8744 14075 8796 14135
rect 8834 14335 8886 14395
rect 9144 14335 9196 14395
rect 8834 14075 8886 14135
rect 9144 14075 9196 14135
rect 9234 14335 9286 14395
rect 9544 14335 9596 14395
rect 9634 14335 9686 14395
rect 9944 14335 9996 14395
rect 10034 14335 10086 14395
rect 10344 14335 10396 14395
rect 10434 14335 10486 14395
rect 10744 14335 10796 14395
rect 10834 14335 10886 14395
rect 11144 14335 11196 14395
rect 11234 14335 11286 14395
rect 11544 14335 11596 14395
rect 11634 14335 11686 14395
rect 11944 14335 11996 14395
rect 12034 14335 12086 14395
rect 12344 14335 12396 14395
rect 12434 14335 12486 14395
rect 12744 14335 12796 14395
rect 12834 14335 12886 14395
rect 13144 14335 13196 14395
rect 9234 14075 9286 14135
rect 9544 14075 9596 14135
rect 9634 14075 9686 14135
rect 9944 14075 9996 14135
rect 10034 14075 10086 14135
rect 10344 14075 10396 14135
rect 10434 14075 10486 14135
rect 10744 14075 10796 14135
rect 10834 14075 10886 14135
rect 11144 14075 11196 14135
rect 11234 14075 11286 14135
rect 11544 14075 11596 14135
rect 11634 14075 11686 14135
rect 11944 14075 11996 14135
rect 12034 14075 12086 14135
rect 12344 14075 12396 14135
rect 12434 14075 12486 14135
rect 12744 14075 12796 14135
rect 12834 14075 12886 14135
rect 13144 14075 13196 14135
rect -366 13965 -330 14025
rect -330 13965 -314 14025
rect -56 13965 -4 14025
rect -366 13705 -330 13765
rect -330 13705 -314 13765
rect -56 13705 -4 13765
rect 34 13965 86 14025
rect 344 13965 396 14025
rect 434 13965 486 14025
rect 744 13965 796 14025
rect 834 13965 886 14025
rect 1144 13965 1196 14025
rect 1234 13965 1286 14025
rect 1544 13965 1596 14025
rect 1634 13965 1686 14025
rect 1944 13965 1996 14025
rect 2034 13965 2086 14025
rect 2344 13965 2396 14025
rect 2434 13965 2486 14025
rect 2744 13965 2796 14025
rect 34 13705 86 13765
rect 344 13705 396 13765
rect 434 13705 486 13765
rect 744 13705 796 13765
rect 834 13705 886 13765
rect 1144 13705 1196 13765
rect 1234 13705 1286 13765
rect 1544 13705 1596 13765
rect 1634 13705 1686 13765
rect 1944 13705 1996 13765
rect 2034 13705 2086 13765
rect 2344 13705 2396 13765
rect 2434 13705 2486 13765
rect 2744 13705 2796 13765
rect 2834 13965 2886 14025
rect 3144 13965 3196 14025
rect 3234 13965 3286 14025
rect 3544 13965 3596 14025
rect 3634 13965 3686 14025
rect 3944 13965 3996 14025
rect 4034 13965 4086 14025
rect 4344 13965 4396 14025
rect 4434 13965 4486 14025
rect 4744 13965 4796 14025
rect 4834 13965 4886 14025
rect 5144 13965 5196 14025
rect 5234 13965 5286 14025
rect 5544 13965 5596 14025
rect 5634 13965 5686 14025
rect 5944 13965 5996 14025
rect 2834 13705 2886 13765
rect 3144 13705 3196 13765
rect 3234 13705 3286 13765
rect 3544 13705 3596 13765
rect 3634 13705 3686 13765
rect 3944 13705 3996 13765
rect 4034 13705 4086 13765
rect 4344 13705 4396 13765
rect 4434 13705 4486 13765
rect 4744 13705 4796 13765
rect 4834 13705 4886 13765
rect 5144 13705 5196 13765
rect 5234 13705 5286 13765
rect 5544 13705 5596 13765
rect 5634 13705 5686 13765
rect 5944 13705 5996 13765
rect 6034 13965 6086 14025
rect 6344 13965 6396 14025
rect 6434 13965 6486 14025
rect 6744 13965 6796 14025
rect 6834 13965 6886 14025
rect 7144 13965 7196 14025
rect 7234 13965 7286 14025
rect 7544 13965 7596 14025
rect 6034 13705 6086 13765
rect 6344 13705 6396 13765
rect 6434 13705 6486 13765
rect 6744 13705 6796 13765
rect 6834 13705 6886 13765
rect 7144 13705 7196 13765
rect 7234 13705 7286 13765
rect 7544 13705 7596 13765
rect 7634 13965 7686 14025
rect 7944 13965 7996 14025
rect 8034 13965 8086 14025
rect 8344 13965 8396 14025
rect 7634 13705 7686 13765
rect 7944 13705 7996 13765
rect 8034 13705 8086 13765
rect 8344 13705 8396 13765
rect 8434 13965 8486 14025
rect 8744 13965 8796 14025
rect 8434 13705 8486 13765
rect 8744 13705 8796 13765
rect 8834 13965 8886 14025
rect 9144 13965 9196 14025
rect 8834 13705 8886 13765
rect 9144 13705 9196 13765
rect 9234 13965 9286 14025
rect 9544 13965 9596 14025
rect 9634 13965 9686 14025
rect 9944 13965 9996 14025
rect 10034 13965 10086 14025
rect 10344 13965 10396 14025
rect 10434 13965 10486 14025
rect 10744 13965 10796 14025
rect 10834 13965 10886 14025
rect 11144 13965 11196 14025
rect 11234 13965 11286 14025
rect 11544 13965 11596 14025
rect 11634 13965 11686 14025
rect 11944 13965 11996 14025
rect 12034 13965 12086 14025
rect 12344 13965 12396 14025
rect 12434 13965 12486 14025
rect 12744 13965 12796 14025
rect 12834 13965 12886 14025
rect 13144 13965 13196 14025
rect 9234 13705 9286 13765
rect 9544 13705 9596 13765
rect 9634 13705 9686 13765
rect 9944 13705 9996 13765
rect 10034 13705 10086 13765
rect 10344 13705 10396 13765
rect 10434 13705 10486 13765
rect 10744 13705 10796 13765
rect 10834 13705 10886 13765
rect 11144 13705 11196 13765
rect 11234 13705 11286 13765
rect 11544 13705 11596 13765
rect 11634 13705 11686 13765
rect 11944 13705 11996 13765
rect 12034 13705 12086 13765
rect 12344 13705 12396 13765
rect 12434 13705 12486 13765
rect 12744 13705 12796 13765
rect 12834 13705 12886 13765
rect 13144 13705 13196 13765
rect -366 13595 -330 13655
rect -330 13595 -314 13655
rect -56 13595 -4 13655
rect -366 13335 -330 13395
rect -330 13335 -314 13395
rect -56 13335 -4 13395
rect 34 13595 86 13655
rect 344 13595 396 13655
rect 434 13595 486 13655
rect 744 13595 796 13655
rect 834 13595 886 13655
rect 1144 13595 1196 13655
rect 1234 13595 1286 13655
rect 1544 13595 1596 13655
rect 1634 13595 1686 13655
rect 1944 13595 1996 13655
rect 2034 13595 2086 13655
rect 2344 13595 2396 13655
rect 2434 13595 2486 13655
rect 2744 13595 2796 13655
rect 34 13335 86 13395
rect 344 13335 396 13395
rect 434 13335 486 13395
rect 744 13335 796 13395
rect 834 13335 886 13395
rect 1144 13335 1196 13395
rect 1234 13335 1286 13395
rect 1544 13335 1596 13395
rect 1634 13335 1686 13395
rect 1944 13335 1996 13395
rect 2034 13335 2086 13395
rect 2344 13335 2396 13395
rect 2434 13335 2486 13395
rect 2744 13335 2796 13395
rect 2834 13595 2886 13655
rect 3144 13595 3196 13655
rect 3234 13595 3286 13655
rect 3544 13595 3596 13655
rect 3634 13595 3686 13655
rect 3944 13595 3996 13655
rect 4034 13595 4086 13655
rect 4344 13595 4396 13655
rect 4434 13595 4486 13655
rect 4744 13595 4796 13655
rect 4834 13595 4886 13655
rect 5144 13595 5196 13655
rect 5234 13595 5286 13655
rect 5544 13595 5596 13655
rect 5634 13595 5686 13655
rect 5944 13595 5996 13655
rect 2834 13335 2886 13395
rect 3144 13335 3196 13395
rect 3234 13335 3286 13395
rect 3544 13335 3596 13395
rect 3634 13335 3686 13395
rect 3944 13335 3996 13395
rect 4034 13335 4086 13395
rect 4344 13335 4396 13395
rect 4434 13335 4486 13395
rect 4744 13335 4796 13395
rect 4834 13335 4886 13395
rect 5144 13335 5196 13395
rect 5234 13335 5286 13395
rect 5544 13335 5596 13395
rect 5634 13335 5686 13395
rect 5944 13335 5996 13395
rect 6034 13595 6086 13655
rect 6344 13595 6396 13655
rect 6434 13595 6486 13655
rect 6744 13595 6796 13655
rect 6834 13595 6886 13655
rect 7144 13595 7196 13655
rect 7234 13595 7286 13655
rect 7544 13595 7596 13655
rect 6034 13335 6086 13395
rect 6344 13335 6396 13395
rect 6434 13335 6486 13395
rect 6744 13335 6796 13395
rect 6834 13335 6886 13395
rect 7144 13335 7196 13395
rect 7234 13335 7286 13395
rect 7544 13335 7596 13395
rect 7634 13595 7686 13655
rect 7944 13595 7996 13655
rect 8034 13595 8086 13655
rect 8344 13595 8396 13655
rect 7634 13335 7686 13395
rect 7944 13335 7996 13395
rect 8034 13335 8086 13395
rect 8344 13335 8396 13395
rect 8434 13595 8486 13655
rect 8744 13595 8796 13655
rect 8434 13335 8486 13395
rect 8744 13335 8796 13395
rect 8834 13595 8886 13655
rect 9144 13595 9196 13655
rect 8834 13335 8886 13395
rect 9144 13335 9196 13395
rect 9234 13595 9286 13655
rect 9544 13595 9596 13655
rect 9634 13595 9686 13655
rect 9944 13595 9996 13655
rect 10034 13595 10086 13655
rect 10344 13595 10396 13655
rect 9234 13335 9286 13395
rect 9544 13335 9596 13395
rect 9634 13335 9686 13395
rect 9944 13335 9996 13395
rect 10034 13335 10086 13395
rect 10344 13335 10396 13395
rect 10434 13595 10486 13655
rect 10744 13595 10796 13655
rect 10834 13595 10886 13655
rect 11144 13595 11196 13655
rect 11234 13595 11286 13655
rect 11544 13595 11596 13655
rect 11634 13595 11686 13655
rect 11944 13595 11996 13655
rect 12034 13595 12086 13655
rect 12344 13595 12396 13655
rect 12434 13595 12486 13655
rect 12744 13595 12796 13655
rect 12834 13595 12886 13655
rect 13144 13595 13196 13655
rect 10434 13335 10486 13395
rect 10744 13335 10796 13395
rect 10834 13335 10886 13395
rect 11144 13335 11196 13395
rect 11234 13335 11286 13395
rect 11544 13335 11596 13395
rect 11634 13335 11686 13395
rect 11944 13335 11996 13395
rect 12034 13335 12086 13395
rect 12344 13335 12396 13395
rect 12434 13335 12486 13395
rect 12744 13335 12796 13395
rect 12834 13335 12886 13395
rect 13144 13335 13196 13395
rect -366 13225 -330 13285
rect -330 13225 -314 13285
rect -56 13225 -4 13285
rect -366 12965 -330 13025
rect -330 12965 -314 13025
rect -56 12965 -4 13025
rect 34 13225 86 13285
rect 344 13225 396 13285
rect 434 13225 486 13285
rect 744 13225 796 13285
rect 834 13225 886 13285
rect 1144 13225 1196 13285
rect 1234 13225 1286 13285
rect 1544 13225 1596 13285
rect 1634 13225 1686 13285
rect 1944 13225 1996 13285
rect 2034 13225 2086 13285
rect 2344 13225 2396 13285
rect 2434 13225 2486 13285
rect 2744 13225 2796 13285
rect 34 12965 86 13025
rect 344 12965 396 13025
rect 434 12965 486 13025
rect 744 12965 796 13025
rect 834 12965 886 13025
rect 1144 12965 1196 13025
rect 1234 12965 1286 13025
rect 1544 12965 1596 13025
rect 1634 12965 1686 13025
rect 1944 12965 1996 13025
rect 2034 12965 2086 13025
rect 2344 12965 2396 13025
rect 2434 12965 2486 13025
rect 2744 12965 2796 13025
rect 2834 13225 2886 13285
rect 3144 13225 3196 13285
rect 3234 13225 3286 13285
rect 3544 13225 3596 13285
rect 3634 13225 3686 13285
rect 3944 13225 3996 13285
rect 4034 13225 4086 13285
rect 4344 13225 4396 13285
rect 4434 13225 4486 13285
rect 4744 13225 4796 13285
rect 4834 13225 4886 13285
rect 5144 13225 5196 13285
rect 5234 13225 5286 13285
rect 5544 13225 5596 13285
rect 5634 13225 5686 13285
rect 5944 13225 5996 13285
rect 2834 12965 2886 13025
rect 3144 12965 3196 13025
rect 3234 12965 3286 13025
rect 3544 12965 3596 13025
rect 3634 12965 3686 13025
rect 3944 12965 3996 13025
rect 4034 12965 4086 13025
rect 4344 12965 4396 13025
rect 4434 12965 4486 13025
rect 4744 12965 4796 13025
rect 4834 12965 4886 13025
rect 5144 12965 5196 13025
rect 5234 12965 5286 13025
rect 5544 12965 5596 13025
rect 5634 12965 5686 13025
rect 5944 12965 5996 13025
rect 6034 13225 6086 13285
rect 6344 13225 6396 13285
rect 6434 13225 6486 13285
rect 6744 13225 6796 13285
rect 6834 13225 6886 13285
rect 7144 13225 7196 13285
rect 7234 13225 7286 13285
rect 7544 13225 7596 13285
rect 6034 12965 6086 13025
rect 6344 12965 6396 13025
rect 6434 12965 6486 13025
rect 6744 12965 6796 13025
rect 6834 12965 6886 13025
rect 7144 12965 7196 13025
rect 7234 12965 7286 13025
rect 7544 12965 7596 13025
rect 7634 13225 7686 13285
rect 7944 13225 7996 13285
rect 8034 13225 8086 13285
rect 8344 13225 8396 13285
rect 7634 12965 7686 13025
rect 7944 12965 7996 13025
rect 8034 12965 8086 13025
rect 8344 12965 8396 13025
rect 8434 13225 8486 13285
rect 8744 13225 8796 13285
rect 8434 12965 8486 13025
rect 8744 12965 8796 13025
rect 8834 13225 8886 13285
rect 9144 13225 9196 13285
rect 8834 12965 8886 13025
rect 9144 12965 9196 13025
rect 9234 13225 9286 13285
rect 9544 13225 9596 13285
rect 9634 13225 9686 13285
rect 9944 13225 9996 13285
rect 10034 13225 10086 13285
rect 10344 13225 10396 13285
rect 9234 12965 9286 13025
rect 9544 12965 9596 13025
rect 9634 12965 9686 13025
rect 9944 12965 9996 13025
rect 10034 12965 10086 13025
rect 10344 12965 10396 13025
rect 10434 13225 10486 13285
rect 10744 13225 10796 13285
rect 10834 13225 10886 13285
rect 11144 13225 11196 13285
rect 10434 12965 10486 13025
rect 10744 12965 10796 13025
rect 10834 12965 10886 13025
rect 11144 12965 11196 13025
rect 11234 13225 11286 13285
rect 11544 13225 11596 13285
rect 11634 13225 11686 13285
rect 11944 13225 11996 13285
rect 12034 13225 12086 13285
rect 12344 13225 12396 13285
rect 12434 13225 12486 13285
rect 12744 13225 12796 13285
rect 12834 13225 12886 13285
rect 13144 13225 13196 13285
rect 11234 12965 11286 13025
rect 11544 12965 11596 13025
rect 11634 12965 11686 13025
rect 11944 12965 11996 13025
rect 12034 12965 12086 13025
rect 12344 12965 12396 13025
rect 12434 12965 12486 13025
rect 12744 12965 12796 13025
rect 12834 12965 12886 13025
rect 13144 12965 13196 13025
rect -366 12855 -330 12915
rect -330 12855 -314 12915
rect -56 12855 -4 12915
rect -366 12595 -330 12655
rect -330 12595 -314 12655
rect -56 12595 -4 12655
rect 34 12855 86 12915
rect 344 12855 396 12915
rect 434 12855 486 12915
rect 744 12855 796 12915
rect 834 12855 886 12915
rect 1144 12855 1196 12915
rect 1234 12855 1286 12915
rect 1544 12855 1596 12915
rect 1634 12855 1686 12915
rect 1944 12855 1996 12915
rect 2034 12855 2086 12915
rect 2344 12855 2396 12915
rect 2434 12855 2486 12915
rect 2744 12855 2796 12915
rect 34 12595 86 12655
rect 344 12595 396 12655
rect 434 12595 486 12655
rect 744 12595 796 12655
rect 834 12595 886 12655
rect 1144 12595 1196 12655
rect 1234 12595 1286 12655
rect 1544 12595 1596 12655
rect 1634 12595 1686 12655
rect 1944 12595 1996 12655
rect 2034 12595 2086 12655
rect 2344 12595 2396 12655
rect 2434 12595 2486 12655
rect 2744 12595 2796 12655
rect 2834 12855 2886 12915
rect 3144 12855 3196 12915
rect 3234 12855 3286 12915
rect 3544 12855 3596 12915
rect 3634 12855 3686 12915
rect 3944 12855 3996 12915
rect 4034 12855 4086 12915
rect 4344 12855 4396 12915
rect 4434 12855 4486 12915
rect 4744 12855 4796 12915
rect 4834 12855 4886 12915
rect 5144 12855 5196 12915
rect 5234 12855 5286 12915
rect 5544 12855 5596 12915
rect 5634 12855 5686 12915
rect 5944 12855 5996 12915
rect 2834 12595 2886 12655
rect 3144 12595 3196 12655
rect 3234 12595 3286 12655
rect 3544 12595 3596 12655
rect 3634 12595 3686 12655
rect 3944 12595 3996 12655
rect 4034 12595 4086 12655
rect 4344 12595 4396 12655
rect 4434 12595 4486 12655
rect 4744 12595 4796 12655
rect 4834 12595 4886 12655
rect 5144 12595 5196 12655
rect 5234 12595 5286 12655
rect 5544 12595 5596 12655
rect 5634 12595 5686 12655
rect 5944 12595 5996 12655
rect 6034 12855 6086 12915
rect 6344 12855 6396 12915
rect 6434 12855 6486 12915
rect 6744 12855 6796 12915
rect 6834 12855 6886 12915
rect 7144 12855 7196 12915
rect 7234 12855 7286 12915
rect 7544 12855 7596 12915
rect 6034 12595 6086 12655
rect 6344 12595 6396 12655
rect 6434 12595 6486 12655
rect 6744 12595 6796 12655
rect 6834 12595 6886 12655
rect 7144 12595 7196 12655
rect 7234 12595 7286 12655
rect 7544 12595 7596 12655
rect 7634 12855 7686 12915
rect 7944 12855 7996 12915
rect 8034 12855 8086 12915
rect 8344 12855 8396 12915
rect 7634 12595 7686 12655
rect 7944 12595 7996 12655
rect 8034 12595 8086 12655
rect 8344 12595 8396 12655
rect 8434 12855 8486 12915
rect 8744 12855 8796 12915
rect 8434 12595 8486 12655
rect 8744 12595 8796 12655
rect 8834 12855 8886 12915
rect 9144 12855 9196 12915
rect 8834 12595 8886 12655
rect 9144 12595 9196 12655
rect 9234 12855 9286 12915
rect 9544 12855 9596 12915
rect 9634 12855 9686 12915
rect 9944 12855 9996 12915
rect 10034 12855 10086 12915
rect 10344 12855 10396 12915
rect 9234 12595 9286 12655
rect 9544 12595 9596 12655
rect 9634 12595 9686 12655
rect 9944 12595 9996 12655
rect 10034 12595 10086 12655
rect 10344 12595 10396 12655
rect 10434 12855 10486 12915
rect 10744 12855 10796 12915
rect 10834 12855 10886 12915
rect 11144 12855 11196 12915
rect 10434 12595 10486 12655
rect 10744 12595 10796 12655
rect 10834 12595 10886 12655
rect 11144 12595 11196 12655
rect 11234 12855 11286 12915
rect 11544 12855 11596 12915
rect 11234 12595 11286 12655
rect 11544 12595 11596 12655
rect 11634 12855 11686 12915
rect 11944 12855 11996 12915
rect 12034 12855 12086 12915
rect 12344 12855 12396 12915
rect 12434 12855 12486 12915
rect 12744 12855 12796 12915
rect 12834 12855 12886 12915
rect 13144 12855 13196 12915
rect 11634 12595 11686 12655
rect 11944 12595 11996 12655
rect 12034 12595 12086 12655
rect 12344 12595 12396 12655
rect 12434 12595 12486 12655
rect 12744 12595 12796 12655
rect 12834 12595 12886 12655
rect 13144 12595 13196 12655
rect -366 12485 -330 12545
rect -330 12485 -314 12545
rect -56 12485 -4 12545
rect -366 12225 -330 12285
rect -330 12225 -314 12285
rect -56 12225 -4 12285
rect 34 12485 86 12545
rect 344 12485 396 12545
rect 434 12485 486 12545
rect 744 12485 796 12545
rect 834 12485 886 12545
rect 1144 12485 1196 12545
rect 1234 12485 1286 12545
rect 1544 12485 1596 12545
rect 1634 12485 1686 12545
rect 1944 12485 1996 12545
rect 2034 12485 2086 12545
rect 2344 12485 2396 12545
rect 2434 12485 2486 12545
rect 2744 12485 2796 12545
rect 34 12225 86 12285
rect 344 12225 396 12285
rect 434 12225 486 12285
rect 744 12225 796 12285
rect 834 12225 886 12285
rect 1144 12225 1196 12285
rect 1234 12225 1286 12285
rect 1544 12225 1596 12285
rect 1634 12225 1686 12285
rect 1944 12225 1996 12285
rect 2034 12225 2086 12285
rect 2344 12225 2396 12285
rect 2434 12225 2486 12285
rect 2744 12225 2796 12285
rect 2834 12485 2886 12545
rect 3144 12485 3196 12545
rect 3234 12485 3286 12545
rect 3544 12485 3596 12545
rect 3634 12485 3686 12545
rect 3944 12485 3996 12545
rect 4034 12485 4086 12545
rect 4344 12485 4396 12545
rect 4434 12485 4486 12545
rect 4744 12485 4796 12545
rect 4834 12485 4886 12545
rect 5144 12485 5196 12545
rect 5234 12485 5286 12545
rect 5544 12485 5596 12545
rect 5634 12485 5686 12545
rect 5944 12485 5996 12545
rect 2834 12225 2886 12285
rect 3144 12225 3196 12285
rect 3234 12225 3286 12285
rect 3544 12225 3596 12285
rect 3634 12225 3686 12285
rect 3944 12225 3996 12285
rect 4034 12225 4086 12285
rect 4344 12225 4396 12285
rect 4434 12225 4486 12285
rect 4744 12225 4796 12285
rect 4834 12225 4886 12285
rect 5144 12225 5196 12285
rect 5234 12225 5286 12285
rect 5544 12225 5596 12285
rect 5634 12225 5686 12285
rect 5944 12225 5996 12285
rect 6034 12485 6086 12545
rect 6344 12485 6396 12545
rect 6434 12485 6486 12545
rect 6744 12485 6796 12545
rect 6834 12485 6886 12545
rect 7144 12485 7196 12545
rect 7234 12485 7286 12545
rect 7544 12485 7596 12545
rect 6034 12225 6086 12285
rect 6344 12225 6396 12285
rect 6434 12225 6486 12285
rect 6744 12225 6796 12285
rect 6834 12225 6886 12285
rect 7144 12225 7196 12285
rect 7234 12225 7286 12285
rect 7544 12225 7596 12285
rect 7634 12485 7686 12545
rect 7944 12485 7996 12545
rect 8034 12485 8086 12545
rect 8344 12485 8396 12545
rect 7634 12225 7686 12285
rect 7944 12225 7996 12285
rect 8034 12225 8086 12285
rect 8344 12225 8396 12285
rect 8434 12485 8486 12545
rect 8744 12485 8796 12545
rect 8434 12225 8486 12285
rect 8744 12225 8796 12285
rect 8834 12485 8886 12545
rect 9144 12485 9196 12545
rect 8834 12225 8886 12285
rect 9144 12225 9196 12285
rect 9234 12485 9286 12545
rect 9544 12485 9596 12545
rect 9634 12485 9686 12545
rect 9944 12485 9996 12545
rect 9234 12225 9286 12285
rect 9544 12225 9596 12285
rect 9634 12225 9686 12285
rect 9944 12225 9996 12285
rect 10034 12485 10086 12545
rect 10344 12485 10396 12545
rect 10434 12485 10486 12545
rect 10744 12485 10796 12545
rect 10834 12485 10886 12545
rect 11144 12485 11196 12545
rect 10034 12225 10086 12285
rect 10344 12225 10396 12285
rect 10434 12225 10486 12285
rect 10744 12225 10796 12285
rect 10834 12225 10886 12285
rect 11144 12225 11196 12285
rect 11234 12485 11286 12545
rect 11544 12485 11596 12545
rect 11234 12225 11286 12285
rect 11544 12225 11596 12285
rect 11634 12485 11686 12545
rect 11944 12485 11996 12545
rect 11634 12225 11686 12285
rect 11944 12225 11996 12285
rect 12034 12485 12086 12545
rect 12344 12485 12396 12545
rect 12434 12485 12486 12545
rect 12744 12485 12796 12545
rect 12834 12485 12886 12545
rect 13144 12485 13196 12545
rect 12034 12225 12086 12285
rect 12344 12225 12396 12285
rect 12434 12225 12486 12285
rect 12744 12225 12796 12285
rect 12834 12225 12886 12285
rect 13144 12225 13196 12285
rect -366 12115 -330 12175
rect -330 12115 -314 12175
rect -56 12115 -4 12175
rect -366 11855 -330 11915
rect -330 11855 -314 11915
rect -56 11855 -4 11915
rect 34 12115 86 12175
rect 344 12115 396 12175
rect 434 12115 486 12175
rect 744 12115 796 12175
rect 834 12115 886 12175
rect 1144 12115 1196 12175
rect 1234 12115 1286 12175
rect 1544 12115 1596 12175
rect 1634 12115 1686 12175
rect 1944 12115 1996 12175
rect 2034 12115 2086 12175
rect 2344 12115 2396 12175
rect 2434 12115 2486 12175
rect 2744 12115 2796 12175
rect 34 11855 86 11915
rect 344 11855 396 11915
rect 434 11855 486 11915
rect 744 11855 796 11915
rect 834 11855 886 11915
rect 1144 11855 1196 11915
rect 1234 11855 1286 11915
rect 1544 11855 1596 11915
rect 1634 11855 1686 11915
rect 1944 11855 1996 11915
rect 2034 11855 2086 11915
rect 2344 11855 2396 11915
rect 2434 11855 2486 11915
rect 2744 11855 2796 11915
rect 2834 12115 2886 12175
rect 3144 12115 3196 12175
rect 3234 12115 3286 12175
rect 3544 12115 3596 12175
rect 3634 12115 3686 12175
rect 3944 12115 3996 12175
rect 4034 12115 4086 12175
rect 4344 12115 4396 12175
rect 4434 12115 4486 12175
rect 4744 12115 4796 12175
rect 4834 12115 4886 12175
rect 5144 12115 5196 12175
rect 5234 12115 5286 12175
rect 5544 12115 5596 12175
rect 2834 11855 2886 11915
rect 3144 11855 3196 11915
rect 3234 11855 3286 11915
rect 3544 11855 3596 11915
rect 3634 11855 3686 11915
rect 3944 11855 3996 11915
rect 4034 11855 4086 11915
rect 4344 11855 4396 11915
rect 4434 11855 4486 11915
rect 4744 11855 4796 11915
rect 4834 11855 4886 11915
rect 5144 11855 5196 11915
rect 5234 11855 5286 11915
rect 5544 11855 5596 11915
rect 5634 12115 5686 12175
rect 5944 12115 5996 12175
rect 6034 12115 6086 12175
rect 6344 12115 6396 12175
rect 6434 12115 6486 12175
rect 6744 12115 6796 12175
rect 6834 12115 6886 12175
rect 7144 12115 7196 12175
rect 7234 12115 7286 12175
rect 7544 12115 7596 12175
rect 5634 11855 5686 11915
rect 5944 11855 5996 11915
rect 6034 11855 6086 11915
rect 6344 11855 6396 11915
rect 6434 11855 6486 11915
rect 6744 11855 6796 11915
rect 6834 11855 6886 11915
rect 7144 11855 7196 11915
rect 7234 11855 7286 11915
rect 7544 11855 7596 11915
rect 7634 12115 7686 12175
rect 7944 12115 7996 12175
rect 8034 12115 8086 12175
rect 8344 12115 8396 12175
rect 7634 11855 7686 11915
rect 7944 11855 7996 11915
rect 8034 11855 8086 11915
rect 8344 11855 8396 11915
rect 8434 12115 8486 12175
rect 8744 12115 8796 12175
rect 8434 11855 8486 11915
rect 8744 11855 8796 11915
rect 8834 12115 8886 12175
rect 9144 12115 9196 12175
rect 9234 12115 9286 12175
rect 9544 12115 9596 12175
rect 9634 12115 9686 12175
rect 9944 12115 9996 12175
rect 8834 11855 8886 11915
rect 9144 11855 9196 11915
rect 9234 11855 9286 11915
rect 9544 11855 9596 11915
rect 9634 11855 9686 11915
rect 9944 11855 9996 11915
rect 10034 12115 10086 12175
rect 10344 12115 10396 12175
rect 10434 12115 10486 12175
rect 10744 12115 10796 12175
rect 10834 12115 10886 12175
rect 11144 12115 11196 12175
rect 10034 11855 10086 11915
rect 10344 11855 10396 11915
rect 10434 11855 10486 11915
rect 10744 11855 10796 11915
rect 10834 11855 10886 11915
rect 11144 11855 11196 11915
rect 11234 12115 11286 12175
rect 11544 12115 11596 12175
rect 11234 11855 11286 11915
rect 11544 11855 11596 11915
rect 11634 12115 11686 12175
rect 11944 12115 11996 12175
rect 11634 11855 11686 11915
rect 11944 11855 11996 11915
rect 12034 12115 12086 12175
rect 12344 12115 12396 12175
rect 12034 11855 12086 11915
rect 12344 11855 12396 11915
rect 12434 12115 12486 12175
rect 12744 12115 12796 12175
rect 12834 12115 12886 12175
rect 13144 12115 13196 12175
rect 12434 11855 12486 11915
rect 12744 11855 12796 11915
rect 12834 11855 12886 11915
rect 13144 11855 13196 11915
rect -366 11745 -330 11805
rect -330 11745 -314 11805
rect -56 11745 -4 11805
rect -366 11485 -330 11545
rect -330 11485 -314 11545
rect -56 11485 -4 11545
rect 34 11745 86 11805
rect 344 11745 396 11805
rect 434 11745 486 11805
rect 744 11745 796 11805
rect 834 11745 886 11805
rect 1144 11745 1196 11805
rect 1234 11745 1286 11805
rect 1544 11745 1596 11805
rect 1634 11745 1686 11805
rect 1944 11745 1996 11805
rect 2034 11745 2086 11805
rect 2344 11745 2396 11805
rect 2434 11745 2486 11805
rect 2744 11745 2796 11805
rect 34 11485 86 11545
rect 344 11485 396 11545
rect 434 11485 486 11545
rect 744 11485 796 11545
rect 834 11485 886 11545
rect 1144 11485 1196 11545
rect 1234 11485 1286 11545
rect 1544 11485 1596 11545
rect 1634 11485 1686 11545
rect 1944 11485 1996 11545
rect 2034 11485 2086 11545
rect 2344 11485 2396 11545
rect 2434 11485 2486 11545
rect 2744 11485 2796 11545
rect 2834 11745 2886 11805
rect 3144 11745 3196 11805
rect 3234 11745 3286 11805
rect 3544 11745 3596 11805
rect 3634 11745 3686 11805
rect 3944 11745 3996 11805
rect 4034 11745 4086 11805
rect 4344 11745 4396 11805
rect 4434 11745 4486 11805
rect 4744 11745 4796 11805
rect 4834 11745 4886 11805
rect 5144 11745 5196 11805
rect 5234 11745 5286 11805
rect 5544 11745 5596 11805
rect 2834 11485 2886 11545
rect 3144 11485 3196 11545
rect 3234 11485 3286 11545
rect 3544 11485 3596 11545
rect 3634 11485 3686 11545
rect 3944 11485 3996 11545
rect 4034 11485 4086 11545
rect 4344 11485 4396 11545
rect 4434 11485 4486 11545
rect 4744 11485 4796 11545
rect 4834 11485 4886 11545
rect 5144 11485 5196 11545
rect 5234 11485 5286 11545
rect 5544 11485 5596 11545
rect 5634 11745 5686 11805
rect 5944 11745 5996 11805
rect 6034 11745 6086 11805
rect 6344 11745 6396 11805
rect 6434 11745 6486 11805
rect 6744 11745 6796 11805
rect 6834 11745 6886 11805
rect 7144 11745 7196 11805
rect 7234 11745 7286 11805
rect 7544 11745 7596 11805
rect 5634 11485 5686 11545
rect 5944 11485 5996 11545
rect 6034 11485 6086 11545
rect 6344 11485 6396 11545
rect 6434 11485 6486 11545
rect 6744 11485 6796 11545
rect 6834 11485 6886 11545
rect 7144 11485 7196 11545
rect 7234 11485 7286 11545
rect 7544 11485 7596 11545
rect 7634 11745 7686 11805
rect 7944 11745 7996 11805
rect 8034 11745 8086 11805
rect 8344 11745 8396 11805
rect 7634 11485 7686 11545
rect 7944 11485 7996 11545
rect 8034 11485 8086 11545
rect 8344 11485 8396 11545
rect 8434 11745 8486 11805
rect 8744 11745 8796 11805
rect 8434 11485 8486 11545
rect 8744 11485 8796 11545
rect 8834 11745 8886 11805
rect 9144 11745 9196 11805
rect 9234 11745 9286 11805
rect 9544 11745 9596 11805
rect 9634 11745 9686 11805
rect 9944 11745 9996 11805
rect 8834 11485 8886 11545
rect 9144 11485 9196 11545
rect 9234 11485 9286 11545
rect 9544 11485 9596 11545
rect 9634 11485 9686 11545
rect 9944 11485 9996 11545
rect 10034 11745 10086 11805
rect 10344 11745 10396 11805
rect 10434 11745 10486 11805
rect 10744 11745 10796 11805
rect 10834 11745 10886 11805
rect 11144 11745 11196 11805
rect 10034 11485 10086 11545
rect 10344 11485 10396 11545
rect 10434 11485 10486 11545
rect 10744 11485 10796 11545
rect 10834 11485 10886 11545
rect 11144 11485 11196 11545
rect 11234 11745 11286 11805
rect 11544 11745 11596 11805
rect 11234 11485 11286 11545
rect 11544 11485 11596 11545
rect 11634 11745 11686 11805
rect 11944 11745 11996 11805
rect 11634 11485 11686 11545
rect 11944 11485 11996 11545
rect 12034 11745 12086 11805
rect 12344 11745 12396 11805
rect 12034 11485 12086 11545
rect 12344 11485 12396 11545
rect 12434 11745 12486 11805
rect 12744 11745 12796 11805
rect 12834 11745 12886 11805
rect 13144 11745 13196 11805
rect 12434 11485 12486 11545
rect 12744 11485 12796 11545
rect 12834 11485 12886 11545
rect 13144 11485 13196 11545
rect -366 11375 -330 11435
rect -330 11375 -314 11435
rect -56 11375 -4 11435
rect -366 11115 -330 11175
rect -330 11115 -314 11175
rect -56 11115 -4 11175
rect 34 11375 86 11435
rect 344 11375 396 11435
rect 434 11375 486 11435
rect 744 11375 796 11435
rect 834 11375 886 11435
rect 1144 11375 1196 11435
rect 1234 11375 1286 11435
rect 1544 11375 1596 11435
rect 1634 11375 1686 11435
rect 1944 11375 1996 11435
rect 2034 11375 2086 11435
rect 2344 11375 2396 11435
rect 2434 11375 2486 11435
rect 2744 11375 2796 11435
rect 34 11115 86 11175
rect 344 11115 396 11175
rect 434 11115 486 11175
rect 744 11115 796 11175
rect 834 11115 886 11175
rect 1144 11115 1196 11175
rect 1234 11115 1286 11175
rect 1544 11115 1596 11175
rect 1634 11115 1686 11175
rect 1944 11115 1996 11175
rect 2034 11115 2086 11175
rect 2344 11115 2396 11175
rect 2434 11115 2486 11175
rect 2744 11115 2796 11175
rect 2834 11375 2886 11435
rect 3144 11375 3196 11435
rect 3234 11375 3286 11435
rect 3544 11375 3596 11435
rect 3634 11375 3686 11435
rect 3944 11375 3996 11435
rect 4034 11375 4086 11435
rect 4344 11375 4396 11435
rect 4434 11375 4486 11435
rect 4744 11375 4796 11435
rect 4834 11375 4886 11435
rect 5144 11375 5196 11435
rect 5234 11375 5286 11435
rect 5544 11375 5596 11435
rect 5634 11375 5686 11435
rect 5944 11375 5996 11435
rect 2834 11115 2886 11175
rect 3144 11115 3196 11175
rect 3234 11115 3286 11175
rect 3544 11115 3596 11175
rect 3634 11115 3686 11175
rect 3944 11115 3996 11175
rect 4034 11115 4086 11175
rect 4344 11115 4396 11175
rect 4434 11115 4486 11175
rect 4744 11115 4796 11175
rect 4834 11115 4886 11175
rect 5144 11115 5196 11175
rect 5234 11115 5286 11175
rect 5544 11115 5596 11175
rect 5634 11115 5686 11175
rect 5944 11115 5996 11175
rect 6034 11375 6086 11435
rect 6344 11375 6396 11435
rect 6434 11375 6486 11435
rect 6744 11375 6796 11435
rect 6834 11375 6886 11435
rect 7144 11375 7196 11435
rect 7234 11375 7286 11435
rect 7544 11375 7596 11435
rect 6034 11115 6086 11175
rect 6344 11115 6396 11175
rect 6434 11115 6486 11175
rect 6744 11115 6796 11175
rect 6834 11115 6886 11175
rect 7144 11115 7196 11175
rect 7234 11115 7286 11175
rect 7544 11115 7596 11175
rect 7634 11375 7686 11435
rect 7944 11375 7996 11435
rect 8034 11375 8086 11435
rect 8344 11375 8396 11435
rect 7634 11115 7686 11175
rect 7944 11115 7996 11175
rect 8034 11115 8086 11175
rect 8344 11115 8396 11175
rect 8434 11375 8486 11435
rect 8744 11375 8796 11435
rect 8434 11115 8486 11175
rect 8744 11115 8796 11175
rect 8834 11375 8886 11435
rect 9144 11375 9196 11435
rect 8834 11115 8886 11175
rect 9144 11115 9196 11175
rect 9234 11375 9286 11435
rect 9544 11375 9596 11435
rect 9634 11375 9686 11435
rect 9944 11375 9996 11435
rect 9234 11115 9286 11175
rect 9544 11115 9596 11175
rect 9634 11115 9686 11175
rect 9944 11115 9996 11175
rect 10034 11375 10086 11435
rect 10344 11375 10396 11435
rect 10434 11375 10486 11435
rect 10744 11375 10796 11435
rect 10834 11375 10886 11435
rect 11144 11375 11196 11435
rect 10034 11115 10086 11175
rect 10344 11115 10396 11175
rect 10434 11115 10486 11175
rect 10744 11115 10796 11175
rect 10834 11115 10886 11175
rect 11144 11115 11196 11175
rect 11234 11375 11286 11435
rect 11544 11375 11596 11435
rect 11234 11115 11286 11175
rect 11544 11115 11596 11175
rect 11634 11375 11686 11435
rect 11944 11375 11996 11435
rect 11634 11115 11686 11175
rect 11944 11115 11996 11175
rect 12034 11375 12086 11435
rect 12344 11375 12396 11435
rect 12434 11375 12486 11435
rect 12744 11375 12796 11435
rect 12834 11375 12886 11435
rect 13144 11375 13196 11435
rect 12034 11115 12086 11175
rect 12344 11115 12396 11175
rect 12434 11115 12486 11175
rect 12744 11115 12796 11175
rect 12834 11115 12886 11175
rect 13144 11115 13196 11175
rect -366 11005 -330 11065
rect -330 11005 -314 11065
rect -56 11005 -4 11065
rect -366 10745 -330 10805
rect -330 10745 -314 10805
rect -56 10745 -4 10805
rect 34 11005 86 11065
rect 344 11005 396 11065
rect 434 11005 486 11065
rect 744 11005 796 11065
rect 834 11005 886 11065
rect 1144 11005 1196 11065
rect 1234 11005 1286 11065
rect 1544 11005 1596 11065
rect 1634 11005 1686 11065
rect 1944 11005 1996 11065
rect 2034 11005 2086 11065
rect 2344 11005 2396 11065
rect 2434 11005 2486 11065
rect 2744 11005 2796 11065
rect 34 10745 86 10805
rect 344 10745 396 10805
rect 434 10745 486 10805
rect 744 10745 796 10805
rect 834 10745 886 10805
rect 1144 10745 1196 10805
rect 1234 10745 1286 10805
rect 1544 10745 1596 10805
rect 1634 10745 1686 10805
rect 1944 10745 1996 10805
rect 2034 10745 2086 10805
rect 2344 10745 2396 10805
rect 2434 10745 2486 10805
rect 2744 10745 2796 10805
rect 2834 11005 2886 11065
rect 3144 11005 3196 11065
rect 3234 11005 3286 11065
rect 3544 11005 3596 11065
rect 3634 11005 3686 11065
rect 3944 11005 3996 11065
rect 4034 11005 4086 11065
rect 4344 11005 4396 11065
rect 4434 11005 4486 11065
rect 4744 11005 4796 11065
rect 4834 11005 4886 11065
rect 5144 11005 5196 11065
rect 5234 11005 5286 11065
rect 5544 11005 5596 11065
rect 5634 11005 5686 11065
rect 5944 11005 5996 11065
rect 2834 10745 2886 10805
rect 3144 10745 3196 10805
rect 3234 10745 3286 10805
rect 3544 10745 3596 10805
rect 3634 10745 3686 10805
rect 3944 10745 3996 10805
rect 4034 10745 4086 10805
rect 4344 10745 4396 10805
rect 4434 10745 4486 10805
rect 4744 10745 4796 10805
rect 4834 10745 4886 10805
rect 5144 10745 5196 10805
rect 5234 10745 5286 10805
rect 5544 10745 5596 10805
rect 5634 10745 5686 10805
rect 5944 10745 5996 10805
rect 6034 11005 6086 11065
rect 6344 11005 6396 11065
rect 6434 11005 6486 11065
rect 6744 11005 6796 11065
rect 6834 11005 6886 11065
rect 7144 11005 7196 11065
rect 7234 11005 7286 11065
rect 7544 11005 7596 11065
rect 6034 10745 6086 10805
rect 6344 10745 6396 10805
rect 6434 10745 6486 10805
rect 6744 10745 6796 10805
rect 6834 10745 6886 10805
rect 7144 10745 7196 10805
rect 7234 10745 7286 10805
rect 7544 10745 7596 10805
rect 7634 11005 7686 11065
rect 7944 11005 7996 11065
rect 8034 11005 8086 11065
rect 8344 11005 8396 11065
rect 7634 10745 7686 10805
rect 7944 10745 7996 10805
rect 8034 10745 8086 10805
rect 8344 10745 8396 10805
rect 8434 11005 8486 11065
rect 8744 11005 8796 11065
rect 8434 10745 8486 10805
rect 8744 10745 8796 10805
rect 8834 11005 8886 11065
rect 9144 11005 9196 11065
rect 8834 10745 8886 10805
rect 9144 10745 9196 10805
rect 9234 11005 9286 11065
rect 9544 11005 9596 11065
rect 9634 11005 9686 11065
rect 9944 11005 9996 11065
rect 10034 11005 10086 11065
rect 10344 11005 10396 11065
rect 9234 10745 9286 10805
rect 9544 10745 9596 10805
rect 9634 10745 9686 10805
rect 9944 10745 9996 10805
rect 10034 10745 10086 10805
rect 10344 10745 10396 10805
rect 10434 11005 10486 11065
rect 10744 11005 10796 11065
rect 10834 11005 10886 11065
rect 11144 11005 11196 11065
rect 10434 10745 10486 10805
rect 10744 10745 10796 10805
rect 10834 10745 10886 10805
rect 11144 10745 11196 10805
rect 11234 11005 11286 11065
rect 11544 11005 11596 11065
rect 11234 10745 11286 10805
rect 11544 10745 11596 10805
rect 11634 11005 11686 11065
rect 11944 11005 11996 11065
rect 11634 10745 11686 10805
rect 11944 10745 11996 10805
rect 12034 11005 12086 11065
rect 12344 11005 12396 11065
rect 12434 11005 12486 11065
rect 12744 11005 12796 11065
rect 12834 11005 12886 11065
rect 13144 11005 13196 11065
rect 12034 10745 12086 10805
rect 12344 10745 12396 10805
rect 12434 10745 12486 10805
rect 12744 10745 12796 10805
rect 12834 10745 12886 10805
rect 13144 10745 13196 10805
rect -366 10635 -330 10695
rect -330 10635 -314 10695
rect -56 10635 -4 10695
rect -366 10375 -330 10435
rect -330 10375 -314 10435
rect -56 10375 -4 10435
rect 34 10635 86 10695
rect 344 10635 396 10695
rect 434 10635 486 10695
rect 744 10635 796 10695
rect 834 10635 886 10695
rect 1144 10635 1196 10695
rect 1234 10635 1286 10695
rect 1544 10635 1596 10695
rect 1634 10635 1686 10695
rect 1944 10635 1996 10695
rect 2034 10635 2086 10695
rect 2344 10635 2396 10695
rect 2434 10635 2486 10695
rect 2744 10635 2796 10695
rect 34 10375 86 10435
rect 344 10375 396 10435
rect 434 10375 486 10435
rect 744 10375 796 10435
rect 834 10375 886 10435
rect 1144 10375 1196 10435
rect 1234 10375 1286 10435
rect 1544 10375 1596 10435
rect 1634 10375 1686 10435
rect 1944 10375 1996 10435
rect 2034 10375 2086 10435
rect 2344 10375 2396 10435
rect 2434 10375 2486 10435
rect 2744 10375 2796 10435
rect 2834 10635 2886 10695
rect 3144 10635 3196 10695
rect 3234 10635 3286 10695
rect 3544 10635 3596 10695
rect 3634 10635 3686 10695
rect 3944 10635 3996 10695
rect 4034 10635 4086 10695
rect 4344 10635 4396 10695
rect 4434 10635 4486 10695
rect 4744 10635 4796 10695
rect 4834 10635 4886 10695
rect 5144 10635 5196 10695
rect 5234 10635 5286 10695
rect 5544 10635 5596 10695
rect 5634 10635 5686 10695
rect 5944 10635 5996 10695
rect 2834 10375 2886 10435
rect 3144 10375 3196 10435
rect 3234 10375 3286 10435
rect 3544 10375 3596 10435
rect 3634 10375 3686 10435
rect 3944 10375 3996 10435
rect 4034 10375 4086 10435
rect 4344 10375 4396 10435
rect 4434 10375 4486 10435
rect 4744 10375 4796 10435
rect 4834 10375 4886 10435
rect 5144 10375 5196 10435
rect 5234 10375 5286 10435
rect 5544 10375 5596 10435
rect 5634 10375 5686 10435
rect 5944 10375 5996 10435
rect 6034 10635 6086 10695
rect 6344 10635 6396 10695
rect 6434 10635 6486 10695
rect 6744 10635 6796 10695
rect 6834 10635 6886 10695
rect 7144 10635 7196 10695
rect 7234 10635 7286 10695
rect 7544 10635 7596 10695
rect 6034 10375 6086 10435
rect 6344 10375 6396 10435
rect 6434 10375 6486 10435
rect 6744 10375 6796 10435
rect 6834 10375 6886 10435
rect 7144 10375 7196 10435
rect 7234 10375 7286 10435
rect 7544 10375 7596 10435
rect 7634 10635 7686 10695
rect 7944 10635 7996 10695
rect 8034 10635 8086 10695
rect 8344 10635 8396 10695
rect 7634 10375 7686 10435
rect 7944 10375 7996 10435
rect 8034 10375 8086 10435
rect 8344 10375 8396 10435
rect 8434 10635 8486 10695
rect 8744 10635 8796 10695
rect 8434 10375 8486 10435
rect 8744 10375 8796 10435
rect 8834 10635 8886 10695
rect 9144 10635 9196 10695
rect 8834 10375 8886 10435
rect 9144 10375 9196 10435
rect 9234 10635 9286 10695
rect 9544 10635 9596 10695
rect 9634 10635 9686 10695
rect 9944 10635 9996 10695
rect 10034 10635 10086 10695
rect 10344 10635 10396 10695
rect 9234 10375 9286 10435
rect 9544 10375 9596 10435
rect 9634 10375 9686 10435
rect 9944 10375 9996 10435
rect 10034 10375 10086 10435
rect 10344 10375 10396 10435
rect 10434 10635 10486 10695
rect 10744 10635 10796 10695
rect 10834 10635 10886 10695
rect 11144 10635 11196 10695
rect 10434 10375 10486 10435
rect 10744 10375 10796 10435
rect 10834 10375 10886 10435
rect 11144 10375 11196 10435
rect 11234 10635 11286 10695
rect 11544 10635 11596 10695
rect 11634 10635 11686 10695
rect 11944 10635 11996 10695
rect 12034 10635 12086 10695
rect 12344 10635 12396 10695
rect 12434 10635 12486 10695
rect 12744 10635 12796 10695
rect 12834 10635 12886 10695
rect 13144 10635 13196 10695
rect 11234 10375 11286 10435
rect 11544 10375 11596 10435
rect 11634 10375 11686 10435
rect 11944 10375 11996 10435
rect 12034 10375 12086 10435
rect 12344 10375 12396 10435
rect 12434 10375 12486 10435
rect 12744 10375 12796 10435
rect 12834 10375 12886 10435
rect 13144 10375 13196 10435
rect -366 10265 -330 10325
rect -330 10265 -314 10325
rect -56 10265 -4 10325
rect -366 10005 -330 10065
rect -330 10005 -314 10065
rect -56 10005 -4 10065
rect 34 10265 86 10325
rect 344 10265 396 10325
rect 434 10265 486 10325
rect 744 10265 796 10325
rect 834 10265 886 10325
rect 1144 10265 1196 10325
rect 1234 10265 1286 10325
rect 1544 10265 1596 10325
rect 1634 10265 1686 10325
rect 1944 10265 1996 10325
rect 2034 10265 2086 10325
rect 2344 10265 2396 10325
rect 2434 10265 2486 10325
rect 2744 10265 2796 10325
rect 34 10005 86 10065
rect 344 10005 396 10065
rect 434 10005 486 10065
rect 744 10005 796 10065
rect 834 10005 886 10065
rect 1144 10005 1196 10065
rect 1234 10005 1286 10065
rect 1544 10005 1596 10065
rect 1634 10005 1686 10065
rect 1944 10005 1996 10065
rect 2034 10005 2086 10065
rect 2344 10005 2396 10065
rect 2434 10005 2486 10065
rect 2744 10005 2796 10065
rect 2834 10265 2886 10325
rect 3144 10265 3196 10325
rect 3234 10265 3286 10325
rect 3544 10265 3596 10325
rect 3634 10265 3686 10325
rect 3944 10265 3996 10325
rect 4034 10265 4086 10325
rect 4344 10265 4396 10325
rect 4434 10265 4486 10325
rect 4744 10265 4796 10325
rect 4834 10265 4886 10325
rect 5144 10265 5196 10325
rect 5234 10265 5286 10325
rect 5544 10265 5596 10325
rect 5634 10265 5686 10325
rect 5944 10265 5996 10325
rect 2834 10005 2886 10065
rect 3144 10005 3196 10065
rect 3234 10005 3286 10065
rect 3544 10005 3596 10065
rect 3634 10005 3686 10065
rect 3944 10005 3996 10065
rect 4034 10005 4086 10065
rect 4344 10005 4396 10065
rect 4434 10005 4486 10065
rect 4744 10005 4796 10065
rect 4834 10005 4886 10065
rect 5144 10005 5196 10065
rect 5234 10005 5286 10065
rect 5544 10005 5596 10065
rect 5634 10005 5686 10065
rect 5944 10005 5996 10065
rect 6034 10265 6086 10325
rect 6344 10265 6396 10325
rect 6434 10265 6486 10325
rect 6744 10265 6796 10325
rect 6834 10265 6886 10325
rect 7144 10265 7196 10325
rect 7234 10265 7286 10325
rect 7544 10265 7596 10325
rect 6034 10005 6086 10065
rect 6344 10005 6396 10065
rect 6434 10005 6486 10065
rect 6744 10005 6796 10065
rect 6834 10005 6886 10065
rect 7144 10005 7196 10065
rect 7234 10005 7286 10065
rect 7544 10005 7596 10065
rect 7634 10265 7686 10325
rect 7944 10265 7996 10325
rect 8034 10265 8086 10325
rect 8344 10265 8396 10325
rect 7634 10005 7686 10065
rect 7944 10005 7996 10065
rect 8034 10005 8086 10065
rect 8344 10005 8396 10065
rect 8434 10265 8486 10325
rect 8744 10265 8796 10325
rect 8434 10005 8486 10065
rect 8744 10005 8796 10065
rect 8834 10265 8886 10325
rect 9144 10265 9196 10325
rect 8834 10005 8886 10065
rect 9144 10005 9196 10065
rect 9234 10265 9286 10325
rect 9544 10265 9596 10325
rect 9634 10265 9686 10325
rect 9944 10265 9996 10325
rect 10034 10265 10086 10325
rect 10344 10265 10396 10325
rect 9234 10005 9286 10065
rect 9544 10005 9596 10065
rect 9634 10005 9686 10065
rect 9944 10005 9996 10065
rect 10034 10005 10086 10065
rect 10344 10005 10396 10065
rect 10434 10265 10486 10325
rect 10744 10265 10796 10325
rect 10834 10265 10886 10325
rect 11144 10265 11196 10325
rect 11234 10265 11286 10325
rect 11544 10265 11596 10325
rect 11634 10265 11686 10325
rect 11944 10265 11996 10325
rect 12034 10265 12086 10325
rect 12344 10265 12396 10325
rect 12434 10265 12486 10325
rect 12744 10265 12796 10325
rect 12834 10265 12886 10325
rect 13144 10265 13196 10325
rect 10434 10005 10486 10065
rect 10744 10005 10796 10065
rect 10834 10005 10886 10065
rect 11144 10005 11196 10065
rect 11234 10005 11286 10065
rect 11544 10005 11596 10065
rect 11634 10005 11686 10065
rect 11944 10005 11996 10065
rect 12034 10005 12086 10065
rect 12344 10005 12396 10065
rect 12434 10005 12486 10065
rect 12744 10005 12796 10065
rect 12834 10005 12886 10065
rect 13144 10005 13196 10065
rect -366 9895 -330 9955
rect -330 9895 -314 9955
rect -56 9895 -4 9955
rect -366 9635 -330 9695
rect -330 9635 -314 9695
rect -56 9635 -4 9695
rect 34 9895 86 9955
rect 344 9895 396 9955
rect 434 9895 486 9955
rect 744 9895 796 9955
rect 834 9895 886 9955
rect 1144 9895 1196 9955
rect 1234 9895 1286 9955
rect 1544 9895 1596 9955
rect 1634 9895 1686 9955
rect 1944 9895 1996 9955
rect 2034 9895 2086 9955
rect 2344 9895 2396 9955
rect 2434 9895 2486 9955
rect 2744 9895 2796 9955
rect 34 9635 86 9695
rect 344 9635 396 9695
rect 434 9635 486 9695
rect 744 9635 796 9695
rect 834 9635 886 9695
rect 1144 9635 1196 9695
rect 1234 9635 1286 9695
rect 1544 9635 1596 9695
rect 1634 9635 1686 9695
rect 1944 9635 1996 9695
rect 2034 9635 2086 9695
rect 2344 9635 2396 9695
rect 2434 9635 2486 9695
rect 2744 9635 2796 9695
rect 2834 9895 2886 9955
rect 3144 9895 3196 9955
rect 3234 9895 3286 9955
rect 3544 9895 3596 9955
rect 3634 9895 3686 9955
rect 3944 9895 3996 9955
rect 4034 9895 4086 9955
rect 4344 9895 4396 9955
rect 4434 9895 4486 9955
rect 4744 9895 4796 9955
rect 4834 9895 4886 9955
rect 5144 9895 5196 9955
rect 5234 9895 5286 9955
rect 5544 9895 5596 9955
rect 5634 9895 5686 9955
rect 5944 9895 5996 9955
rect 2834 9635 2886 9695
rect 3144 9635 3196 9695
rect 3234 9635 3286 9695
rect 3544 9635 3596 9695
rect 3634 9635 3686 9695
rect 3944 9635 3996 9695
rect 4034 9635 4086 9695
rect 4344 9635 4396 9695
rect 4434 9635 4486 9695
rect 4744 9635 4796 9695
rect 4834 9635 4886 9695
rect 5144 9635 5196 9695
rect 5234 9635 5286 9695
rect 5544 9635 5596 9695
rect 5634 9635 5686 9695
rect 5944 9635 5996 9695
rect 6034 9895 6086 9955
rect 6344 9895 6396 9955
rect 6434 9895 6486 9955
rect 6744 9895 6796 9955
rect 6834 9895 6886 9955
rect 7144 9895 7196 9955
rect 7234 9895 7286 9955
rect 7544 9895 7596 9955
rect 6034 9635 6086 9695
rect 6344 9635 6396 9695
rect 6434 9635 6486 9695
rect 6744 9635 6796 9695
rect 6834 9635 6886 9695
rect 7144 9635 7196 9695
rect 7234 9635 7286 9695
rect 7544 9635 7596 9695
rect 7634 9895 7686 9955
rect 7944 9895 7996 9955
rect 8034 9895 8086 9955
rect 8344 9895 8396 9955
rect 7634 9635 7686 9695
rect 7944 9635 7996 9695
rect 8034 9635 8086 9695
rect 8344 9635 8396 9695
rect 8434 9895 8486 9955
rect 8744 9895 8796 9955
rect 8434 9635 8486 9695
rect 8744 9635 8796 9695
rect 8834 9895 8886 9955
rect 9144 9895 9196 9955
rect 8834 9635 8886 9695
rect 9144 9635 9196 9695
rect 9234 9895 9286 9955
rect 9544 9895 9596 9955
rect 9634 9895 9686 9955
rect 9944 9895 9996 9955
rect 10034 9895 10086 9955
rect 10344 9895 10396 9955
rect 10434 9895 10486 9955
rect 10744 9895 10796 9955
rect 10834 9895 10886 9955
rect 11144 9895 11196 9955
rect 11234 9895 11286 9955
rect 11544 9895 11596 9955
rect 11634 9895 11686 9955
rect 11944 9895 11996 9955
rect 12034 9895 12086 9955
rect 12344 9895 12396 9955
rect 12434 9895 12486 9955
rect 12744 9895 12796 9955
rect 12834 9895 12886 9955
rect 13144 9895 13196 9955
rect 9234 9635 9286 9695
rect 9544 9635 9596 9695
rect 9634 9635 9686 9695
rect 9944 9635 9996 9695
rect 10034 9635 10086 9695
rect 10344 9635 10396 9695
rect 10434 9635 10486 9695
rect 10744 9635 10796 9695
rect 10834 9635 10886 9695
rect 11144 9635 11196 9695
rect 11234 9635 11286 9695
rect 11544 9635 11596 9695
rect 11634 9635 11686 9695
rect 11944 9635 11996 9695
rect 12034 9635 12086 9695
rect 12344 9635 12396 9695
rect 12434 9635 12486 9695
rect 12744 9635 12796 9695
rect 12834 9635 12886 9695
rect 13144 9635 13196 9695
rect -366 9525 -330 9585
rect -330 9525 -314 9585
rect -56 9525 -4 9585
rect -366 9265 -330 9325
rect -330 9265 -314 9325
rect -56 9265 -4 9325
rect 34 9525 86 9585
rect 344 9525 396 9585
rect 434 9525 486 9585
rect 744 9525 796 9585
rect 834 9525 886 9585
rect 1144 9525 1196 9585
rect 1234 9525 1286 9585
rect 1544 9525 1596 9585
rect 1634 9525 1686 9585
rect 1944 9525 1996 9585
rect 2034 9525 2086 9585
rect 2344 9525 2396 9585
rect 2434 9525 2486 9585
rect 2744 9525 2796 9585
rect 34 9265 86 9325
rect 344 9265 396 9325
rect 434 9265 486 9325
rect 744 9265 796 9325
rect 834 9265 886 9325
rect 1144 9265 1196 9325
rect 1234 9265 1286 9325
rect 1544 9265 1596 9325
rect 1634 9265 1686 9325
rect 1944 9265 1996 9325
rect 2034 9265 2086 9325
rect 2344 9265 2396 9325
rect 2434 9265 2486 9325
rect 2744 9265 2796 9325
rect 2834 9525 2886 9585
rect 3144 9525 3196 9585
rect 3234 9525 3286 9585
rect 3544 9525 3596 9585
rect 3634 9525 3686 9585
rect 3944 9525 3996 9585
rect 4034 9525 4086 9585
rect 4344 9525 4396 9585
rect 4434 9525 4486 9585
rect 4744 9525 4796 9585
rect 4834 9525 4886 9585
rect 5144 9525 5196 9585
rect 5234 9525 5286 9585
rect 5544 9525 5596 9585
rect 5634 9525 5686 9585
rect 5944 9525 5996 9585
rect 2834 9265 2886 9325
rect 3144 9265 3196 9325
rect 3234 9265 3286 9325
rect 3544 9265 3596 9325
rect 3634 9265 3686 9325
rect 3944 9265 3996 9325
rect 4034 9265 4086 9325
rect 4344 9265 4396 9325
rect 4434 9265 4486 9325
rect 4744 9265 4796 9325
rect 4834 9265 4886 9325
rect 5144 9265 5196 9325
rect 5234 9265 5286 9325
rect 5544 9265 5596 9325
rect 5634 9265 5686 9325
rect 5944 9265 5996 9325
rect 6034 9525 6086 9585
rect 6344 9525 6396 9585
rect 6434 9525 6486 9585
rect 6744 9525 6796 9585
rect 6834 9525 6886 9585
rect 7144 9525 7196 9585
rect 7234 9525 7286 9585
rect 7544 9525 7596 9585
rect 6034 9265 6086 9325
rect 6344 9265 6396 9325
rect 6434 9265 6486 9325
rect 6744 9265 6796 9325
rect 6834 9265 6886 9325
rect 7144 9265 7196 9325
rect 7234 9265 7286 9325
rect 7544 9265 7596 9325
rect 7634 9525 7686 9585
rect 7944 9525 7996 9585
rect 8034 9525 8086 9585
rect 8344 9525 8396 9585
rect 7634 9265 7686 9325
rect 7944 9265 7996 9325
rect 8034 9265 8086 9325
rect 8344 9265 8396 9325
rect 8434 9525 8486 9585
rect 8744 9525 8796 9585
rect 8434 9265 8486 9325
rect 8744 9265 8796 9325
rect 8834 9525 8886 9585
rect 9144 9525 9196 9585
rect 8834 9265 8886 9325
rect 9144 9265 9196 9325
rect 9234 9525 9286 9585
rect 9544 9525 9596 9585
rect 9634 9525 9686 9585
rect 9944 9525 9996 9585
rect 10034 9525 10086 9585
rect 10344 9525 10396 9585
rect 10434 9525 10486 9585
rect 10744 9525 10796 9585
rect 10834 9525 10886 9585
rect 11144 9525 11196 9585
rect 11234 9525 11286 9585
rect 11544 9525 11596 9585
rect 11634 9525 11686 9585
rect 11944 9525 11996 9585
rect 12034 9525 12086 9585
rect 12344 9525 12396 9585
rect 12434 9525 12486 9585
rect 12744 9525 12796 9585
rect 12834 9525 12886 9585
rect 13144 9525 13196 9585
rect 9234 9265 9286 9325
rect 9544 9265 9596 9325
rect 9634 9265 9686 9325
rect 9944 9265 9996 9325
rect 10034 9265 10086 9325
rect 10344 9265 10396 9325
rect 10434 9265 10486 9325
rect 10744 9265 10796 9325
rect 10834 9265 10886 9325
rect 11144 9265 11196 9325
rect 11234 9265 11286 9325
rect 11544 9265 11596 9325
rect 11634 9265 11686 9325
rect 11944 9265 11996 9325
rect 12034 9265 12086 9325
rect 12344 9265 12396 9325
rect 12434 9265 12486 9325
rect 12744 9265 12796 9325
rect 12834 9265 12886 9325
rect 13144 9265 13196 9325
rect -366 9155 -330 9215
rect -330 9155 -314 9215
rect -56 9155 -4 9215
rect -366 8895 -330 8955
rect -330 8895 -314 8955
rect -56 8895 -4 8955
rect 34 9155 86 9215
rect 344 9155 396 9215
rect 434 9155 486 9215
rect 744 9155 796 9215
rect 834 9155 886 9215
rect 1144 9155 1196 9215
rect 1234 9155 1286 9215
rect 1544 9155 1596 9215
rect 1634 9155 1686 9215
rect 1944 9155 1996 9215
rect 2034 9155 2086 9215
rect 2344 9155 2396 9215
rect 2434 9155 2486 9215
rect 2744 9155 2796 9215
rect 34 8895 86 8955
rect 344 8895 396 8955
rect 434 8895 486 8955
rect 744 8895 796 8955
rect 834 8895 886 8955
rect 1144 8895 1196 8955
rect 1234 8895 1286 8955
rect 1544 8895 1596 8955
rect 1634 8895 1686 8955
rect 1944 8895 1996 8955
rect 2034 8895 2086 8955
rect 2344 8895 2396 8955
rect 2434 8895 2486 8955
rect 2744 8895 2796 8955
rect 2834 9155 2886 9215
rect 3144 9155 3196 9215
rect 3234 9155 3286 9215
rect 3544 9155 3596 9215
rect 3634 9155 3686 9215
rect 3944 9155 3996 9215
rect 4034 9155 4086 9215
rect 4344 9155 4396 9215
rect 4434 9155 4486 9215
rect 4744 9155 4796 9215
rect 4834 9155 4886 9215
rect 5144 9155 5196 9215
rect 5234 9155 5286 9215
rect 5544 9155 5596 9215
rect 5634 9155 5686 9215
rect 5944 9155 5996 9215
rect 2834 8895 2886 8955
rect 3144 8895 3196 8955
rect 3234 8895 3286 8955
rect 3544 8895 3596 8955
rect 3634 8895 3686 8955
rect 3944 8895 3996 8955
rect 4034 8895 4086 8955
rect 4344 8895 4396 8955
rect 4434 8895 4486 8955
rect 4744 8895 4796 8955
rect 4834 8895 4886 8955
rect 5144 8895 5196 8955
rect 5234 8895 5286 8955
rect 5544 8895 5596 8955
rect 5634 8895 5686 8955
rect 5944 8895 5996 8955
rect 6034 9155 6086 9215
rect 6344 9155 6396 9215
rect 6434 9155 6486 9215
rect 6744 9155 6796 9215
rect 6834 9155 6886 9215
rect 7144 9155 7196 9215
rect 7234 9155 7286 9215
rect 7544 9155 7596 9215
rect 6034 8895 6086 8955
rect 6344 8895 6396 8955
rect 6434 8895 6486 8955
rect 6744 8895 6796 8955
rect 6834 8895 6886 8955
rect 7144 8895 7196 8955
rect 7234 8895 7286 8955
rect 7544 8895 7596 8955
rect 7634 9155 7686 9215
rect 7944 9155 7996 9215
rect 8034 9155 8086 9215
rect 8344 9155 8396 9215
rect 8434 9155 8486 9215
rect 8744 9155 8796 9215
rect 8834 9155 8886 9215
rect 9144 9155 9196 9215
rect 9234 9155 9286 9215
rect 9544 9155 9596 9215
rect 9634 9155 9686 9215
rect 9944 9155 9996 9215
rect 10034 9155 10086 9215
rect 10344 9155 10396 9215
rect 10434 9155 10486 9215
rect 10744 9155 10796 9215
rect 10834 9155 10886 9215
rect 11144 9155 11196 9215
rect 11234 9155 11286 9215
rect 11544 9155 11596 9215
rect 11634 9155 11686 9215
rect 11944 9155 11996 9215
rect 12034 9155 12086 9215
rect 12344 9155 12396 9215
rect 12434 9155 12486 9215
rect 12744 9155 12796 9215
rect 12834 9155 12886 9215
rect 13144 9155 13196 9215
rect 7634 8895 7686 8955
rect 7944 8895 7996 8955
rect 8034 8895 8086 8955
rect 8344 8895 8396 8955
rect 8434 8895 8486 8955
rect 8744 8895 8796 8955
rect 8834 8895 8886 8955
rect 9144 8895 9196 8955
rect 9234 8895 9286 8955
rect 9544 8895 9596 8955
rect 9634 8895 9686 8955
rect 9944 8895 9996 8955
rect 10034 8895 10086 8955
rect 10344 8895 10396 8955
rect 10434 8895 10486 8955
rect 10744 8895 10796 8955
rect 10834 8895 10886 8955
rect 11144 8895 11196 8955
rect 11234 8895 11286 8955
rect 11544 8895 11596 8955
rect 11634 8895 11686 8955
rect 11944 8895 11996 8955
rect 12034 8895 12086 8955
rect 12344 8895 12396 8955
rect 12434 8895 12486 8955
rect 12744 8895 12796 8955
rect 12834 8895 12886 8955
rect 13144 8895 13196 8955
rect -366 8785 -330 8845
rect -330 8785 -314 8845
rect -56 8785 -4 8845
rect -366 8525 -330 8585
rect -330 8525 -314 8585
rect -56 8525 -4 8585
rect 34 8785 86 8845
rect 344 8785 396 8845
rect 434 8785 486 8845
rect 744 8785 796 8845
rect 834 8785 886 8845
rect 1144 8785 1196 8845
rect 1234 8785 1286 8845
rect 1544 8785 1596 8845
rect 1634 8785 1686 8845
rect 1944 8785 1996 8845
rect 2034 8785 2086 8845
rect 2344 8785 2396 8845
rect 2434 8785 2486 8845
rect 2744 8785 2796 8845
rect 2834 8785 2886 8845
rect 3144 8785 3196 8845
rect 34 8525 86 8585
rect 344 8525 396 8585
rect 434 8525 486 8585
rect 744 8525 796 8585
rect 834 8525 886 8585
rect 1144 8525 1196 8585
rect 1234 8525 1286 8585
rect 1544 8525 1596 8585
rect 1634 8525 1686 8585
rect 1944 8525 1996 8585
rect 2034 8525 2086 8585
rect 2344 8525 2396 8585
rect 2434 8525 2486 8585
rect 2744 8525 2796 8585
rect 2834 8525 2886 8585
rect 3144 8525 3196 8585
rect 3234 8785 3286 8845
rect 3544 8785 3596 8845
rect 3634 8785 3686 8845
rect 3944 8785 3996 8845
rect 4034 8785 4086 8845
rect 4344 8785 4396 8845
rect 4434 8785 4486 8845
rect 4744 8785 4796 8845
rect 4834 8785 4886 8845
rect 5144 8785 5196 8845
rect 5234 8785 5286 8845
rect 5544 8785 5596 8845
rect 5634 8785 5686 8845
rect 5944 8785 5996 8845
rect 3234 8525 3286 8585
rect 3544 8525 3596 8585
rect 3634 8525 3686 8585
rect 3944 8525 3996 8585
rect 4034 8525 4086 8585
rect 4344 8525 4396 8585
rect 4434 8525 4486 8585
rect 4744 8525 4796 8585
rect 4834 8525 4886 8585
rect 5144 8525 5196 8585
rect 5234 8525 5286 8585
rect 5544 8525 5596 8585
rect 5634 8525 5686 8585
rect 5944 8525 5996 8585
rect 6034 8785 6086 8845
rect 6344 8785 6396 8845
rect 6434 8785 6486 8845
rect 6744 8785 6796 8845
rect 6834 8785 6886 8845
rect 7144 8785 7196 8845
rect 7234 8785 7286 8845
rect 7544 8785 7596 8845
rect 7634 8785 7686 8845
rect 7944 8785 7996 8845
rect 6034 8525 6086 8585
rect 6344 8525 6396 8585
rect 6434 8525 6486 8585
rect 6744 8525 6796 8585
rect 6834 8525 6886 8585
rect 7144 8525 7196 8585
rect 7234 8525 7286 8585
rect 7544 8525 7596 8585
rect 7634 8525 7686 8585
rect 7944 8525 7996 8585
rect 8034 8785 8086 8845
rect 8344 8785 8396 8845
rect 8434 8785 8486 8845
rect 8744 8785 8796 8845
rect 8834 8785 8886 8845
rect 9144 8785 9196 8845
rect 9234 8785 9286 8845
rect 9544 8785 9596 8845
rect 9634 8785 9686 8845
rect 9944 8785 9996 8845
rect 10034 8785 10086 8845
rect 10344 8785 10396 8845
rect 10434 8785 10486 8845
rect 10744 8785 10796 8845
rect 10834 8785 10886 8845
rect 11144 8785 11196 8845
rect 11234 8785 11286 8845
rect 11544 8785 11596 8845
rect 11634 8785 11686 8845
rect 11944 8785 11996 8845
rect 12034 8785 12086 8845
rect 12344 8785 12396 8845
rect 12434 8785 12486 8845
rect 12744 8785 12796 8845
rect 12834 8785 12886 8845
rect 13144 8785 13196 8845
rect 8034 8525 8086 8585
rect 8344 8525 8396 8585
rect 8434 8525 8486 8585
rect 8744 8525 8796 8585
rect 8834 8525 8886 8585
rect 9144 8525 9196 8585
rect 9234 8525 9286 8585
rect 9544 8525 9596 8585
rect 9634 8525 9686 8585
rect 9944 8525 9996 8585
rect 10034 8525 10086 8585
rect 10344 8525 10396 8585
rect 10434 8525 10486 8585
rect 10744 8525 10796 8585
rect 10834 8525 10886 8585
rect 11144 8525 11196 8585
rect 11234 8525 11286 8585
rect 11544 8525 11596 8585
rect 11634 8525 11686 8585
rect 11944 8525 11996 8585
rect 12034 8525 12086 8585
rect 12344 8525 12396 8585
rect 12434 8525 12486 8585
rect 12744 8525 12796 8585
rect 12834 8525 12886 8585
rect 13144 8525 13196 8585
rect -366 8415 -330 8475
rect -330 8415 -314 8475
rect -56 8415 -4 8475
rect -366 8155 -330 8215
rect -330 8155 -314 8215
rect -56 8155 -4 8215
rect 34 8415 86 8475
rect 344 8415 396 8475
rect 434 8415 486 8475
rect 744 8415 796 8475
rect 834 8415 886 8475
rect 1144 8415 1196 8475
rect 1234 8415 1286 8475
rect 1544 8415 1596 8475
rect 1634 8415 1686 8475
rect 1944 8415 1996 8475
rect 2034 8415 2086 8475
rect 2344 8415 2396 8475
rect 2434 8415 2486 8475
rect 2744 8415 2796 8475
rect 2834 8415 2886 8475
rect 3144 8415 3196 8475
rect 34 8155 86 8215
rect 344 8155 396 8215
rect 434 8155 486 8215
rect 744 8155 796 8215
rect 834 8155 886 8215
rect 1144 8155 1196 8215
rect 1234 8155 1286 8215
rect 1544 8155 1596 8215
rect 1634 8155 1686 8215
rect 1944 8155 1996 8215
rect 2034 8155 2086 8215
rect 2344 8155 2396 8215
rect 2434 8155 2486 8215
rect 2744 8155 2796 8215
rect 2834 8155 2886 8215
rect 3144 8155 3196 8215
rect 3234 8415 3286 8475
rect 3544 8415 3596 8475
rect 3634 8415 3686 8475
rect 3944 8415 3996 8475
rect 4034 8415 4086 8475
rect 4344 8415 4396 8475
rect 4434 8415 4486 8475
rect 4744 8415 4796 8475
rect 4834 8415 4886 8475
rect 5144 8415 5196 8475
rect 5234 8415 5286 8475
rect 5544 8415 5596 8475
rect 5634 8415 5686 8475
rect 5944 8415 5996 8475
rect 3234 8155 3286 8215
rect 3544 8155 3596 8215
rect 3634 8155 3686 8215
rect 3944 8155 3996 8215
rect 4034 8155 4086 8215
rect 4344 8155 4396 8215
rect 4434 8155 4486 8215
rect 4744 8155 4796 8215
rect 4834 8155 4886 8215
rect 5144 8155 5196 8215
rect 5234 8155 5286 8215
rect 5544 8155 5596 8215
rect 5634 8155 5686 8215
rect 5944 8155 5996 8215
rect 6034 8415 6086 8475
rect 6344 8415 6396 8475
rect 6434 8415 6486 8475
rect 6744 8415 6796 8475
rect 6834 8415 6886 8475
rect 7144 8415 7196 8475
rect 7234 8415 7286 8475
rect 7544 8415 7596 8475
rect 7634 8415 7686 8475
rect 7944 8415 7996 8475
rect 6034 8155 6086 8215
rect 6344 8155 6396 8215
rect 6434 8155 6486 8215
rect 6744 8155 6796 8215
rect 6834 8155 6886 8215
rect 7144 8155 7196 8215
rect 7234 8155 7286 8215
rect 7544 8155 7596 8215
rect 7634 8155 7686 8215
rect 7944 8155 7996 8215
rect 8034 8415 8086 8475
rect 8344 8415 8396 8475
rect 8434 8415 8486 8475
rect 8744 8415 8796 8475
rect 8834 8415 8886 8475
rect 9144 8415 9196 8475
rect 9234 8415 9286 8475
rect 9544 8415 9596 8475
rect 9634 8415 9686 8475
rect 9944 8415 9996 8475
rect 10034 8415 10086 8475
rect 10344 8415 10396 8475
rect 10434 8415 10486 8475
rect 10744 8415 10796 8475
rect 10834 8415 10886 8475
rect 11144 8415 11196 8475
rect 11234 8415 11286 8475
rect 11544 8415 11596 8475
rect 11634 8415 11686 8475
rect 11944 8415 11996 8475
rect 12034 8415 12086 8475
rect 12344 8415 12396 8475
rect 12434 8415 12486 8475
rect 12744 8415 12796 8475
rect 12834 8415 12886 8475
rect 13144 8415 13196 8475
rect 8034 8155 8086 8215
rect 8344 8155 8396 8215
rect 8434 8155 8486 8215
rect 8744 8155 8796 8215
rect 8834 8155 8886 8215
rect 9144 8155 9196 8215
rect 9234 8155 9286 8215
rect 9544 8155 9596 8215
rect 9634 8155 9686 8215
rect 9944 8155 9996 8215
rect 10034 8155 10086 8215
rect 10344 8155 10396 8215
rect 10434 8155 10486 8215
rect 10744 8155 10796 8215
rect 10834 8155 10886 8215
rect 11144 8155 11196 8215
rect 11234 8155 11286 8215
rect 11544 8155 11596 8215
rect 11634 8155 11686 8215
rect 11944 8155 11996 8215
rect 12034 8155 12086 8215
rect 12344 8155 12396 8215
rect 12434 8155 12486 8215
rect 12744 8155 12796 8215
rect 12834 8155 12886 8215
rect 13144 8155 13196 8215
rect -366 8045 -330 8105
rect -330 8045 -314 8105
rect -56 8045 -4 8105
rect -366 7785 -330 7845
rect -330 7785 -314 7845
rect -56 7785 -4 7845
rect 34 8045 86 8105
rect 344 8045 396 8105
rect 434 8045 486 8105
rect 744 8045 796 8105
rect 834 8045 886 8105
rect 1144 8045 1196 8105
rect 1234 8045 1286 8105
rect 1544 8045 1596 8105
rect 1634 8045 1686 8105
rect 1944 8045 1996 8105
rect 2034 8045 2086 8105
rect 2344 8045 2396 8105
rect 2434 8045 2486 8105
rect 2744 8045 2796 8105
rect 2834 8045 2886 8105
rect 3144 8045 3196 8105
rect 34 7785 86 7845
rect 344 7785 396 7845
rect 434 7785 486 7845
rect 744 7785 796 7845
rect 834 7785 886 7845
rect 1144 7785 1196 7845
rect 1234 7785 1286 7845
rect 1544 7785 1596 7845
rect 1634 7785 1686 7845
rect 1944 7785 1996 7845
rect 2034 7785 2086 7845
rect 2344 7785 2396 7845
rect 2434 7785 2486 7845
rect 2744 7785 2796 7845
rect 2834 7785 2886 7845
rect 3144 7785 3196 7845
rect 3234 8045 3286 8105
rect 3544 8045 3596 8105
rect 3634 8045 3686 8105
rect 3944 8045 3996 8105
rect 4034 8045 4086 8105
rect 4344 8045 4396 8105
rect 4434 8045 4486 8105
rect 4744 8045 4796 8105
rect 4834 8045 4886 8105
rect 5144 8045 5196 8105
rect 5234 8045 5286 8105
rect 5544 8045 5596 8105
rect 5634 8045 5686 8105
rect 5944 8045 5996 8105
rect 3234 7785 3286 7845
rect 3544 7785 3596 7845
rect 3634 7785 3686 7845
rect 3944 7785 3996 7845
rect 4034 7785 4086 7845
rect 4344 7785 4396 7845
rect 4434 7785 4486 7845
rect 4744 7785 4796 7845
rect 4834 7785 4886 7845
rect 5144 7785 5196 7845
rect 5234 7785 5286 7845
rect 5544 7785 5596 7845
rect 5634 7785 5686 7845
rect 5944 7785 5996 7845
rect 6034 8045 6086 8105
rect 6344 8045 6396 8105
rect 6434 8045 6486 8105
rect 6744 8045 6796 8105
rect 6834 8045 6886 8105
rect 7144 8045 7196 8105
rect 7234 8045 7286 8105
rect 7544 8045 7596 8105
rect 7634 8045 7686 8105
rect 7944 8045 7996 8105
rect 8034 8045 8086 8105
rect 8344 8045 8396 8105
rect 8434 8045 8486 8105
rect 8744 8045 8796 8105
rect 8834 8045 8886 8105
rect 9144 8045 9196 8105
rect 9234 8045 9286 8105
rect 9544 8045 9596 8105
rect 9634 8045 9686 8105
rect 9944 8045 9996 8105
rect 10034 8045 10086 8105
rect 10344 8045 10396 8105
rect 10434 8045 10486 8105
rect 10744 8045 10796 8105
rect 10834 8045 10886 8105
rect 11144 8045 11196 8105
rect 11234 8045 11286 8105
rect 11544 8045 11596 8105
rect 11634 8045 11686 8105
rect 11944 8045 11996 8105
rect 12034 8045 12086 8105
rect 12344 8045 12396 8105
rect 12434 8045 12486 8105
rect 12744 8045 12796 8105
rect 12834 8045 12886 8105
rect 13144 8045 13196 8105
rect 6034 7785 6086 7845
rect 6344 7785 6396 7845
rect 6434 7785 6486 7845
rect 6744 7785 6796 7845
rect 6834 7785 6886 7845
rect 7144 7785 7196 7845
rect 7234 7785 7286 7845
rect 7544 7785 7596 7845
rect 7634 7785 7686 7845
rect 7944 7785 7996 7845
rect 8034 7785 8086 7845
rect 8344 7785 8396 7845
rect 8434 7785 8486 7845
rect 8744 7785 8796 7845
rect 8834 7785 8886 7845
rect 9144 7785 9196 7845
rect 9234 7785 9286 7845
rect 9544 7785 9596 7845
rect 9634 7785 9686 7845
rect 9944 7785 9996 7845
rect 10034 7785 10086 7845
rect 10344 7785 10396 7845
rect 10434 7785 10486 7845
rect 10744 7785 10796 7845
rect 10834 7785 10886 7845
rect 11144 7785 11196 7845
rect 11234 7785 11286 7845
rect 11544 7785 11596 7845
rect 11634 7785 11686 7845
rect 11944 7785 11996 7845
rect 12034 7785 12086 7845
rect 12344 7785 12396 7845
rect 12434 7785 12486 7845
rect 12744 7785 12796 7845
rect 12834 7785 12886 7845
rect 13144 7785 13196 7845
rect -366 7675 -330 7735
rect -330 7675 -314 7735
rect -56 7675 -4 7735
rect -366 7415 -330 7475
rect -330 7415 -314 7475
rect -56 7415 -4 7475
rect 34 7675 86 7735
rect 344 7675 396 7735
rect 434 7675 486 7735
rect 744 7675 796 7735
rect 834 7675 886 7735
rect 1144 7675 1196 7735
rect 1234 7675 1286 7735
rect 1544 7675 1596 7735
rect 1634 7675 1686 7735
rect 1944 7675 1996 7735
rect 2034 7675 2086 7735
rect 2344 7675 2396 7735
rect 2434 7675 2486 7735
rect 2744 7675 2796 7735
rect 2834 7675 2886 7735
rect 3144 7675 3196 7735
rect 34 7415 86 7475
rect 344 7415 396 7475
rect 434 7415 486 7475
rect 744 7415 796 7475
rect 834 7415 886 7475
rect 1144 7415 1196 7475
rect 1234 7415 1286 7475
rect 1544 7415 1596 7475
rect 1634 7415 1686 7475
rect 1944 7415 1996 7475
rect 2034 7415 2086 7475
rect 2344 7415 2396 7475
rect 2434 7415 2486 7475
rect 2744 7415 2796 7475
rect 2834 7415 2886 7475
rect 3144 7415 3196 7475
rect 3234 7675 3286 7735
rect 3544 7675 3596 7735
rect 3634 7675 3686 7735
rect 3944 7675 3996 7735
rect 4034 7675 4086 7735
rect 4344 7675 4396 7735
rect 4434 7675 4486 7735
rect 4744 7675 4796 7735
rect 4834 7675 4886 7735
rect 5144 7675 5196 7735
rect 5234 7675 5286 7735
rect 5544 7675 5596 7735
rect 5634 7675 5686 7735
rect 5944 7675 5996 7735
rect 3234 7415 3286 7475
rect 3544 7415 3596 7475
rect 3634 7415 3686 7475
rect 3944 7415 3996 7475
rect 4034 7415 4086 7475
rect 4344 7415 4396 7475
rect 4434 7415 4486 7475
rect 4744 7415 4796 7475
rect 4834 7415 4886 7475
rect 5144 7415 5196 7475
rect 5234 7415 5286 7475
rect 5544 7415 5596 7475
rect 5634 7415 5686 7475
rect 5944 7415 5996 7475
rect 6034 7675 6086 7735
rect 6344 7675 6396 7735
rect 6434 7675 6486 7735
rect 6744 7675 6796 7735
rect 6834 7675 6886 7735
rect 7144 7675 7196 7735
rect 7234 7675 7286 7735
rect 7544 7675 7596 7735
rect 7634 7675 7686 7735
rect 7944 7675 7996 7735
rect 8034 7675 8086 7735
rect 8344 7675 8396 7735
rect 8434 7675 8486 7735
rect 8744 7675 8796 7735
rect 8834 7675 8886 7735
rect 9144 7675 9196 7735
rect 9234 7675 9286 7735
rect 9544 7675 9596 7735
rect 9634 7675 9686 7735
rect 9944 7675 9996 7735
rect 10034 7675 10086 7735
rect 10344 7675 10396 7735
rect 10434 7675 10486 7735
rect 10744 7675 10796 7735
rect 10834 7675 10886 7735
rect 11144 7675 11196 7735
rect 11234 7675 11286 7735
rect 11544 7675 11596 7735
rect 11634 7675 11686 7735
rect 11944 7675 11996 7735
rect 12034 7675 12086 7735
rect 12344 7675 12396 7735
rect 12434 7675 12486 7735
rect 12744 7675 12796 7735
rect 12834 7675 12886 7735
rect 13144 7675 13196 7735
rect 6034 7415 6086 7475
rect 6344 7415 6396 7475
rect 6434 7415 6486 7475
rect 6744 7415 6796 7475
rect 6834 7415 6886 7475
rect 7144 7415 7196 7475
rect 7234 7415 7286 7475
rect 7544 7415 7596 7475
rect 7634 7415 7686 7475
rect 7944 7415 7996 7475
rect 8034 7415 8086 7475
rect 8344 7415 8396 7475
rect 8434 7415 8486 7475
rect 8744 7415 8796 7475
rect 8834 7415 8886 7475
rect 9144 7415 9196 7475
rect 9234 7415 9286 7475
rect 9544 7415 9596 7475
rect 9634 7415 9686 7475
rect 9944 7415 9996 7475
rect 10034 7415 10086 7475
rect 10344 7415 10396 7475
rect 10434 7415 10486 7475
rect 10744 7415 10796 7475
rect 10834 7415 10886 7475
rect 11144 7415 11196 7475
rect 11234 7415 11286 7475
rect 11544 7415 11596 7475
rect 11634 7415 11686 7475
rect 11944 7415 11996 7475
rect 12034 7415 12086 7475
rect 12344 7415 12396 7475
rect 12434 7415 12486 7475
rect 12744 7415 12796 7475
rect 12834 7415 12886 7475
rect 13144 7415 13196 7475
rect -366 7305 -330 7365
rect -330 7305 -314 7365
rect -56 7305 -4 7365
rect -366 7045 -330 7105
rect -330 7045 -314 7105
rect -56 7045 -4 7105
rect 34 7305 86 7365
rect 344 7305 396 7365
rect 434 7305 486 7365
rect 744 7305 796 7365
rect 834 7305 886 7365
rect 1144 7305 1196 7365
rect 1234 7305 1286 7365
rect 1544 7305 1596 7365
rect 1634 7305 1686 7365
rect 1944 7305 1996 7365
rect 2034 7305 2086 7365
rect 2344 7305 2396 7365
rect 2434 7305 2486 7365
rect 2744 7305 2796 7365
rect 2834 7305 2886 7365
rect 3144 7305 3196 7365
rect 34 7045 86 7105
rect 344 7045 396 7105
rect 434 7045 486 7105
rect 744 7045 796 7105
rect 834 7045 886 7105
rect 1144 7045 1196 7105
rect 1234 7045 1286 7105
rect 1544 7045 1596 7105
rect 1634 7045 1686 7105
rect 1944 7045 1996 7105
rect 2034 7045 2086 7105
rect 2344 7045 2396 7105
rect 2434 7045 2486 7105
rect 2744 7045 2796 7105
rect 2834 7045 2886 7105
rect 3144 7045 3196 7105
rect 3234 7305 3286 7365
rect 3544 7305 3596 7365
rect 3634 7305 3686 7365
rect 3944 7305 3996 7365
rect 4034 7305 4086 7365
rect 4344 7305 4396 7365
rect 4434 7305 4486 7365
rect 4744 7305 4796 7365
rect 4834 7305 4886 7365
rect 5144 7305 5196 7365
rect 5234 7305 5286 7365
rect 5544 7305 5596 7365
rect 5634 7305 5686 7365
rect 5944 7305 5996 7365
rect 3234 7045 3286 7105
rect 3544 7045 3596 7105
rect 3634 7045 3686 7105
rect 3944 7045 3996 7105
rect 4034 7045 4086 7105
rect 4344 7045 4396 7105
rect 4434 7045 4486 7105
rect 4744 7045 4796 7105
rect 4834 7045 4886 7105
rect 5144 7045 5196 7105
rect 5234 7045 5286 7105
rect 5544 7045 5596 7105
rect 5634 7045 5686 7105
rect 5944 7045 5996 7105
rect 6034 7305 6086 7365
rect 6344 7305 6396 7365
rect 6434 7305 6486 7365
rect 6744 7305 6796 7365
rect 6834 7305 6886 7365
rect 7144 7305 7196 7365
rect 7234 7305 7286 7365
rect 7544 7305 7596 7365
rect 7634 7305 7686 7365
rect 7944 7305 7996 7365
rect 8034 7305 8086 7365
rect 8344 7305 8396 7365
rect 8434 7305 8486 7365
rect 8744 7305 8796 7365
rect 8834 7305 8886 7365
rect 9144 7305 9196 7365
rect 9234 7305 9286 7365
rect 9544 7305 9596 7365
rect 9634 7305 9686 7365
rect 9944 7305 9996 7365
rect 10034 7305 10086 7365
rect 10344 7305 10396 7365
rect 10434 7305 10486 7365
rect 10744 7305 10796 7365
rect 10834 7305 10886 7365
rect 11144 7305 11196 7365
rect 11234 7305 11286 7365
rect 11544 7305 11596 7365
rect 11634 7305 11686 7365
rect 11944 7305 11996 7365
rect 12034 7305 12086 7365
rect 12344 7305 12396 7365
rect 12434 7305 12486 7365
rect 12744 7305 12796 7365
rect 12834 7305 12886 7365
rect 13144 7305 13196 7365
rect 6034 7045 6086 7105
rect 6344 7045 6396 7105
rect 6434 7045 6486 7105
rect 6744 7045 6796 7105
rect 6834 7045 6886 7105
rect 7144 7045 7196 7105
rect 7234 7045 7286 7105
rect 7544 7045 7596 7105
rect 7634 7045 7686 7105
rect 7944 7045 7996 7105
rect 8034 7045 8086 7105
rect 8344 7045 8396 7105
rect 8434 7045 8486 7105
rect 8744 7045 8796 7105
rect 8834 7045 8886 7105
rect 9144 7045 9196 7105
rect 9234 7045 9286 7105
rect 9544 7045 9596 7105
rect 9634 7045 9686 7105
rect 9944 7045 9996 7105
rect 10034 7045 10086 7105
rect 10344 7045 10396 7105
rect 10434 7045 10486 7105
rect 10744 7045 10796 7105
rect 10834 7045 10886 7105
rect 11144 7045 11196 7105
rect 11234 7045 11286 7105
rect 11544 7045 11596 7105
rect 11634 7045 11686 7105
rect 11944 7045 11996 7105
rect 12034 7045 12086 7105
rect 12344 7045 12396 7105
rect 12434 7045 12486 7105
rect 12744 7045 12796 7105
rect 12834 7045 12886 7105
rect 13144 7045 13196 7105
rect -366 6935 -330 6995
rect -330 6935 -314 6995
rect -56 6935 -4 6995
rect -366 6675 -330 6735
rect -330 6675 -314 6735
rect -56 6675 -4 6735
rect 34 6935 86 6995
rect 344 6935 396 6995
rect 434 6935 486 6995
rect 744 6935 796 6995
rect 834 6935 886 6995
rect 1144 6935 1196 6995
rect 1234 6935 1286 6995
rect 1544 6935 1596 6995
rect 1634 6935 1686 6995
rect 1944 6935 1996 6995
rect 2034 6935 2086 6995
rect 2344 6935 2396 6995
rect 2434 6935 2486 6995
rect 2744 6935 2796 6995
rect 2834 6935 2886 6995
rect 3144 6935 3196 6995
rect 34 6675 86 6735
rect 344 6675 396 6735
rect 434 6675 486 6735
rect 744 6675 796 6735
rect 834 6675 886 6735
rect 1144 6675 1196 6735
rect 1234 6675 1286 6735
rect 1544 6675 1596 6735
rect 1634 6675 1686 6735
rect 1944 6675 1996 6735
rect 2034 6675 2086 6735
rect 2344 6675 2396 6735
rect 2434 6675 2486 6735
rect 2744 6675 2796 6735
rect 2834 6675 2886 6735
rect 3144 6675 3196 6735
rect 3234 6935 3286 6995
rect 3544 6935 3596 6995
rect 3634 6935 3686 6995
rect 3944 6935 3996 6995
rect 4034 6935 4086 6995
rect 4344 6935 4396 6995
rect 4434 6935 4486 6995
rect 4744 6935 4796 6995
rect 4834 6935 4886 6995
rect 5144 6935 5196 6995
rect 5234 6935 5286 6995
rect 5544 6935 5596 6995
rect 5634 6935 5686 6995
rect 5944 6935 5996 6995
rect 3234 6675 3286 6735
rect 3544 6675 3596 6735
rect 3634 6675 3686 6735
rect 3944 6675 3996 6735
rect 4034 6675 4086 6735
rect 4344 6675 4396 6735
rect 4434 6675 4486 6735
rect 4744 6675 4796 6735
rect 4834 6675 4886 6735
rect 5144 6675 5196 6735
rect 5234 6675 5286 6735
rect 5544 6675 5596 6735
rect 5634 6675 5686 6735
rect 5944 6675 5996 6735
rect 6034 6935 6086 6995
rect 6344 6935 6396 6995
rect 6434 6935 6486 6995
rect 6744 6935 6796 6995
rect 6834 6935 6886 6995
rect 7144 6935 7196 6995
rect 7234 6935 7286 6995
rect 7544 6935 7596 6995
rect 7634 6935 7686 6995
rect 7944 6935 7996 6995
rect 8034 6935 8086 6995
rect 8344 6935 8396 6995
rect 8434 6935 8486 6995
rect 8744 6935 8796 6995
rect 8834 6935 8886 6995
rect 9144 6935 9196 6995
rect 9234 6935 9286 6995
rect 9544 6935 9596 6995
rect 9634 6935 9686 6995
rect 9944 6935 9996 6995
rect 10034 6935 10086 6995
rect 10344 6935 10396 6995
rect 10434 6935 10486 6995
rect 10744 6935 10796 6995
rect 10834 6935 10886 6995
rect 11144 6935 11196 6995
rect 11234 6935 11286 6995
rect 11544 6935 11596 6995
rect 11634 6935 11686 6995
rect 11944 6935 11996 6995
rect 12034 6935 12086 6995
rect 12344 6935 12396 6995
rect 12434 6935 12486 6995
rect 12744 6935 12796 6995
rect 12834 6935 12886 6995
rect 13144 6935 13196 6995
rect 6034 6675 6086 6735
rect 6344 6675 6396 6735
rect 6434 6675 6486 6735
rect 6744 6675 6796 6735
rect 6834 6675 6886 6735
rect 7144 6675 7196 6735
rect 7234 6675 7286 6735
rect 7544 6675 7596 6735
rect 7634 6675 7686 6735
rect 7944 6675 7996 6735
rect 8034 6675 8086 6735
rect 8344 6675 8396 6735
rect 8434 6675 8486 6735
rect 8744 6675 8796 6735
rect 8834 6675 8886 6735
rect 9144 6675 9196 6735
rect 9234 6675 9286 6735
rect 9544 6675 9596 6735
rect 9634 6675 9686 6735
rect 9944 6675 9996 6735
rect 10034 6675 10086 6735
rect 10344 6675 10396 6735
rect 10434 6675 10486 6735
rect 10744 6675 10796 6735
rect 10834 6675 10886 6735
rect 11144 6675 11196 6735
rect 11234 6675 11286 6735
rect 11544 6675 11596 6735
rect 11634 6675 11686 6735
rect 11944 6675 11996 6735
rect 12034 6675 12086 6735
rect 12344 6675 12396 6735
rect 12434 6675 12486 6735
rect 12744 6675 12796 6735
rect 12834 6675 12886 6735
rect 13144 6675 13196 6735
rect -366 6565 -330 6625
rect -330 6565 -314 6625
rect -56 6565 -4 6625
rect -366 6305 -330 6365
rect -330 6305 -314 6365
rect -56 6305 -4 6365
rect 34 6565 86 6625
rect 344 6565 396 6625
rect 434 6565 486 6625
rect 744 6565 796 6625
rect 834 6565 886 6625
rect 1144 6565 1196 6625
rect 1234 6565 1286 6625
rect 1544 6565 1596 6625
rect 1634 6565 1686 6625
rect 1944 6565 1996 6625
rect 2034 6565 2086 6625
rect 2344 6565 2396 6625
rect 2434 6565 2486 6625
rect 2744 6565 2796 6625
rect 2834 6565 2886 6625
rect 3144 6565 3196 6625
rect 34 6305 86 6365
rect 344 6305 396 6365
rect 434 6305 486 6365
rect 744 6305 796 6365
rect 834 6305 886 6365
rect 1144 6305 1196 6365
rect 1234 6305 1286 6365
rect 1544 6305 1596 6365
rect 1634 6305 1686 6365
rect 1944 6305 1996 6365
rect 2034 6305 2086 6365
rect 2344 6305 2396 6365
rect 2434 6305 2486 6365
rect 2744 6305 2796 6365
rect 2834 6305 2886 6365
rect 3144 6305 3196 6365
rect 3234 6565 3286 6625
rect 3544 6565 3596 6625
rect 3634 6565 3686 6625
rect 3944 6565 3996 6625
rect 4034 6565 4086 6625
rect 4344 6565 4396 6625
rect 4434 6565 4486 6625
rect 4744 6565 4796 6625
rect 4834 6565 4886 6625
rect 5144 6565 5196 6625
rect 5234 6565 5286 6625
rect 5544 6565 5596 6625
rect 5634 6565 5686 6625
rect 5944 6565 5996 6625
rect 3234 6305 3286 6365
rect 3544 6305 3596 6365
rect 3634 6305 3686 6365
rect 3944 6305 3996 6365
rect 4034 6305 4086 6365
rect 4344 6305 4396 6365
rect 4434 6305 4486 6365
rect 4744 6305 4796 6365
rect 4834 6305 4886 6365
rect 5144 6305 5196 6365
rect 5234 6305 5286 6365
rect 5544 6305 5596 6365
rect 5634 6305 5686 6365
rect 5944 6305 5996 6365
rect 6034 6565 6086 6625
rect 6344 6565 6396 6625
rect 6434 6565 6486 6625
rect 6744 6565 6796 6625
rect 6834 6565 6886 6625
rect 7144 6565 7196 6625
rect 7234 6565 7286 6625
rect 7544 6565 7596 6625
rect 7634 6565 7686 6625
rect 7944 6565 7996 6625
rect 8034 6565 8086 6625
rect 8344 6565 8396 6625
rect 8434 6565 8486 6625
rect 8744 6565 8796 6625
rect 8834 6565 8886 6625
rect 9144 6565 9196 6625
rect 9234 6565 9286 6625
rect 9544 6565 9596 6625
rect 9634 6565 9686 6625
rect 9944 6565 9996 6625
rect 10034 6565 10086 6625
rect 10344 6565 10396 6625
rect 10434 6565 10486 6625
rect 10744 6565 10796 6625
rect 10834 6565 10886 6625
rect 11144 6565 11196 6625
rect 11234 6565 11286 6625
rect 11544 6565 11596 6625
rect 11634 6565 11686 6625
rect 11944 6565 11996 6625
rect 12034 6565 12086 6625
rect 12344 6565 12396 6625
rect 12434 6565 12486 6625
rect 12744 6565 12796 6625
rect 12834 6565 12886 6625
rect 13144 6565 13196 6625
rect 6034 6305 6086 6365
rect 6344 6305 6396 6365
rect 6434 6305 6486 6365
rect 6744 6305 6796 6365
rect 6834 6305 6886 6365
rect 7144 6305 7196 6365
rect 7234 6305 7286 6365
rect 7544 6305 7596 6365
rect 7634 6305 7686 6365
rect 7944 6305 7996 6365
rect 8034 6305 8086 6365
rect 8344 6305 8396 6365
rect 8434 6305 8486 6365
rect 8744 6305 8796 6365
rect 8834 6305 8886 6365
rect 9144 6305 9196 6365
rect 9234 6305 9286 6365
rect 9544 6305 9596 6365
rect 9634 6305 9686 6365
rect 9944 6305 9996 6365
rect 10034 6305 10086 6365
rect 10344 6305 10396 6365
rect 10434 6305 10486 6365
rect 10744 6305 10796 6365
rect 10834 6305 10886 6365
rect 11144 6305 11196 6365
rect 11234 6305 11286 6365
rect 11544 6305 11596 6365
rect 11634 6305 11686 6365
rect 11944 6305 11996 6365
rect 12034 6305 12086 6365
rect 12344 6305 12396 6365
rect 12434 6305 12486 6365
rect 12744 6305 12796 6365
rect 12834 6305 12886 6365
rect 13144 6305 13196 6365
rect -366 6195 -330 6255
rect -330 6195 -314 6255
rect -56 6195 -4 6255
rect -366 5935 -330 5995
rect -330 5935 -314 5995
rect -56 5935 -4 5995
rect 34 6195 86 6255
rect 344 6195 396 6255
rect 434 6195 486 6255
rect 744 6195 796 6255
rect 834 6195 886 6255
rect 1144 6195 1196 6255
rect 1234 6195 1286 6255
rect 1544 6195 1596 6255
rect 1634 6195 1686 6255
rect 1944 6195 1996 6255
rect 2034 6195 2086 6255
rect 2344 6195 2396 6255
rect 2434 6195 2486 6255
rect 2744 6195 2796 6255
rect 2834 6195 2886 6255
rect 3144 6195 3196 6255
rect 34 5935 86 5995
rect 344 5935 396 5995
rect 434 5935 486 5995
rect 744 5935 796 5995
rect 834 5935 886 5995
rect 1144 5935 1196 5995
rect 1234 5935 1286 5995
rect 1544 5935 1596 5995
rect 1634 5935 1686 5995
rect 1944 5935 1996 5995
rect 2034 5935 2086 5995
rect 2344 5935 2396 5995
rect 2434 5935 2486 5995
rect 2744 5935 2796 5995
rect 2834 5935 2886 5995
rect 3144 5935 3196 5995
rect 3234 6195 3286 6255
rect 3544 6195 3596 6255
rect 3634 6195 3686 6255
rect 3944 6195 3996 6255
rect 4034 6195 4086 6255
rect 4344 6195 4396 6255
rect 4434 6195 4486 6255
rect 4744 6195 4796 6255
rect 4834 6195 4886 6255
rect 5144 6195 5196 6255
rect 5234 6195 5286 6255
rect 5544 6195 5596 6255
rect 5634 6195 5686 6255
rect 5944 6195 5996 6255
rect 6034 6195 6086 6255
rect 6344 6195 6396 6255
rect 6434 6195 6486 6255
rect 6744 6195 6796 6255
rect 6834 6195 6886 6255
rect 7144 6195 7196 6255
rect 7234 6195 7286 6255
rect 7544 6195 7596 6255
rect 7634 6195 7686 6255
rect 7944 6195 7996 6255
rect 8034 6195 8086 6255
rect 8344 6195 8396 6255
rect 8434 6195 8486 6255
rect 8744 6195 8796 6255
rect 8834 6195 8886 6255
rect 9144 6195 9196 6255
rect 9234 6195 9286 6255
rect 9544 6195 9596 6255
rect 9634 6195 9686 6255
rect 9944 6195 9996 6255
rect 10034 6195 10086 6255
rect 10344 6195 10396 6255
rect 10434 6195 10486 6255
rect 10744 6195 10796 6255
rect 10834 6195 10886 6255
rect 11144 6195 11196 6255
rect 11234 6195 11286 6255
rect 11544 6195 11596 6255
rect 11634 6195 11686 6255
rect 11944 6195 11996 6255
rect 12034 6195 12086 6255
rect 12344 6195 12396 6255
rect 12434 6195 12486 6255
rect 12744 6195 12796 6255
rect 12834 6195 12886 6255
rect 13144 6195 13196 6255
rect 3234 5935 3286 5995
rect 3544 5935 3596 5995
rect 3634 5935 3686 5995
rect 3944 5935 3996 5995
rect 4034 5935 4086 5995
rect 4344 5935 4396 5995
rect 4434 5935 4486 5995
rect 4744 5935 4796 5995
rect 4834 5935 4886 5995
rect 5144 5935 5196 5995
rect 5234 5935 5286 5995
rect 5544 5935 5596 5995
rect 5634 5935 5686 5995
rect 5944 5935 5996 5995
rect 6034 5935 6086 5995
rect 6344 5935 6396 5995
rect 6434 5935 6486 5995
rect 6744 5935 6796 5995
rect 6834 5935 6886 5995
rect 7144 5935 7196 5995
rect 7234 5935 7286 5995
rect 7544 5935 7596 5995
rect 7634 5935 7686 5995
rect 7944 5935 7996 5995
rect 8034 5935 8086 5995
rect 8344 5935 8396 5995
rect 8434 5935 8486 5995
rect 8744 5935 8796 5995
rect 8834 5935 8886 5995
rect 9144 5935 9196 5995
rect 9234 5935 9286 5995
rect 9544 5935 9596 5995
rect 9634 5935 9686 5995
rect 9944 5935 9996 5995
rect 10034 5935 10086 5995
rect 10344 5935 10396 5995
rect 10434 5935 10486 5995
rect 10744 5935 10796 5995
rect 10834 5935 10886 5995
rect 11144 5935 11196 5995
rect 11234 5935 11286 5995
rect 11544 5935 11596 5995
rect 11634 5935 11686 5995
rect 11944 5935 11996 5995
rect 12034 5935 12086 5995
rect 12344 5935 12396 5995
rect 12434 5935 12486 5995
rect 12744 5935 12796 5995
rect 12834 5935 12886 5995
rect 13144 5935 13196 5995
rect -366 5825 -330 5885
rect -330 5825 -314 5885
rect -56 5825 -4 5885
rect -366 5565 -330 5625
rect -330 5565 -314 5625
rect -56 5565 -4 5625
rect 34 5825 86 5885
rect 344 5825 396 5885
rect 434 5825 486 5885
rect 744 5825 796 5885
rect 834 5825 886 5885
rect 1144 5825 1196 5885
rect 1234 5825 1286 5885
rect 1544 5825 1596 5885
rect 1634 5825 1686 5885
rect 1944 5825 1996 5885
rect 2034 5825 2086 5885
rect 2344 5825 2396 5885
rect 2434 5825 2486 5885
rect 2744 5825 2796 5885
rect 2834 5825 2886 5885
rect 3144 5825 3196 5885
rect 34 5565 86 5625
rect 344 5565 396 5625
rect 434 5565 486 5625
rect 744 5565 796 5625
rect 834 5565 886 5625
rect 1144 5565 1196 5625
rect 1234 5565 1286 5625
rect 1544 5565 1596 5625
rect 1634 5565 1686 5625
rect 1944 5565 1996 5625
rect 2034 5565 2086 5625
rect 2344 5565 2396 5625
rect 2434 5565 2486 5625
rect 2744 5565 2796 5625
rect 2834 5565 2886 5625
rect 3144 5565 3196 5625
rect 3234 5825 3286 5885
rect 3544 5825 3596 5885
rect 3634 5825 3686 5885
rect 3944 5825 3996 5885
rect 4034 5825 4086 5885
rect 4344 5825 4396 5885
rect 4434 5825 4486 5885
rect 4744 5825 4796 5885
rect 4834 5825 4886 5885
rect 5144 5825 5196 5885
rect 5234 5825 5286 5885
rect 5544 5825 5596 5885
rect 5634 5825 5686 5885
rect 5944 5825 5996 5885
rect 6034 5825 6086 5885
rect 6344 5825 6396 5885
rect 6434 5825 6486 5885
rect 6744 5825 6796 5885
rect 6834 5825 6886 5885
rect 7144 5825 7196 5885
rect 7234 5825 7286 5885
rect 7544 5825 7596 5885
rect 7634 5825 7686 5885
rect 7944 5825 7996 5885
rect 8034 5825 8086 5885
rect 8344 5825 8396 5885
rect 8434 5825 8486 5885
rect 8744 5825 8796 5885
rect 8834 5825 8886 5885
rect 9144 5825 9196 5885
rect 9234 5825 9286 5885
rect 9544 5825 9596 5885
rect 9634 5825 9686 5885
rect 9944 5825 9996 5885
rect 10034 5825 10086 5885
rect 10344 5825 10396 5885
rect 10434 5825 10486 5885
rect 10744 5825 10796 5885
rect 10834 5825 10886 5885
rect 11144 5825 11196 5885
rect 11234 5825 11286 5885
rect 11544 5825 11596 5885
rect 11634 5825 11686 5885
rect 11944 5825 11996 5885
rect 12034 5825 12086 5885
rect 12344 5825 12396 5885
rect 12434 5825 12486 5885
rect 12744 5825 12796 5885
rect 12834 5825 12886 5885
rect 13144 5825 13196 5885
rect 3234 5565 3286 5625
rect 3544 5565 3596 5625
rect 3634 5565 3686 5625
rect 3944 5565 3996 5625
rect 4034 5565 4086 5625
rect 4344 5565 4396 5625
rect 4434 5565 4486 5625
rect 4744 5565 4796 5625
rect 4834 5565 4886 5625
rect 5144 5565 5196 5625
rect 5234 5565 5286 5625
rect 5544 5565 5596 5625
rect 5634 5565 5686 5625
rect 5944 5565 5996 5625
rect 6034 5565 6086 5625
rect 6344 5565 6396 5625
rect 6434 5565 6486 5625
rect 6744 5565 6796 5625
rect 6834 5565 6886 5625
rect 7144 5565 7196 5625
rect 7234 5565 7286 5625
rect 7544 5565 7596 5625
rect 7634 5565 7686 5625
rect 7944 5565 7996 5625
rect 8034 5565 8086 5625
rect 8344 5565 8396 5625
rect 8434 5565 8486 5625
rect 8744 5565 8796 5625
rect 8834 5565 8886 5625
rect 9144 5565 9196 5625
rect 9234 5565 9286 5625
rect 9544 5565 9596 5625
rect 9634 5565 9686 5625
rect 9944 5565 9996 5625
rect 10034 5565 10086 5625
rect 10344 5565 10396 5625
rect 10434 5565 10486 5625
rect 10744 5565 10796 5625
rect 10834 5565 10886 5625
rect 11144 5565 11196 5625
rect 11234 5565 11286 5625
rect 11544 5565 11596 5625
rect 11634 5565 11686 5625
rect 11944 5565 11996 5625
rect 12034 5565 12086 5625
rect 12344 5565 12396 5625
rect 12434 5565 12486 5625
rect 12744 5565 12796 5625
rect 12834 5565 12886 5625
rect 13144 5565 13196 5625
rect -366 5455 -330 5515
rect -330 5455 -314 5515
rect -56 5455 -4 5515
rect -366 5195 -330 5255
rect -330 5195 -314 5255
rect -56 5195 -4 5255
rect 34 5455 86 5515
rect 344 5455 396 5515
rect 434 5455 486 5515
rect 744 5455 796 5515
rect 834 5455 886 5515
rect 1144 5455 1196 5515
rect 1234 5455 1286 5515
rect 1544 5455 1596 5515
rect 1634 5455 1686 5515
rect 1944 5455 1996 5515
rect 2034 5455 2086 5515
rect 2344 5455 2396 5515
rect 2434 5455 2486 5515
rect 2744 5455 2796 5515
rect 2834 5455 2886 5515
rect 3144 5455 3196 5515
rect 34 5195 86 5255
rect 344 5195 396 5255
rect 434 5195 486 5255
rect 744 5195 796 5255
rect 834 5195 886 5255
rect 1144 5195 1196 5255
rect 1234 5195 1286 5255
rect 1544 5195 1596 5255
rect 1634 5195 1686 5255
rect 1944 5195 1996 5255
rect 2034 5195 2086 5255
rect 2344 5195 2396 5255
rect 2434 5195 2486 5255
rect 2744 5195 2796 5255
rect 2834 5195 2886 5255
rect 3144 5195 3196 5255
rect 3234 5455 3286 5515
rect 3544 5455 3596 5515
rect 3634 5455 3686 5515
rect 3944 5455 3996 5515
rect 4034 5455 4086 5515
rect 4344 5455 4396 5515
rect 4434 5455 4486 5515
rect 4744 5455 4796 5515
rect 4834 5455 4886 5515
rect 5144 5455 5196 5515
rect 5234 5455 5286 5515
rect 5544 5455 5596 5515
rect 5634 5455 5686 5515
rect 5944 5455 5996 5515
rect 6034 5455 6086 5515
rect 6344 5455 6396 5515
rect 6434 5455 6486 5515
rect 6744 5455 6796 5515
rect 6834 5455 6886 5515
rect 7144 5455 7196 5515
rect 7234 5455 7286 5515
rect 7544 5455 7596 5515
rect 7634 5455 7686 5515
rect 7944 5455 7996 5515
rect 8034 5455 8086 5515
rect 8344 5455 8396 5515
rect 8434 5455 8486 5515
rect 8744 5455 8796 5515
rect 8834 5455 8886 5515
rect 9144 5455 9196 5515
rect 9234 5455 9286 5515
rect 9544 5455 9596 5515
rect 9634 5455 9686 5515
rect 9944 5455 9996 5515
rect 10034 5455 10086 5515
rect 10344 5455 10396 5515
rect 10434 5455 10486 5515
rect 10744 5455 10796 5515
rect 10834 5455 10886 5515
rect 11144 5455 11196 5515
rect 11234 5455 11286 5515
rect 11544 5455 11596 5515
rect 11634 5455 11686 5515
rect 11944 5455 11996 5515
rect 12034 5455 12086 5515
rect 12344 5455 12396 5515
rect 12434 5455 12486 5515
rect 12744 5455 12796 5515
rect 12834 5455 12886 5515
rect 13144 5455 13196 5515
rect 3234 5195 3286 5255
rect 3544 5195 3596 5255
rect 3634 5195 3686 5255
rect 3944 5195 3996 5255
rect 4034 5195 4086 5255
rect 4344 5195 4396 5255
rect 4434 5195 4486 5255
rect 4744 5195 4796 5255
rect 4834 5195 4886 5255
rect 5144 5195 5196 5255
rect 5234 5195 5286 5255
rect 5544 5195 5596 5255
rect 5634 5195 5686 5255
rect 5944 5195 5996 5255
rect 6034 5195 6086 5255
rect 6344 5195 6396 5255
rect 6434 5195 6486 5255
rect 6744 5195 6796 5255
rect 6834 5195 6886 5255
rect 7144 5195 7196 5255
rect 7234 5195 7286 5255
rect 7544 5195 7596 5255
rect 7634 5195 7686 5255
rect 7944 5195 7996 5255
rect 8034 5195 8086 5255
rect 8344 5195 8396 5255
rect 8434 5195 8486 5255
rect 8744 5195 8796 5255
rect 8834 5195 8886 5255
rect 9144 5195 9196 5255
rect 9234 5195 9286 5255
rect 9544 5195 9596 5255
rect 9634 5195 9686 5255
rect 9944 5195 9996 5255
rect 10034 5195 10086 5255
rect 10344 5195 10396 5255
rect 10434 5195 10486 5255
rect 10744 5195 10796 5255
rect 10834 5195 10886 5255
rect 11144 5195 11196 5255
rect 11234 5195 11286 5255
rect 11544 5195 11596 5255
rect 11634 5195 11686 5255
rect 11944 5195 11996 5255
rect 12034 5195 12086 5255
rect 12344 5195 12396 5255
rect 12434 5195 12486 5255
rect 12744 5195 12796 5255
rect 12834 5195 12886 5255
rect 13144 5195 13196 5255
rect -366 5085 -330 5145
rect -330 5085 -314 5145
rect -56 5085 -4 5145
rect -366 4825 -330 4885
rect -330 4825 -314 4885
rect -56 4825 -4 4885
rect 34 5085 86 5145
rect 344 5085 396 5145
rect 434 5085 486 5145
rect 744 5085 796 5145
rect 834 5085 886 5145
rect 1144 5085 1196 5145
rect 1234 5085 1286 5145
rect 1544 5085 1596 5145
rect 1634 5085 1686 5145
rect 1944 5085 1996 5145
rect 2034 5085 2086 5145
rect 2344 5085 2396 5145
rect 2434 5085 2486 5145
rect 2744 5085 2796 5145
rect 2834 5085 2886 5145
rect 3144 5085 3196 5145
rect 34 4825 86 4885
rect 344 4825 396 4885
rect 434 4825 486 4885
rect 744 4825 796 4885
rect 834 4825 886 4885
rect 1144 4825 1196 4885
rect 1234 4825 1286 4885
rect 1544 4825 1596 4885
rect 1634 4825 1686 4885
rect 1944 4825 1996 4885
rect 2034 4825 2086 4885
rect 2344 4825 2396 4885
rect 2434 4825 2486 4885
rect 2744 4825 2796 4885
rect 2834 4825 2886 4885
rect 3144 4825 3196 4885
rect 3234 5085 3286 5145
rect 3544 5085 3596 5145
rect 3634 5085 3686 5145
rect 3944 5085 3996 5145
rect 4034 5085 4086 5145
rect 4344 5085 4396 5145
rect 4434 5085 4486 5145
rect 4744 5085 4796 5145
rect 4834 5085 4886 5145
rect 5144 5085 5196 5145
rect 5234 5085 5286 5145
rect 5544 5085 5596 5145
rect 5634 5085 5686 5145
rect 5944 5085 5996 5145
rect 6034 5085 6086 5145
rect 6344 5085 6396 5145
rect 6434 5085 6486 5145
rect 6744 5085 6796 5145
rect 6834 5085 6886 5145
rect 7144 5085 7196 5145
rect 7234 5085 7286 5145
rect 7544 5085 7596 5145
rect 7634 5085 7686 5145
rect 7944 5085 7996 5145
rect 8034 5085 8086 5145
rect 8344 5085 8396 5145
rect 8434 5085 8486 5145
rect 8744 5085 8796 5145
rect 8834 5085 8886 5145
rect 9144 5085 9196 5145
rect 9234 5085 9286 5145
rect 9544 5085 9596 5145
rect 9634 5085 9686 5145
rect 9944 5085 9996 5145
rect 10034 5085 10086 5145
rect 10344 5085 10396 5145
rect 10434 5085 10486 5145
rect 10744 5085 10796 5145
rect 10834 5085 10886 5145
rect 11144 5085 11196 5145
rect 11234 5085 11286 5145
rect 11544 5085 11596 5145
rect 11634 5085 11686 5145
rect 11944 5085 11996 5145
rect 12034 5085 12086 5145
rect 12344 5085 12396 5145
rect 12434 5085 12486 5145
rect 12744 5085 12796 5145
rect 12834 5085 12886 5145
rect 13144 5085 13196 5145
rect 3234 4825 3286 4885
rect 3544 4825 3596 4885
rect 3634 4825 3686 4885
rect 3944 4825 3996 4885
rect 4034 4825 4086 4885
rect 4344 4825 4396 4885
rect 4434 4825 4486 4885
rect 4744 4825 4796 4885
rect 4834 4825 4886 4885
rect 5144 4825 5196 4885
rect 5234 4825 5286 4885
rect 5544 4825 5596 4885
rect 5634 4825 5686 4885
rect 5944 4825 5996 4885
rect 6034 4825 6086 4885
rect 6344 4825 6396 4885
rect 6434 4825 6486 4885
rect 6744 4825 6796 4885
rect 6834 4825 6886 4885
rect 7144 4825 7196 4885
rect 7234 4825 7286 4885
rect 7544 4825 7596 4885
rect 7634 4825 7686 4885
rect 7944 4825 7996 4885
rect 8034 4825 8086 4885
rect 8344 4825 8396 4885
rect 8434 4825 8486 4885
rect 8744 4825 8796 4885
rect 8834 4825 8886 4885
rect 9144 4825 9196 4885
rect 9234 4825 9286 4885
rect 9544 4825 9596 4885
rect 9634 4825 9686 4885
rect 9944 4825 9996 4885
rect 10034 4825 10086 4885
rect 10344 4825 10396 4885
rect 10434 4825 10486 4885
rect 10744 4825 10796 4885
rect 10834 4825 10886 4885
rect 11144 4825 11196 4885
rect 11234 4825 11286 4885
rect 11544 4825 11596 4885
rect 11634 4825 11686 4885
rect 11944 4825 11996 4885
rect 12034 4825 12086 4885
rect 12344 4825 12396 4885
rect 12434 4825 12486 4885
rect 12744 4825 12796 4885
rect 12834 4825 12886 4885
rect 13144 4825 13196 4885
rect -366 4715 -330 4775
rect -330 4715 -314 4775
rect -56 4715 -4 4775
rect -366 4455 -330 4515
rect -330 4455 -314 4515
rect -56 4455 -4 4515
rect 34 4715 86 4775
rect 344 4715 396 4775
rect 434 4715 486 4775
rect 744 4715 796 4775
rect 834 4715 886 4775
rect 1144 4715 1196 4775
rect 1234 4715 1286 4775
rect 1544 4715 1596 4775
rect 1634 4715 1686 4775
rect 1944 4715 1996 4775
rect 2034 4715 2086 4775
rect 2344 4715 2396 4775
rect 2434 4715 2486 4775
rect 2744 4715 2796 4775
rect 2834 4715 2886 4775
rect 3144 4715 3196 4775
rect 34 4455 86 4515
rect 344 4455 396 4515
rect 434 4455 486 4515
rect 744 4455 796 4515
rect 834 4455 886 4515
rect 1144 4455 1196 4515
rect 1234 4455 1286 4515
rect 1544 4455 1596 4515
rect 1634 4455 1686 4515
rect 1944 4455 1996 4515
rect 2034 4455 2086 4515
rect 2344 4455 2396 4515
rect 2434 4455 2486 4515
rect 2744 4455 2796 4515
rect 2834 4455 2886 4515
rect 3144 4455 3196 4515
rect 3234 4715 3286 4775
rect 3544 4715 3596 4775
rect 3634 4715 3686 4775
rect 3944 4715 3996 4775
rect 4034 4715 4086 4775
rect 4344 4715 4396 4775
rect 4434 4715 4486 4775
rect 4744 4715 4796 4775
rect 4834 4715 4886 4775
rect 5144 4715 5196 4775
rect 5234 4715 5286 4775
rect 5544 4715 5596 4775
rect 5634 4715 5686 4775
rect 5944 4715 5996 4775
rect 6034 4715 6086 4775
rect 6344 4715 6396 4775
rect 6434 4715 6486 4775
rect 6744 4715 6796 4775
rect 6834 4715 6886 4775
rect 7144 4715 7196 4775
rect 7234 4715 7286 4775
rect 7544 4715 7596 4775
rect 7634 4715 7686 4775
rect 7944 4715 7996 4775
rect 8034 4715 8086 4775
rect 8344 4715 8396 4775
rect 8434 4715 8486 4775
rect 8744 4715 8796 4775
rect 8834 4715 8886 4775
rect 9144 4715 9196 4775
rect 9234 4715 9286 4775
rect 9544 4715 9596 4775
rect 9634 4715 9686 4775
rect 9944 4715 9996 4775
rect 10034 4715 10086 4775
rect 10344 4715 10396 4775
rect 10434 4715 10486 4775
rect 10744 4715 10796 4775
rect 10834 4715 10886 4775
rect 11144 4715 11196 4775
rect 11234 4715 11286 4775
rect 11544 4715 11596 4775
rect 11634 4715 11686 4775
rect 11944 4715 11996 4775
rect 12034 4715 12086 4775
rect 12344 4715 12396 4775
rect 12434 4715 12486 4775
rect 12744 4715 12796 4775
rect 12834 4715 12886 4775
rect 13144 4715 13196 4775
rect 3234 4455 3286 4515
rect 3544 4455 3596 4515
rect 3634 4455 3686 4515
rect 3944 4455 3996 4515
rect 4034 4455 4086 4515
rect 4344 4455 4396 4515
rect 4434 4455 4486 4515
rect 4744 4455 4796 4515
rect 4834 4455 4886 4515
rect 5144 4455 5196 4515
rect 5234 4455 5286 4515
rect 5544 4455 5596 4515
rect 5634 4455 5686 4515
rect 5944 4455 5996 4515
rect 6034 4455 6086 4515
rect 6344 4455 6396 4515
rect 6434 4455 6486 4515
rect 6744 4455 6796 4515
rect 6834 4455 6886 4515
rect 7144 4455 7196 4515
rect 7234 4455 7286 4515
rect 7544 4455 7596 4515
rect 7634 4455 7686 4515
rect 7944 4455 7996 4515
rect 8034 4455 8086 4515
rect 8344 4455 8396 4515
rect 8434 4455 8486 4515
rect 8744 4455 8796 4515
rect 8834 4455 8886 4515
rect 9144 4455 9196 4515
rect 9234 4455 9286 4515
rect 9544 4455 9596 4515
rect 9634 4455 9686 4515
rect 9944 4455 9996 4515
rect 10034 4455 10086 4515
rect 10344 4455 10396 4515
rect 10434 4455 10486 4515
rect 10744 4455 10796 4515
rect 10834 4455 10886 4515
rect 11144 4455 11196 4515
rect 11234 4455 11286 4515
rect 11544 4455 11596 4515
rect 11634 4455 11686 4515
rect 11944 4455 11996 4515
rect 12034 4455 12086 4515
rect 12344 4455 12396 4515
rect 12434 4455 12486 4515
rect 12744 4455 12796 4515
rect 12834 4455 12886 4515
rect 13144 4455 13196 4515
rect -366 4345 -330 4405
rect -330 4345 -314 4405
rect -56 4345 -4 4405
rect -366 4085 -330 4145
rect -330 4085 -314 4145
rect -56 4085 -4 4145
rect 34 4345 86 4405
rect 344 4345 396 4405
rect 434 4345 486 4405
rect 744 4345 796 4405
rect 834 4345 886 4405
rect 1144 4345 1196 4405
rect 1234 4345 1286 4405
rect 1544 4345 1596 4405
rect 1634 4345 1686 4405
rect 1944 4345 1996 4405
rect 2034 4345 2086 4405
rect 2344 4345 2396 4405
rect 2434 4345 2486 4405
rect 2744 4345 2796 4405
rect 2834 4345 2886 4405
rect 3144 4345 3196 4405
rect 34 4085 86 4145
rect 344 4085 396 4145
rect 434 4085 486 4145
rect 744 4085 796 4145
rect 834 4085 886 4145
rect 1144 4085 1196 4145
rect 1234 4085 1286 4145
rect 1544 4085 1596 4145
rect 1634 4085 1686 4145
rect 1944 4085 1996 4145
rect 2034 4085 2086 4145
rect 2344 4085 2396 4145
rect 2434 4085 2486 4145
rect 2744 4085 2796 4145
rect 2834 4085 2886 4145
rect 3144 4085 3196 4145
rect 3234 4345 3286 4405
rect 3544 4345 3596 4405
rect 3634 4345 3686 4405
rect 3944 4345 3996 4405
rect 4034 4345 4086 4405
rect 4344 4345 4396 4405
rect 4434 4345 4486 4405
rect 4744 4345 4796 4405
rect 4834 4345 4886 4405
rect 5144 4345 5196 4405
rect 5234 4345 5286 4405
rect 5544 4345 5596 4405
rect 5634 4345 5686 4405
rect 5944 4345 5996 4405
rect 6034 4345 6086 4405
rect 6344 4345 6396 4405
rect 6434 4345 6486 4405
rect 6744 4345 6796 4405
rect 6834 4345 6886 4405
rect 7144 4345 7196 4405
rect 7234 4345 7286 4405
rect 7544 4345 7596 4405
rect 7634 4345 7686 4405
rect 7944 4345 7996 4405
rect 8034 4345 8086 4405
rect 8344 4345 8396 4405
rect 8434 4345 8486 4405
rect 8744 4345 8796 4405
rect 8834 4345 8886 4405
rect 9144 4345 9196 4405
rect 9234 4345 9286 4405
rect 9544 4345 9596 4405
rect 9634 4345 9686 4405
rect 9944 4345 9996 4405
rect 10034 4345 10086 4405
rect 10344 4345 10396 4405
rect 10434 4345 10486 4405
rect 10744 4345 10796 4405
rect 10834 4345 10886 4405
rect 11144 4345 11196 4405
rect 11234 4345 11286 4405
rect 11544 4345 11596 4405
rect 11634 4345 11686 4405
rect 11944 4345 11996 4405
rect 12034 4345 12086 4405
rect 12344 4345 12396 4405
rect 12434 4345 12486 4405
rect 12744 4345 12796 4405
rect 12834 4345 12886 4405
rect 13144 4345 13196 4405
rect 3234 4085 3286 4145
rect 3544 4085 3596 4145
rect 3634 4085 3686 4145
rect 3944 4085 3996 4145
rect 4034 4085 4086 4145
rect 4344 4085 4396 4145
rect 4434 4085 4486 4145
rect 4744 4085 4796 4145
rect 4834 4085 4886 4145
rect 5144 4085 5196 4145
rect 5234 4085 5286 4145
rect 5544 4085 5596 4145
rect 5634 4085 5686 4145
rect 5944 4085 5996 4145
rect 6034 4085 6086 4145
rect 6344 4085 6396 4145
rect 6434 4085 6486 4145
rect 6744 4085 6796 4145
rect 6834 4085 6886 4145
rect 7144 4085 7196 4145
rect 7234 4085 7286 4145
rect 7544 4085 7596 4145
rect 7634 4085 7686 4145
rect 7944 4085 7996 4145
rect 8034 4085 8086 4145
rect 8344 4085 8396 4145
rect 8434 4085 8486 4145
rect 8744 4085 8796 4145
rect 8834 4085 8886 4145
rect 9144 4085 9196 4145
rect 9234 4085 9286 4145
rect 9544 4085 9596 4145
rect 9634 4085 9686 4145
rect 9944 4085 9996 4145
rect 10034 4085 10086 4145
rect 10344 4085 10396 4145
rect 10434 4085 10486 4145
rect 10744 4085 10796 4145
rect 10834 4085 10886 4145
rect 11144 4085 11196 4145
rect 11234 4085 11286 4145
rect 11544 4085 11596 4145
rect 11634 4085 11686 4145
rect 11944 4085 11996 4145
rect 12034 4085 12086 4145
rect 12344 4085 12396 4145
rect 12434 4085 12486 4145
rect 12744 4085 12796 4145
rect 12834 4085 12886 4145
rect 13144 4085 13196 4145
rect -366 3975 -330 4035
rect -330 3975 -314 4035
rect -56 3975 -4 4035
rect -366 3715 -330 3775
rect -330 3715 -314 3775
rect -56 3715 -4 3775
rect 34 3975 86 4035
rect 344 3975 396 4035
rect 434 3975 486 4035
rect 744 3975 796 4035
rect 834 3975 886 4035
rect 1144 3975 1196 4035
rect 1234 3975 1286 4035
rect 1544 3975 1596 4035
rect 1634 3975 1686 4035
rect 1944 3975 1996 4035
rect 2034 3975 2086 4035
rect 2344 3975 2396 4035
rect 2434 3975 2486 4035
rect 2744 3975 2796 4035
rect 2834 3975 2886 4035
rect 3144 3975 3196 4035
rect 3234 3975 3286 4035
rect 3544 3975 3596 4035
rect 3634 3975 3686 4035
rect 3944 3975 3996 4035
rect 4034 3975 4086 4035
rect 4344 3975 4396 4035
rect 4434 3975 4486 4035
rect 4744 3975 4796 4035
rect 4834 3975 4886 4035
rect 5144 3975 5196 4035
rect 5234 3975 5286 4035
rect 5544 3975 5596 4035
rect 5634 3975 5686 4035
rect 5944 3975 5996 4035
rect 6034 3975 6086 4035
rect 6344 3975 6396 4035
rect 6434 3975 6486 4035
rect 6744 3975 6796 4035
rect 6834 3975 6886 4035
rect 7144 3975 7196 4035
rect 7234 3975 7286 4035
rect 7544 3975 7596 4035
rect 7634 3975 7686 4035
rect 7944 3975 7996 4035
rect 8034 3975 8086 4035
rect 8344 3975 8396 4035
rect 8434 3975 8486 4035
rect 8744 3975 8796 4035
rect 8834 3975 8886 4035
rect 9144 3975 9196 4035
rect 9234 3975 9286 4035
rect 9544 3975 9596 4035
rect 9634 3975 9686 4035
rect 9944 3975 9996 4035
rect 10034 3975 10086 4035
rect 10344 3975 10396 4035
rect 10434 3975 10486 4035
rect 10744 3975 10796 4035
rect 10834 3975 10886 4035
rect 11144 3975 11196 4035
rect 11234 3975 11286 4035
rect 11544 3975 11596 4035
rect 11634 3975 11686 4035
rect 11944 3975 11996 4035
rect 12034 3975 12086 4035
rect 12344 3975 12396 4035
rect 12434 3975 12486 4035
rect 12744 3975 12796 4035
rect 12834 3975 12886 4035
rect 13144 3975 13196 4035
rect 34 3715 86 3775
rect 344 3715 396 3775
rect 434 3715 486 3775
rect 744 3715 796 3775
rect 834 3715 886 3775
rect 1144 3715 1196 3775
rect 1234 3715 1286 3775
rect 1544 3715 1596 3775
rect 1634 3715 1686 3775
rect 1944 3715 1996 3775
rect 2034 3715 2086 3775
rect 2344 3715 2396 3775
rect 2434 3715 2486 3775
rect 2744 3715 2796 3775
rect 2834 3715 2886 3775
rect 3144 3715 3196 3775
rect 3234 3715 3286 3775
rect 3544 3715 3596 3775
rect 3634 3715 3686 3775
rect 3944 3715 3996 3775
rect 4034 3715 4086 3775
rect 4344 3715 4396 3775
rect 4434 3715 4486 3775
rect 4744 3715 4796 3775
rect 4834 3715 4886 3775
rect 5144 3715 5196 3775
rect 5234 3715 5286 3775
rect 5544 3715 5596 3775
rect 5634 3715 5686 3775
rect 5944 3715 5996 3775
rect 6034 3715 6086 3775
rect 6344 3715 6396 3775
rect 6434 3715 6486 3775
rect 6744 3715 6796 3775
rect 6834 3715 6886 3775
rect 7144 3715 7196 3775
rect 7234 3715 7286 3775
rect 7544 3715 7596 3775
rect 7634 3715 7686 3775
rect 7944 3715 7996 3775
rect 8034 3715 8086 3775
rect 8344 3715 8396 3775
rect 8434 3715 8486 3775
rect 8744 3715 8796 3775
rect 8834 3715 8886 3775
rect 9144 3715 9196 3775
rect 9234 3715 9286 3775
rect 9544 3715 9596 3775
rect 9634 3715 9686 3775
rect 9944 3715 9996 3775
rect 10034 3715 10086 3775
rect 10344 3715 10396 3775
rect 10434 3715 10486 3775
rect 10744 3715 10796 3775
rect 10834 3715 10886 3775
rect 11144 3715 11196 3775
rect 11234 3715 11286 3775
rect 11544 3715 11596 3775
rect 11634 3715 11686 3775
rect 11944 3715 11996 3775
rect 12034 3715 12086 3775
rect 12344 3715 12396 3775
rect 12434 3715 12486 3775
rect 12744 3715 12796 3775
rect 12834 3715 12886 3775
rect 13144 3715 13196 3775
rect -366 3605 -330 3665
rect -330 3605 -314 3665
rect -56 3605 -4 3665
rect -366 3345 -330 3405
rect -330 3345 -314 3405
rect -56 3345 -4 3405
rect 34 3605 86 3665
rect 344 3605 396 3665
rect 434 3605 486 3665
rect 744 3605 796 3665
rect 834 3605 886 3665
rect 1144 3605 1196 3665
rect 1234 3605 1286 3665
rect 1544 3605 1596 3665
rect 1634 3605 1686 3665
rect 1944 3605 1996 3665
rect 2034 3605 2086 3665
rect 2344 3605 2396 3665
rect 2434 3605 2486 3665
rect 2744 3605 2796 3665
rect 2834 3605 2886 3665
rect 3144 3605 3196 3665
rect 3234 3605 3286 3665
rect 3544 3605 3596 3665
rect 3634 3605 3686 3665
rect 3944 3605 3996 3665
rect 4034 3605 4086 3665
rect 4344 3605 4396 3665
rect 4434 3605 4486 3665
rect 4744 3605 4796 3665
rect 4834 3605 4886 3665
rect 5144 3605 5196 3665
rect 5234 3605 5286 3665
rect 5544 3605 5596 3665
rect 5634 3605 5686 3665
rect 5944 3605 5996 3665
rect 6034 3605 6086 3665
rect 6344 3605 6396 3665
rect 6434 3605 6486 3665
rect 6744 3605 6796 3665
rect 6834 3605 6886 3665
rect 7144 3605 7196 3665
rect 7234 3605 7286 3665
rect 7544 3605 7596 3665
rect 7634 3605 7686 3665
rect 7944 3605 7996 3665
rect 8034 3605 8086 3665
rect 8344 3605 8396 3665
rect 8434 3605 8486 3665
rect 8744 3605 8796 3665
rect 8834 3605 8886 3665
rect 9144 3605 9196 3665
rect 9234 3605 9286 3665
rect 9544 3605 9596 3665
rect 9634 3605 9686 3665
rect 9944 3605 9996 3665
rect 10034 3605 10086 3665
rect 10344 3605 10396 3665
rect 10434 3605 10486 3665
rect 10744 3605 10796 3665
rect 10834 3605 10886 3665
rect 11144 3605 11196 3665
rect 11234 3605 11286 3665
rect 11544 3605 11596 3665
rect 11634 3605 11686 3665
rect 11944 3605 11996 3665
rect 12034 3605 12086 3665
rect 12344 3605 12396 3665
rect 12434 3605 12486 3665
rect 12744 3605 12796 3665
rect 12834 3605 12886 3665
rect 13144 3605 13196 3665
rect 34 3345 86 3405
rect 344 3345 396 3405
rect 434 3345 486 3405
rect 744 3345 796 3405
rect 834 3345 886 3405
rect 1144 3345 1196 3405
rect 1234 3345 1286 3405
rect 1544 3345 1596 3405
rect 1634 3345 1686 3405
rect 1944 3345 1996 3405
rect 2034 3345 2086 3405
rect 2344 3345 2396 3405
rect 2434 3345 2486 3405
rect 2744 3345 2796 3405
rect 2834 3345 2886 3405
rect 3144 3345 3196 3405
rect 3234 3345 3286 3405
rect 3544 3345 3596 3405
rect 3634 3345 3686 3405
rect 3944 3345 3996 3405
rect 4034 3345 4086 3405
rect 4344 3345 4396 3405
rect 4434 3345 4486 3405
rect 4744 3345 4796 3405
rect 4834 3345 4886 3405
rect 5144 3345 5196 3405
rect 5234 3345 5286 3405
rect 5544 3345 5596 3405
rect 5634 3345 5686 3405
rect 5944 3345 5996 3405
rect 6034 3345 6086 3405
rect 6344 3345 6396 3405
rect 6434 3345 6486 3405
rect 6744 3345 6796 3405
rect 6834 3345 6886 3405
rect 7144 3345 7196 3405
rect 7234 3345 7286 3405
rect 7544 3345 7596 3405
rect 7634 3345 7686 3405
rect 7944 3345 7996 3405
rect 8034 3345 8086 3405
rect 8344 3345 8396 3405
rect 8434 3345 8486 3405
rect 8744 3345 8796 3405
rect 8834 3345 8886 3405
rect 9144 3345 9196 3405
rect 9234 3345 9286 3405
rect 9544 3345 9596 3405
rect 9634 3345 9686 3405
rect 9944 3345 9996 3405
rect 10034 3345 10086 3405
rect 10344 3345 10396 3405
rect 10434 3345 10486 3405
rect 10744 3345 10796 3405
rect 10834 3345 10886 3405
rect 11144 3345 11196 3405
rect 11234 3345 11286 3405
rect 11544 3345 11596 3405
rect 11634 3345 11686 3405
rect 11944 3345 11996 3405
rect 12034 3345 12086 3405
rect 12344 3345 12396 3405
rect 12434 3345 12486 3405
rect 12744 3345 12796 3405
rect 12834 3345 12886 3405
rect 13144 3345 13196 3405
rect -366 3235 -330 3295
rect -330 3235 -314 3295
rect -56 3235 -4 3295
rect -366 2975 -330 3035
rect -330 2975 -314 3035
rect -56 2975 -4 3035
rect 34 3235 86 3295
rect 344 3235 396 3295
rect 434 3235 486 3295
rect 744 3235 796 3295
rect 834 3235 886 3295
rect 1144 3235 1196 3295
rect 1234 3235 1286 3295
rect 1544 3235 1596 3295
rect 1634 3235 1686 3295
rect 1944 3235 1996 3295
rect 2034 3235 2086 3295
rect 2344 3235 2396 3295
rect 2434 3235 2486 3295
rect 2744 3235 2796 3295
rect 2834 3235 2886 3295
rect 3144 3235 3196 3295
rect 3234 3235 3286 3295
rect 3544 3235 3596 3295
rect 3634 3235 3686 3295
rect 3944 3235 3996 3295
rect 4034 3235 4086 3295
rect 4344 3235 4396 3295
rect 4434 3235 4486 3295
rect 4744 3235 4796 3295
rect 4834 3235 4886 3295
rect 5144 3235 5196 3295
rect 5234 3235 5286 3295
rect 5544 3235 5596 3295
rect 5634 3235 5686 3295
rect 5944 3235 5996 3295
rect 6034 3235 6086 3295
rect 6344 3235 6396 3295
rect 6434 3235 6486 3295
rect 6744 3235 6796 3295
rect 6834 3235 6886 3295
rect 7144 3235 7196 3295
rect 7234 3235 7286 3295
rect 7544 3235 7596 3295
rect 7634 3235 7686 3295
rect 7944 3235 7996 3295
rect 8034 3235 8086 3295
rect 8344 3235 8396 3295
rect 8434 3235 8486 3295
rect 8744 3235 8796 3295
rect 8834 3235 8886 3295
rect 9144 3235 9196 3295
rect 9234 3235 9286 3295
rect 9544 3235 9596 3295
rect 9634 3235 9686 3295
rect 9944 3235 9996 3295
rect 10034 3235 10086 3295
rect 10344 3235 10396 3295
rect 10434 3235 10486 3295
rect 10744 3235 10796 3295
rect 10834 3235 10886 3295
rect 11144 3235 11196 3295
rect 11234 3235 11286 3295
rect 11544 3235 11596 3295
rect 11634 3235 11686 3295
rect 11944 3235 11996 3295
rect 12034 3235 12086 3295
rect 12344 3235 12396 3295
rect 12434 3235 12486 3295
rect 12744 3235 12796 3295
rect 12834 3235 12886 3295
rect 13144 3235 13196 3295
rect 34 2975 86 3035
rect 344 2975 396 3035
rect 434 2975 486 3035
rect 744 2975 796 3035
rect 834 2975 886 3035
rect 1144 2975 1196 3035
rect 1234 2975 1286 3035
rect 1544 2975 1596 3035
rect 1634 2975 1686 3035
rect 1944 2975 1996 3035
rect 2034 2975 2086 3035
rect 2344 2975 2396 3035
rect 2434 2975 2486 3035
rect 2744 2975 2796 3035
rect 2834 2975 2886 3035
rect 3144 2975 3196 3035
rect 3234 2975 3286 3035
rect 3544 2975 3596 3035
rect 3634 2975 3686 3035
rect 3944 2975 3996 3035
rect 4034 2975 4086 3035
rect 4344 2975 4396 3035
rect 4434 2975 4486 3035
rect 4744 2975 4796 3035
rect 4834 2975 4886 3035
rect 5144 2975 5196 3035
rect 5234 2975 5286 3035
rect 5544 2975 5596 3035
rect 5634 2975 5686 3035
rect 5944 2975 5996 3035
rect 6034 2975 6086 3035
rect 6344 2975 6396 3035
rect 6434 2975 6486 3035
rect 6744 2975 6796 3035
rect 6834 2975 6886 3035
rect 7144 2975 7196 3035
rect 7234 2975 7286 3035
rect 7544 2975 7596 3035
rect 7634 2975 7686 3035
rect 7944 2975 7996 3035
rect 8034 2975 8086 3035
rect 8344 2975 8396 3035
rect 8434 2975 8486 3035
rect 8744 2975 8796 3035
rect 8834 2975 8886 3035
rect 9144 2975 9196 3035
rect 9234 2975 9286 3035
rect 9544 2975 9596 3035
rect 9634 2975 9686 3035
rect 9944 2975 9996 3035
rect 10034 2975 10086 3035
rect 10344 2975 10396 3035
rect 10434 2975 10486 3035
rect 10744 2975 10796 3035
rect 10834 2975 10886 3035
rect 11144 2975 11196 3035
rect 11234 2975 11286 3035
rect 11544 2975 11596 3035
rect 11634 2975 11686 3035
rect 11944 2975 11996 3035
rect 12034 2975 12086 3035
rect 12344 2975 12396 3035
rect 12434 2975 12486 3035
rect 12744 2975 12796 3035
rect 12834 2975 12886 3035
rect 13144 2975 13196 3035
rect -366 2865 -330 2925
rect -330 2865 -314 2925
rect -56 2865 -4 2925
rect -366 2605 -330 2665
rect -330 2605 -314 2665
rect -56 2605 -4 2665
rect 34 2865 86 2925
rect 344 2865 396 2925
rect 434 2865 486 2925
rect 744 2865 796 2925
rect 834 2865 886 2925
rect 1144 2865 1196 2925
rect 1234 2865 1286 2925
rect 1544 2865 1596 2925
rect 1634 2865 1686 2925
rect 1944 2865 1996 2925
rect 2034 2865 2086 2925
rect 2344 2865 2396 2925
rect 2434 2865 2486 2925
rect 2744 2865 2796 2925
rect 2834 2865 2886 2925
rect 3144 2865 3196 2925
rect 3234 2865 3286 2925
rect 3544 2865 3596 2925
rect 3634 2865 3686 2925
rect 3944 2865 3996 2925
rect 4034 2865 4086 2925
rect 4344 2865 4396 2925
rect 4434 2865 4486 2925
rect 4744 2865 4796 2925
rect 4834 2865 4886 2925
rect 5144 2865 5196 2925
rect 5234 2865 5286 2925
rect 5544 2865 5596 2925
rect 5634 2865 5686 2925
rect 5944 2865 5996 2925
rect 6034 2865 6086 2925
rect 6344 2865 6396 2925
rect 6434 2865 6486 2925
rect 6744 2865 6796 2925
rect 6834 2865 6886 2925
rect 7144 2865 7196 2925
rect 7234 2865 7286 2925
rect 7544 2865 7596 2925
rect 7634 2865 7686 2925
rect 7944 2865 7996 2925
rect 8034 2865 8086 2925
rect 8344 2865 8396 2925
rect 8434 2865 8486 2925
rect 8744 2865 8796 2925
rect 8834 2865 8886 2925
rect 9144 2865 9196 2925
rect 9234 2865 9286 2925
rect 9544 2865 9596 2925
rect 9634 2865 9686 2925
rect 9944 2865 9996 2925
rect 10034 2865 10086 2925
rect 10344 2865 10396 2925
rect 10434 2865 10486 2925
rect 10744 2865 10796 2925
rect 10834 2865 10886 2925
rect 11144 2865 11196 2925
rect 11234 2865 11286 2925
rect 11544 2865 11596 2925
rect 11634 2865 11686 2925
rect 11944 2865 11996 2925
rect 12034 2865 12086 2925
rect 12344 2865 12396 2925
rect 12434 2865 12486 2925
rect 12744 2865 12796 2925
rect 12834 2865 12886 2925
rect 13144 2865 13196 2925
rect 34 2605 86 2665
rect 344 2605 396 2665
rect 434 2605 486 2665
rect 744 2605 796 2665
rect 834 2605 886 2665
rect 1144 2605 1196 2665
rect 1234 2605 1286 2665
rect 1544 2605 1596 2665
rect 1634 2605 1686 2665
rect 1944 2605 1996 2665
rect 2034 2605 2086 2665
rect 2344 2605 2396 2665
rect 2434 2605 2486 2665
rect 2744 2605 2796 2665
rect 2834 2605 2886 2665
rect 3144 2605 3196 2665
rect 3234 2605 3286 2665
rect 3544 2605 3596 2665
rect 3634 2605 3686 2665
rect 3944 2605 3996 2665
rect 4034 2605 4086 2665
rect 4344 2605 4396 2665
rect 4434 2605 4486 2665
rect 4744 2605 4796 2665
rect 4834 2605 4886 2665
rect 5144 2605 5196 2665
rect 5234 2605 5286 2665
rect 5544 2605 5596 2665
rect 5634 2605 5686 2665
rect 5944 2605 5996 2665
rect 6034 2605 6086 2665
rect 6344 2605 6396 2665
rect 6434 2605 6486 2665
rect 6744 2605 6796 2665
rect 6834 2605 6886 2665
rect 7144 2605 7196 2665
rect 7234 2605 7286 2665
rect 7544 2605 7596 2665
rect 7634 2605 7686 2665
rect 7944 2605 7996 2665
rect 8034 2605 8086 2665
rect 8344 2605 8396 2665
rect 8434 2605 8486 2665
rect 8744 2605 8796 2665
rect 8834 2605 8886 2665
rect 9144 2605 9196 2665
rect 9234 2605 9286 2665
rect 9544 2605 9596 2665
rect 9634 2605 9686 2665
rect 9944 2605 9996 2665
rect 10034 2605 10086 2665
rect 10344 2605 10396 2665
rect 10434 2605 10486 2665
rect 10744 2605 10796 2665
rect 10834 2605 10886 2665
rect 11144 2605 11196 2665
rect 11234 2605 11286 2665
rect 11544 2605 11596 2665
rect 11634 2605 11686 2665
rect 11944 2605 11996 2665
rect 12034 2605 12086 2665
rect 12344 2605 12396 2665
rect 12434 2605 12486 2665
rect 12744 2605 12796 2665
rect 12834 2605 12886 2665
rect 13144 2605 13196 2665
rect -366 2495 -330 2555
rect -330 2495 -314 2555
rect -56 2495 -4 2555
rect -366 2235 -330 2295
rect -330 2235 -314 2295
rect -56 2235 -4 2295
rect 34 2495 86 2555
rect 344 2495 396 2555
rect 434 2495 486 2555
rect 744 2495 796 2555
rect 834 2495 886 2555
rect 1144 2495 1196 2555
rect 1234 2495 1286 2555
rect 1544 2495 1596 2555
rect 1634 2495 1686 2555
rect 1944 2495 1996 2555
rect 2034 2495 2086 2555
rect 2344 2495 2396 2555
rect 2434 2495 2486 2555
rect 2744 2495 2796 2555
rect 2834 2495 2886 2555
rect 3144 2495 3196 2555
rect 3234 2495 3286 2555
rect 3544 2495 3596 2555
rect 3634 2495 3686 2555
rect 3944 2495 3996 2555
rect 4034 2495 4086 2555
rect 4344 2495 4396 2555
rect 4434 2495 4486 2555
rect 4744 2495 4796 2555
rect 4834 2495 4886 2555
rect 5144 2495 5196 2555
rect 5234 2495 5286 2555
rect 5544 2495 5596 2555
rect 5634 2495 5686 2555
rect 5944 2495 5996 2555
rect 6034 2495 6086 2555
rect 6344 2495 6396 2555
rect 6434 2495 6486 2555
rect 6744 2495 6796 2555
rect 6834 2495 6886 2555
rect 7144 2495 7196 2555
rect 7234 2495 7286 2555
rect 7544 2495 7596 2555
rect 7634 2495 7686 2555
rect 7944 2495 7996 2555
rect 8034 2495 8086 2555
rect 8344 2495 8396 2555
rect 8434 2495 8486 2555
rect 8744 2495 8796 2555
rect 8834 2495 8886 2555
rect 9144 2495 9196 2555
rect 9234 2495 9286 2555
rect 9544 2495 9596 2555
rect 9634 2495 9686 2555
rect 9944 2495 9996 2555
rect 10034 2495 10086 2555
rect 10344 2495 10396 2555
rect 10434 2495 10486 2555
rect 10744 2495 10796 2555
rect 10834 2495 10886 2555
rect 11144 2495 11196 2555
rect 11234 2495 11286 2555
rect 11544 2495 11596 2555
rect 11634 2495 11686 2555
rect 11944 2495 11996 2555
rect 12034 2495 12086 2555
rect 12344 2495 12396 2555
rect 12434 2495 12486 2555
rect 12744 2495 12796 2555
rect 12834 2495 12886 2555
rect 13144 2495 13196 2555
rect 34 2235 86 2295
rect 344 2235 396 2295
rect 434 2235 486 2295
rect 744 2235 796 2295
rect 834 2235 886 2295
rect 1144 2235 1196 2295
rect 1234 2235 1286 2295
rect 1544 2235 1596 2295
rect 1634 2235 1686 2295
rect 1944 2235 1996 2295
rect 2034 2235 2086 2295
rect 2344 2235 2396 2295
rect 2434 2235 2486 2295
rect 2744 2235 2796 2295
rect 2834 2235 2886 2295
rect 3144 2235 3196 2295
rect 3234 2235 3286 2295
rect 3544 2235 3596 2295
rect 3634 2235 3686 2295
rect 3944 2235 3996 2295
rect 4034 2235 4086 2295
rect 4344 2235 4396 2295
rect 4434 2235 4486 2295
rect 4744 2235 4796 2295
rect 4834 2235 4886 2295
rect 5144 2235 5196 2295
rect 5234 2235 5286 2295
rect 5544 2235 5596 2295
rect 5634 2235 5686 2295
rect 5944 2235 5996 2295
rect 6034 2235 6086 2295
rect 6344 2235 6396 2295
rect 6434 2235 6486 2295
rect 6744 2235 6796 2295
rect 6834 2235 6886 2295
rect 7144 2235 7196 2295
rect 7234 2235 7286 2295
rect 7544 2235 7596 2295
rect 7634 2235 7686 2295
rect 7944 2235 7996 2295
rect 8034 2235 8086 2295
rect 8344 2235 8396 2295
rect 8434 2235 8486 2295
rect 8744 2235 8796 2295
rect 8834 2235 8886 2295
rect 9144 2235 9196 2295
rect 9234 2235 9286 2295
rect 9544 2235 9596 2295
rect 9634 2235 9686 2295
rect 9944 2235 9996 2295
rect 10034 2235 10086 2295
rect 10344 2235 10396 2295
rect 10434 2235 10486 2295
rect 10744 2235 10796 2295
rect 10834 2235 10886 2295
rect 11144 2235 11196 2295
rect 11234 2235 11286 2295
rect 11544 2235 11596 2295
rect 11634 2235 11686 2295
rect 11944 2235 11996 2295
rect 12034 2235 12086 2295
rect 12344 2235 12396 2295
rect 12434 2235 12486 2295
rect 12744 2235 12796 2295
rect 12834 2235 12886 2295
rect 13144 2235 13196 2295
rect -366 2125 -330 2185
rect -330 2125 -314 2185
rect -56 2125 -4 2185
rect -366 1865 -330 1925
rect -330 1865 -314 1925
rect -56 1865 -4 1925
rect 34 2125 86 2185
rect 344 2125 396 2185
rect 434 2125 486 2185
rect 744 2125 796 2185
rect 834 2125 886 2185
rect 1144 2125 1196 2185
rect 1234 2125 1286 2185
rect 1544 2125 1596 2185
rect 1634 2125 1686 2185
rect 1944 2125 1996 2185
rect 2034 2125 2086 2185
rect 2344 2125 2396 2185
rect 2434 2125 2486 2185
rect 2744 2125 2796 2185
rect 2834 2125 2886 2185
rect 3144 2125 3196 2185
rect 3234 2125 3286 2185
rect 3544 2125 3596 2185
rect 3634 2125 3686 2185
rect 3944 2125 3996 2185
rect 4034 2125 4086 2185
rect 4344 2125 4396 2185
rect 4434 2125 4486 2185
rect 4744 2125 4796 2185
rect 4834 2125 4886 2185
rect 5144 2125 5196 2185
rect 5234 2125 5286 2185
rect 5544 2125 5596 2185
rect 5634 2125 5686 2185
rect 5944 2125 5996 2185
rect 6034 2125 6086 2185
rect 6344 2125 6396 2185
rect 6434 2125 6486 2185
rect 6744 2125 6796 2185
rect 6834 2125 6886 2185
rect 7144 2125 7196 2185
rect 7234 2125 7286 2185
rect 7544 2125 7596 2185
rect 7634 2125 7686 2185
rect 7944 2125 7996 2185
rect 8034 2125 8086 2185
rect 8344 2125 8396 2185
rect 8434 2125 8486 2185
rect 8744 2125 8796 2185
rect 8834 2125 8886 2185
rect 9144 2125 9196 2185
rect 9234 2125 9286 2185
rect 9544 2125 9596 2185
rect 9634 2125 9686 2185
rect 9944 2125 9996 2185
rect 10034 2125 10086 2185
rect 10344 2125 10396 2185
rect 10434 2125 10486 2185
rect 10744 2125 10796 2185
rect 10834 2125 10886 2185
rect 11144 2125 11196 2185
rect 11234 2125 11286 2185
rect 11544 2125 11596 2185
rect 11634 2125 11686 2185
rect 11944 2125 11996 2185
rect 12034 2125 12086 2185
rect 12344 2125 12396 2185
rect 12434 2125 12486 2185
rect 12744 2125 12796 2185
rect 12834 2125 12886 2185
rect 13144 2125 13196 2185
rect 34 1865 86 1925
rect 344 1865 396 1925
rect 434 1865 486 1925
rect 744 1865 796 1925
rect 834 1865 886 1925
rect 1144 1865 1196 1925
rect 1234 1865 1286 1925
rect 1544 1865 1596 1925
rect 1634 1865 1686 1925
rect 1944 1865 1996 1925
rect 2034 1865 2086 1925
rect 2344 1865 2396 1925
rect 2434 1865 2486 1925
rect 2744 1865 2796 1925
rect 2834 1865 2886 1925
rect 3144 1865 3196 1925
rect 3234 1865 3286 1925
rect 3544 1865 3596 1925
rect 3634 1865 3686 1925
rect 3944 1865 3996 1925
rect 4034 1865 4086 1925
rect 4344 1865 4396 1925
rect 4434 1865 4486 1925
rect 4744 1865 4796 1925
rect 4834 1865 4886 1925
rect 5144 1865 5196 1925
rect 5234 1865 5286 1925
rect 5544 1865 5596 1925
rect 5634 1865 5686 1925
rect 5944 1865 5996 1925
rect 6034 1865 6086 1925
rect 6344 1865 6396 1925
rect 6434 1865 6486 1925
rect 6744 1865 6796 1925
rect 6834 1865 6886 1925
rect 7144 1865 7196 1925
rect 7234 1865 7286 1925
rect 7544 1865 7596 1925
rect 7634 1865 7686 1925
rect 7944 1865 7996 1925
rect 8034 1865 8086 1925
rect 8344 1865 8396 1925
rect 8434 1865 8486 1925
rect 8744 1865 8796 1925
rect 8834 1865 8886 1925
rect 9144 1865 9196 1925
rect 9234 1865 9286 1925
rect 9544 1865 9596 1925
rect 9634 1865 9686 1925
rect 9944 1865 9996 1925
rect 10034 1865 10086 1925
rect 10344 1865 10396 1925
rect 10434 1865 10486 1925
rect 10744 1865 10796 1925
rect 10834 1865 10886 1925
rect 11144 1865 11196 1925
rect 11234 1865 11286 1925
rect 11544 1865 11596 1925
rect 11634 1865 11686 1925
rect 11944 1865 11996 1925
rect 12034 1865 12086 1925
rect 12344 1865 12396 1925
rect 12434 1865 12486 1925
rect 12744 1865 12796 1925
rect 12834 1865 12886 1925
rect 13144 1865 13196 1925
rect -366 1755 -330 1815
rect -330 1755 -314 1815
rect -56 1755 -4 1815
rect -366 1495 -330 1555
rect -330 1495 -314 1555
rect -56 1495 -4 1555
rect 34 1755 86 1815
rect 344 1755 396 1815
rect 434 1755 486 1815
rect 744 1755 796 1815
rect 834 1755 886 1815
rect 1144 1755 1196 1815
rect 1234 1755 1286 1815
rect 1544 1755 1596 1815
rect 1634 1755 1686 1815
rect 1944 1755 1996 1815
rect 2034 1755 2086 1815
rect 2344 1755 2396 1815
rect 2434 1755 2486 1815
rect 2744 1755 2796 1815
rect 2834 1755 2886 1815
rect 3144 1755 3196 1815
rect 3234 1755 3286 1815
rect 3544 1755 3596 1815
rect 3634 1755 3686 1815
rect 3944 1755 3996 1815
rect 4034 1755 4086 1815
rect 4344 1755 4396 1815
rect 4434 1755 4486 1815
rect 4744 1755 4796 1815
rect 4834 1755 4886 1815
rect 5144 1755 5196 1815
rect 5234 1755 5286 1815
rect 5544 1755 5596 1815
rect 5634 1755 5686 1815
rect 5944 1755 5996 1815
rect 6034 1755 6086 1815
rect 6344 1755 6396 1815
rect 6434 1755 6486 1815
rect 6744 1755 6796 1815
rect 6834 1755 6886 1815
rect 7144 1755 7196 1815
rect 7234 1755 7286 1815
rect 7544 1755 7596 1815
rect 7634 1755 7686 1815
rect 7944 1755 7996 1815
rect 8034 1755 8086 1815
rect 8344 1755 8396 1815
rect 8434 1755 8486 1815
rect 8744 1755 8796 1815
rect 8834 1755 8886 1815
rect 9144 1755 9196 1815
rect 9234 1755 9286 1815
rect 9544 1755 9596 1815
rect 9634 1755 9686 1815
rect 9944 1755 9996 1815
rect 10034 1755 10086 1815
rect 10344 1755 10396 1815
rect 10434 1755 10486 1815
rect 10744 1755 10796 1815
rect 10834 1755 10886 1815
rect 11144 1755 11196 1815
rect 11234 1755 11286 1815
rect 11544 1755 11596 1815
rect 11634 1755 11686 1815
rect 11944 1755 11996 1815
rect 12034 1755 12086 1815
rect 12344 1755 12396 1815
rect 12434 1755 12486 1815
rect 12744 1755 12796 1815
rect 12834 1755 12886 1815
rect 13144 1755 13196 1815
rect 34 1495 86 1555
rect 344 1495 396 1555
rect 434 1495 486 1555
rect 744 1495 796 1555
rect 834 1495 886 1555
rect 1144 1495 1196 1555
rect 1234 1495 1286 1555
rect 1544 1495 1596 1555
rect 1634 1495 1686 1555
rect 1944 1495 1996 1555
rect 2034 1495 2086 1555
rect 2344 1495 2396 1555
rect 2434 1495 2486 1555
rect 2744 1495 2796 1555
rect 2834 1495 2886 1555
rect 3144 1495 3196 1555
rect 3234 1495 3286 1555
rect 3544 1495 3596 1555
rect 3634 1495 3686 1555
rect 3944 1495 3996 1555
rect 4034 1495 4086 1555
rect 4344 1495 4396 1555
rect 4434 1495 4486 1555
rect 4744 1495 4796 1555
rect 4834 1495 4886 1555
rect 5144 1495 5196 1555
rect 5234 1495 5286 1555
rect 5544 1495 5596 1555
rect 5634 1495 5686 1555
rect 5944 1495 5996 1555
rect 6034 1495 6086 1555
rect 6344 1495 6396 1555
rect 6434 1495 6486 1555
rect 6744 1495 6796 1555
rect 6834 1495 6886 1555
rect 7144 1495 7196 1555
rect 7234 1495 7286 1555
rect 7544 1495 7596 1555
rect 7634 1495 7686 1555
rect 7944 1495 7996 1555
rect 8034 1495 8086 1555
rect 8344 1495 8396 1555
rect 8434 1495 8486 1555
rect 8744 1495 8796 1555
rect 8834 1495 8886 1555
rect 9144 1495 9196 1555
rect 9234 1495 9286 1555
rect 9544 1495 9596 1555
rect 9634 1495 9686 1555
rect 9944 1495 9996 1555
rect 10034 1495 10086 1555
rect 10344 1495 10396 1555
rect 10434 1495 10486 1555
rect 10744 1495 10796 1555
rect 10834 1495 10886 1555
rect 11144 1495 11196 1555
rect 11234 1495 11286 1555
rect 11544 1495 11596 1555
rect 11634 1495 11686 1555
rect 11944 1495 11996 1555
rect 12034 1495 12086 1555
rect 12344 1495 12396 1555
rect 12434 1495 12486 1555
rect 12744 1495 12796 1555
rect 12834 1495 12886 1555
rect 13144 1495 13196 1555
rect -366 1385 -330 1445
rect -330 1385 -314 1445
rect -56 1385 -4 1445
rect -366 1125 -330 1185
rect -330 1125 -314 1185
rect -56 1125 -4 1185
rect 34 1385 86 1445
rect 344 1385 396 1445
rect 434 1385 486 1445
rect 744 1385 796 1445
rect 834 1385 886 1445
rect 1144 1385 1196 1445
rect 1234 1385 1286 1445
rect 1544 1385 1596 1445
rect 1634 1385 1686 1445
rect 1944 1385 1996 1445
rect 2034 1385 2086 1445
rect 2344 1385 2396 1445
rect 2434 1385 2486 1445
rect 2744 1385 2796 1445
rect 2834 1385 2886 1445
rect 3144 1385 3196 1445
rect 3234 1385 3286 1445
rect 3544 1385 3596 1445
rect 3634 1385 3686 1445
rect 3944 1385 3996 1445
rect 4034 1385 4086 1445
rect 4344 1385 4396 1445
rect 4434 1385 4486 1445
rect 4744 1385 4796 1445
rect 4834 1385 4886 1445
rect 5144 1385 5196 1445
rect 5234 1385 5286 1445
rect 5544 1385 5596 1445
rect 5634 1385 5686 1445
rect 5944 1385 5996 1445
rect 6034 1385 6086 1445
rect 6344 1385 6396 1445
rect 6434 1385 6486 1445
rect 6744 1385 6796 1445
rect 6834 1385 6886 1445
rect 7144 1385 7196 1445
rect 7234 1385 7286 1445
rect 7544 1385 7596 1445
rect 7634 1385 7686 1445
rect 7944 1385 7996 1445
rect 8034 1385 8086 1445
rect 8344 1385 8396 1445
rect 8434 1385 8486 1445
rect 8744 1385 8796 1445
rect 8834 1385 8886 1445
rect 9144 1385 9196 1445
rect 9234 1385 9286 1445
rect 9544 1385 9596 1445
rect 9634 1385 9686 1445
rect 9944 1385 9996 1445
rect 10034 1385 10086 1445
rect 10344 1385 10396 1445
rect 10434 1385 10486 1445
rect 10744 1385 10796 1445
rect 10834 1385 10886 1445
rect 11144 1385 11196 1445
rect 11234 1385 11286 1445
rect 11544 1385 11596 1445
rect 11634 1385 11686 1445
rect 11944 1385 11996 1445
rect 12034 1385 12086 1445
rect 12344 1385 12396 1445
rect 12434 1385 12486 1445
rect 12744 1385 12796 1445
rect 12834 1385 12886 1445
rect 13144 1385 13196 1445
rect 34 1125 86 1185
rect 344 1125 396 1185
rect 434 1125 486 1185
rect 744 1125 796 1185
rect 834 1125 886 1185
rect 1144 1125 1196 1185
rect 1234 1125 1286 1185
rect 1544 1125 1596 1185
rect 1634 1125 1686 1185
rect 1944 1125 1996 1185
rect 2034 1125 2086 1185
rect 2344 1125 2396 1185
rect 2434 1125 2486 1185
rect 2744 1125 2796 1185
rect 2834 1125 2886 1185
rect 3144 1125 3196 1185
rect 3234 1125 3286 1185
rect 3544 1125 3596 1185
rect 3634 1125 3686 1185
rect 3944 1125 3996 1185
rect 4034 1125 4086 1185
rect 4344 1125 4396 1185
rect 4434 1125 4486 1185
rect 4744 1125 4796 1185
rect 4834 1125 4886 1185
rect 5144 1125 5196 1185
rect 5234 1125 5286 1185
rect 5544 1125 5596 1185
rect 5634 1125 5686 1185
rect 5944 1125 5996 1185
rect 6034 1125 6086 1185
rect 6344 1125 6396 1185
rect 6434 1125 6486 1185
rect 6744 1125 6796 1185
rect 6834 1125 6886 1185
rect 7144 1125 7196 1185
rect 7234 1125 7286 1185
rect 7544 1125 7596 1185
rect 7634 1125 7686 1185
rect 7944 1125 7996 1185
rect 8034 1125 8086 1185
rect 8344 1125 8396 1185
rect 8434 1125 8486 1185
rect 8744 1125 8796 1185
rect 8834 1125 8886 1185
rect 9144 1125 9196 1185
rect 9234 1125 9286 1185
rect 9544 1125 9596 1185
rect 9634 1125 9686 1185
rect 9944 1125 9996 1185
rect 10034 1125 10086 1185
rect 10344 1125 10396 1185
rect 10434 1125 10486 1185
rect 10744 1125 10796 1185
rect 10834 1125 10886 1185
rect 11144 1125 11196 1185
rect 11234 1125 11286 1185
rect 11544 1125 11596 1185
rect 11634 1125 11686 1185
rect 11944 1125 11996 1185
rect 12034 1125 12086 1185
rect 12344 1125 12396 1185
rect 12434 1125 12486 1185
rect 12744 1125 12796 1185
rect 12834 1125 12886 1185
rect 13144 1125 13196 1185
rect -366 1015 -330 1075
rect -330 1015 -314 1075
rect -56 1015 -4 1075
rect -366 755 -330 815
rect -330 755 -314 815
rect -56 755 -4 815
rect 34 1015 86 1075
rect 344 1015 396 1075
rect 434 1015 486 1075
rect 744 1015 796 1075
rect 834 1015 886 1075
rect 1144 1015 1196 1075
rect 1234 1015 1286 1075
rect 1544 1015 1596 1075
rect 1634 1015 1686 1075
rect 1944 1015 1996 1075
rect 2034 1015 2086 1075
rect 2344 1015 2396 1075
rect 2434 1015 2486 1075
rect 2744 1015 2796 1075
rect 2834 1015 2886 1075
rect 3144 1015 3196 1075
rect 3234 1015 3286 1075
rect 3544 1015 3596 1075
rect 3634 1015 3686 1075
rect 3944 1015 3996 1075
rect 4034 1015 4086 1075
rect 4344 1015 4396 1075
rect 4434 1015 4486 1075
rect 4744 1015 4796 1075
rect 4834 1015 4886 1075
rect 5144 1015 5196 1075
rect 5234 1015 5286 1075
rect 5544 1015 5596 1075
rect 5634 1015 5686 1075
rect 5944 1015 5996 1075
rect 6034 1015 6086 1075
rect 6344 1015 6396 1075
rect 6434 1015 6486 1075
rect 6744 1015 6796 1075
rect 6834 1015 6886 1075
rect 7144 1015 7196 1075
rect 7234 1015 7286 1075
rect 7544 1015 7596 1075
rect 7634 1015 7686 1075
rect 7944 1015 7996 1075
rect 8034 1015 8086 1075
rect 8344 1015 8396 1075
rect 8434 1015 8486 1075
rect 8744 1015 8796 1075
rect 8834 1015 8886 1075
rect 9144 1015 9196 1075
rect 9234 1015 9286 1075
rect 9544 1015 9596 1075
rect 9634 1015 9686 1075
rect 9944 1015 9996 1075
rect 10034 1015 10086 1075
rect 10344 1015 10396 1075
rect 10434 1015 10486 1075
rect 10744 1015 10796 1075
rect 10834 1015 10886 1075
rect 11144 1015 11196 1075
rect 11234 1015 11286 1075
rect 11544 1015 11596 1075
rect 11634 1015 11686 1075
rect 11944 1015 11996 1075
rect 12034 1015 12086 1075
rect 12344 1015 12396 1075
rect 12434 1015 12486 1075
rect 12744 1015 12796 1075
rect 12834 1015 12886 1075
rect 13144 1015 13196 1075
rect 34 755 86 815
rect 344 755 396 815
rect 434 755 486 815
rect 744 755 796 815
rect 834 755 886 815
rect 1144 755 1196 815
rect 1234 755 1286 815
rect 1544 755 1596 815
rect 1634 755 1686 815
rect 1944 755 1996 815
rect 2034 755 2086 815
rect 2344 755 2396 815
rect 2434 755 2486 815
rect 2744 755 2796 815
rect 2834 755 2886 815
rect 3144 755 3196 815
rect 3234 755 3286 815
rect 3544 755 3596 815
rect 3634 755 3686 815
rect 3944 755 3996 815
rect 4034 755 4086 815
rect 4344 755 4396 815
rect 4434 755 4486 815
rect 4744 755 4796 815
rect 4834 755 4886 815
rect 5144 755 5196 815
rect 5234 755 5286 815
rect 5544 755 5596 815
rect 5634 755 5686 815
rect 5944 755 5996 815
rect 6034 755 6086 815
rect 6344 755 6396 815
rect 6434 755 6486 815
rect 6744 755 6796 815
rect 6834 755 6886 815
rect 7144 755 7196 815
rect 7234 755 7286 815
rect 7544 755 7596 815
rect 7634 755 7686 815
rect 7944 755 7996 815
rect 8034 755 8086 815
rect 8344 755 8396 815
rect 8434 755 8486 815
rect 8744 755 8796 815
rect 8834 755 8886 815
rect 9144 755 9196 815
rect 9234 755 9286 815
rect 9544 755 9596 815
rect 9634 755 9686 815
rect 9944 755 9996 815
rect 10034 755 10086 815
rect 10344 755 10396 815
rect 10434 755 10486 815
rect 10744 755 10796 815
rect 10834 755 10886 815
rect 11144 755 11196 815
rect 11234 755 11286 815
rect 11544 755 11596 815
rect 11634 755 11686 815
rect 11944 755 11996 815
rect 12034 755 12086 815
rect 12344 755 12396 815
rect 12434 755 12486 815
rect 12744 755 12796 815
rect 12834 755 12886 815
rect 13144 755 13196 815
rect -366 645 -330 705
rect -330 645 -314 705
rect -56 645 -4 705
rect -366 385 -330 445
rect -330 385 -314 445
rect -56 385 -4 445
rect 34 645 86 705
rect 344 645 396 705
rect 434 645 486 705
rect 744 645 796 705
rect 834 645 886 705
rect 1144 645 1196 705
rect 1234 645 1286 705
rect 1544 645 1596 705
rect 1634 645 1686 705
rect 1944 645 1996 705
rect 2034 645 2086 705
rect 2344 645 2396 705
rect 2434 645 2486 705
rect 2744 645 2796 705
rect 2834 645 2886 705
rect 3144 645 3196 705
rect 3234 645 3286 705
rect 3544 645 3596 705
rect 3634 645 3686 705
rect 3944 645 3996 705
rect 4034 645 4086 705
rect 4344 645 4396 705
rect 4434 645 4486 705
rect 4744 645 4796 705
rect 4834 645 4886 705
rect 5144 645 5196 705
rect 5234 645 5286 705
rect 5544 645 5596 705
rect 5634 645 5686 705
rect 5944 645 5996 705
rect 6034 645 6086 705
rect 6344 645 6396 705
rect 6434 645 6486 705
rect 6744 645 6796 705
rect 6834 645 6886 705
rect 7144 645 7196 705
rect 7234 645 7286 705
rect 7544 645 7596 705
rect 7634 645 7686 705
rect 7944 645 7996 705
rect 8034 645 8086 705
rect 8344 645 8396 705
rect 8434 645 8486 705
rect 8744 645 8796 705
rect 8834 645 8886 705
rect 9144 645 9196 705
rect 9234 645 9286 705
rect 9544 645 9596 705
rect 9634 645 9686 705
rect 9944 645 9996 705
rect 10034 645 10086 705
rect 10344 645 10396 705
rect 10434 645 10486 705
rect 10744 645 10796 705
rect 10834 645 10886 705
rect 11144 645 11196 705
rect 11234 645 11286 705
rect 11544 645 11596 705
rect 11634 645 11686 705
rect 11944 645 11996 705
rect 12034 645 12086 705
rect 12344 645 12396 705
rect 12434 645 12486 705
rect 12744 645 12796 705
rect 12834 645 12886 705
rect 13144 645 13196 705
rect 34 385 86 445
rect 344 385 396 445
rect 434 385 486 445
rect 744 385 796 445
rect 834 385 886 445
rect 1144 385 1196 445
rect 1234 385 1286 445
rect 1544 385 1596 445
rect 1634 385 1686 445
rect 1944 385 1996 445
rect 2034 385 2086 445
rect 2344 385 2396 445
rect 2434 385 2486 445
rect 2744 385 2796 445
rect 2834 385 2886 445
rect 3144 385 3196 445
rect 3234 385 3286 445
rect 3544 385 3596 445
rect 3634 385 3686 445
rect 3944 385 3996 445
rect 4034 385 4086 445
rect 4344 385 4396 445
rect 4434 385 4486 445
rect 4744 385 4796 445
rect 4834 385 4886 445
rect 5144 385 5196 445
rect 5234 385 5286 445
rect 5544 385 5596 445
rect 5634 385 5686 445
rect 5944 385 5996 445
rect 6034 385 6086 445
rect 6344 385 6396 445
rect 6434 385 6486 445
rect 6744 385 6796 445
rect 6834 385 6886 445
rect 7144 385 7196 445
rect 7234 385 7286 445
rect 7544 385 7596 445
rect 7634 385 7686 445
rect 7944 385 7996 445
rect 8034 385 8086 445
rect 8344 385 8396 445
rect 8434 385 8486 445
rect 8744 385 8796 445
rect 8834 385 8886 445
rect 9144 385 9196 445
rect 9234 385 9286 445
rect 9544 385 9596 445
rect 9634 385 9686 445
rect 9944 385 9996 445
rect 10034 385 10086 445
rect 10344 385 10396 445
rect 10434 385 10486 445
rect 10744 385 10796 445
rect 10834 385 10886 445
rect 11144 385 11196 445
rect 11234 385 11286 445
rect 11544 385 11596 445
rect 11634 385 11686 445
rect 11944 385 11996 445
rect 12034 385 12086 445
rect 12344 385 12396 445
rect 12434 385 12486 445
rect 12744 385 12796 445
rect 12834 385 12886 445
rect 13144 385 13196 445
rect -366 275 -330 335
rect -330 275 -314 335
rect -56 275 -4 335
rect -366 15 -330 75
rect -330 15 -314 75
rect -56 15 -4 75
rect 34 275 86 335
rect 344 275 396 335
rect 434 275 486 335
rect 744 275 796 335
rect 834 275 886 335
rect 1144 275 1196 335
rect 1234 275 1286 335
rect 1544 275 1596 335
rect 1634 275 1686 335
rect 1944 275 1996 335
rect 2034 275 2086 335
rect 2344 275 2396 335
rect 2434 275 2486 335
rect 2744 275 2796 335
rect 2834 275 2886 335
rect 3144 275 3196 335
rect 3234 275 3286 335
rect 3544 275 3596 335
rect 3634 275 3686 335
rect 3944 275 3996 335
rect 4034 275 4086 335
rect 4344 275 4396 335
rect 4434 275 4486 335
rect 4744 275 4796 335
rect 4834 275 4886 335
rect 5144 275 5196 335
rect 5234 275 5286 335
rect 5544 275 5596 335
rect 5634 275 5686 335
rect 5944 275 5996 335
rect 6034 275 6086 335
rect 6344 275 6396 335
rect 6434 275 6486 335
rect 6744 275 6796 335
rect 6834 275 6886 335
rect 7144 275 7196 335
rect 7234 275 7286 335
rect 7544 275 7596 335
rect 7634 275 7686 335
rect 7944 275 7996 335
rect 8034 275 8086 335
rect 8344 275 8396 335
rect 8434 275 8486 335
rect 8744 275 8796 335
rect 8834 275 8886 335
rect 9144 275 9196 335
rect 9234 275 9286 335
rect 9544 275 9596 335
rect 9634 275 9686 335
rect 9944 275 9996 335
rect 10034 275 10086 335
rect 10344 275 10396 335
rect 10434 275 10486 335
rect 10744 275 10796 335
rect 10834 275 10886 335
rect 11144 275 11196 335
rect 11234 275 11286 335
rect 11544 275 11596 335
rect 11634 275 11686 335
rect 11944 275 11996 335
rect 12034 275 12086 335
rect 12344 275 12396 335
rect 12434 275 12486 335
rect 12744 275 12796 335
rect 12834 275 12886 335
rect 13144 275 13196 335
rect 34 15 86 75
rect 344 15 396 75
rect 434 15 486 75
rect 744 15 796 75
rect 834 15 886 75
rect 1144 15 1196 75
rect 1234 15 1286 75
rect 1544 15 1596 75
rect 1634 15 1686 75
rect 1944 15 1996 75
rect 2034 15 2086 75
rect 2344 15 2396 75
rect 2434 15 2486 75
rect 2744 15 2796 75
rect 2834 15 2886 75
rect 3144 15 3196 75
rect 3234 15 3286 75
rect 3544 15 3596 75
rect 3634 15 3686 75
rect 3944 15 3996 75
rect 4034 15 4086 75
rect 4344 15 4396 75
rect 4434 15 4486 75
rect 4744 15 4796 75
rect 4834 15 4886 75
rect 5144 15 5196 75
rect 5234 15 5286 75
rect 5544 15 5596 75
rect 5634 15 5686 75
rect 5944 15 5996 75
rect 6034 15 6086 75
rect 6344 15 6396 75
rect 6434 15 6486 75
rect 6744 15 6796 75
rect 6834 15 6886 75
rect 7144 15 7196 75
rect 7234 15 7286 75
rect 7544 15 7596 75
rect 7634 15 7686 75
rect 7944 15 7996 75
rect 8034 15 8086 75
rect 8344 15 8396 75
rect 8434 15 8486 75
rect 8744 15 8796 75
rect 8834 15 8886 75
rect 9144 15 9196 75
rect 9234 15 9286 75
rect 9544 15 9596 75
rect 9634 15 9686 75
rect 9944 15 9996 75
rect 10034 15 10086 75
rect 10344 15 10396 75
rect 10434 15 10486 75
rect 10744 15 10796 75
rect 10834 15 10886 75
rect 11144 15 11196 75
rect 11234 15 11286 75
rect 11544 15 11596 75
rect 11634 15 11686 75
rect 11944 15 11996 75
rect 12034 15 12086 75
rect 12344 15 12396 75
rect 12434 15 12486 75
rect 12744 15 12796 75
rect 12834 15 12886 75
rect 13144 15 13196 75
rect -366 -50 -330 -35
rect -330 -50 -314 -35
rect -366 -95 -314 -50
rect -56 -95 -4 -35
rect 34 -95 86 -35
rect 344 -95 396 -35
rect 434 -95 486 -35
rect 744 -95 796 -35
rect 834 -95 886 -35
rect 1144 -95 1196 -35
rect 1234 -95 1286 -35
rect 1544 -95 1596 -35
rect 1634 -95 1686 -35
rect 1944 -95 1996 -35
rect 2034 -95 2086 -35
rect 2344 -95 2396 -35
rect 2434 -95 2486 -35
rect 2744 -95 2796 -35
rect 2834 -95 2886 -35
rect 3144 -95 3196 -35
rect 3234 -95 3286 -35
rect 3544 -95 3596 -35
rect 3634 -95 3686 -35
rect 3944 -95 3996 -35
rect 4034 -95 4086 -35
rect 4344 -95 4396 -35
rect 4434 -95 4486 -35
rect 4744 -95 4796 -35
rect 4834 -95 4886 -35
rect 5144 -95 5196 -35
rect 5234 -95 5286 -35
rect 5544 -95 5596 -35
rect 5634 -95 5686 -35
rect 5944 -95 5996 -35
rect 6034 -95 6086 -35
rect 6344 -95 6396 -35
rect 6434 -95 6486 -35
rect 6744 -95 6796 -35
rect 6834 -95 6886 -35
rect 7144 -95 7196 -35
rect 7234 -95 7286 -35
rect 7544 -95 7596 -35
rect 7634 -95 7686 -35
rect 7944 -95 7996 -35
rect 8034 -95 8086 -35
rect 8344 -95 8396 -35
rect 8434 -95 8486 -35
rect 8744 -95 8796 -35
rect 8834 -95 8886 -35
rect 9144 -95 9196 -35
rect 9234 -95 9286 -35
rect 9544 -95 9596 -35
rect 9634 -95 9686 -35
rect 9944 -95 9996 -35
rect 10034 -95 10086 -35
rect 10344 -95 10396 -35
rect 10434 -95 10486 -35
rect 10744 -95 10796 -35
rect 10834 -95 10886 -35
rect 11144 -95 11196 -35
rect 11234 -95 11286 -35
rect 11544 -95 11596 -35
rect 11634 -95 11686 -35
rect 11944 -95 11996 -35
rect 12034 -95 12086 -35
rect 12344 -95 12396 -35
rect 12434 -95 12486 -35
rect 12744 -95 12796 -35
rect 12834 -95 12886 -35
rect 13144 -95 13196 -35
rect -366 -355 -314 -295
rect -56 -355 -4 -295
rect 34 -355 86 -295
rect 344 -355 396 -295
rect 434 -355 486 -295
rect 744 -355 796 -295
rect 834 -355 886 -295
rect 1144 -355 1196 -295
rect 1234 -355 1286 -295
rect 1544 -355 1596 -295
rect 1634 -355 1686 -295
rect 1944 -355 1996 -295
rect 2034 -355 2086 -295
rect 2344 -355 2396 -295
rect 2434 -355 2486 -295
rect 2744 -355 2796 -295
rect 2834 -355 2886 -295
rect 3144 -355 3196 -295
rect 3234 -355 3286 -295
rect 3544 -355 3596 -295
rect 3634 -355 3686 -295
rect 3944 -355 3996 -295
rect 4034 -355 4086 -295
rect 4344 -355 4396 -295
rect 4434 -355 4486 -295
rect 4744 -355 4796 -295
rect 4834 -355 4886 -295
rect 5144 -355 5196 -295
rect 5234 -355 5286 -295
rect 5544 -355 5596 -295
rect 5634 -355 5686 -295
rect 5944 -355 5996 -295
rect 6034 -355 6086 -295
rect 6344 -355 6396 -295
rect 6434 -355 6486 -295
rect 6744 -355 6796 -295
rect 6834 -355 6886 -295
rect 7144 -355 7196 -295
rect 7234 -355 7286 -295
rect 7544 -355 7596 -295
rect 7634 -355 7686 -295
rect 7944 -355 7996 -295
rect 8034 -355 8086 -295
rect 8344 -355 8396 -295
rect 8434 -355 8486 -295
rect 8744 -355 8796 -295
rect 8834 -355 8886 -295
rect 9144 -355 9196 -295
rect 9234 -355 9286 -295
rect 9544 -355 9596 -295
rect 9634 -355 9686 -295
rect 9944 -355 9996 -295
rect 10034 -355 10086 -295
rect 10344 -355 10396 -295
rect 10434 -355 10486 -295
rect 10744 -355 10796 -295
rect 10834 -355 10886 -295
rect 11144 -355 11196 -295
rect 11234 -355 11286 -295
rect 11544 -355 11596 -295
rect 11634 -355 11686 -295
rect 11944 -355 11996 -295
rect 12034 -355 12086 -295
rect 12344 -355 12396 -295
rect 12434 -355 12486 -295
rect 12744 -355 12796 -295
rect 12834 -355 12886 -295
rect 13144 -355 13196 -295
<< metal2 >>
rect -275 24180 -95 24190
rect -275 24120 -265 24180
rect -205 24120 -165 24180
rect -105 24120 -95 24180
rect -275 24110 -95 24120
rect 12915 24125 13105 24135
rect 12990 24065 13030 24125
rect 12915 24055 13105 24065
rect -370 24015 0 24025
rect -370 23955 -366 24015
rect -314 23995 -56 24015
rect -370 23949 -314 23955
rect -370 23761 -340 23949
rect -285 23940 -85 23965
rect -4 23955 0 24015
rect -56 23949 0 23955
rect -285 23920 -215 23940
rect -310 23880 -215 23920
rect -155 23920 -85 23940
rect -155 23880 -60 23920
rect -310 23830 -60 23880
rect -310 23790 -215 23830
rect -285 23770 -215 23790
rect -155 23790 -60 23830
rect -155 23770 -85 23790
rect -370 23755 -314 23761
rect -370 23695 -366 23755
rect -285 23745 -85 23770
rect -30 23761 0 23949
rect -56 23755 0 23761
rect -314 23695 -56 23715
rect -4 23695 0 23755
rect -370 23685 0 23695
rect 30 24015 400 24025
rect 30 23955 34 24015
rect 86 23995 344 24015
rect 30 23949 86 23955
rect 30 23761 60 23949
rect 115 23940 315 23965
rect 396 23955 400 24015
rect 344 23949 400 23955
rect 115 23920 185 23940
rect 90 23880 185 23920
rect 245 23920 315 23940
rect 245 23880 340 23920
rect 90 23830 340 23880
rect 90 23790 185 23830
rect 115 23770 185 23790
rect 245 23790 340 23830
rect 245 23770 315 23790
rect 30 23755 86 23761
rect 30 23695 34 23755
rect 115 23745 315 23770
rect 370 23761 400 23949
rect 344 23755 400 23761
rect 86 23695 344 23715
rect 396 23695 400 23755
rect 30 23685 400 23695
rect 430 24015 800 24025
rect 430 23955 434 24015
rect 486 23995 744 24015
rect 430 23949 486 23955
rect 430 23761 460 23949
rect 515 23940 715 23965
rect 796 23955 800 24015
rect 744 23949 800 23955
rect 515 23920 585 23940
rect 490 23880 585 23920
rect 645 23920 715 23940
rect 645 23880 740 23920
rect 490 23830 740 23880
rect 490 23790 585 23830
rect 515 23770 585 23790
rect 645 23790 740 23830
rect 645 23770 715 23790
rect 430 23755 486 23761
rect 430 23695 434 23755
rect 515 23745 715 23770
rect 770 23761 800 23949
rect 744 23755 800 23761
rect 486 23695 744 23715
rect 796 23695 800 23755
rect 430 23685 800 23695
rect 830 24015 1200 24025
rect 830 23955 834 24015
rect 886 23995 1144 24015
rect 830 23949 886 23955
rect 830 23761 860 23949
rect 915 23940 1115 23965
rect 1196 23955 1200 24015
rect 1144 23949 1200 23955
rect 915 23920 985 23940
rect 890 23880 985 23920
rect 1045 23920 1115 23940
rect 1045 23880 1140 23920
rect 890 23830 1140 23880
rect 890 23790 985 23830
rect 915 23770 985 23790
rect 1045 23790 1140 23830
rect 1045 23770 1115 23790
rect 830 23755 886 23761
rect 830 23695 834 23755
rect 915 23745 1115 23770
rect 1170 23761 1200 23949
rect 1144 23755 1200 23761
rect 886 23695 1144 23715
rect 1196 23695 1200 23755
rect 830 23685 1200 23695
rect 1230 24015 1600 24025
rect 1230 23955 1234 24015
rect 1286 23995 1544 24015
rect 1230 23949 1286 23955
rect 1230 23761 1260 23949
rect 1315 23940 1515 23965
rect 1596 23955 1600 24015
rect 1544 23949 1600 23955
rect 1315 23920 1385 23940
rect 1290 23880 1385 23920
rect 1445 23920 1515 23940
rect 1445 23880 1540 23920
rect 1290 23830 1540 23880
rect 1290 23790 1385 23830
rect 1315 23770 1385 23790
rect 1445 23790 1540 23830
rect 1445 23770 1515 23790
rect 1230 23755 1286 23761
rect 1230 23695 1234 23755
rect 1315 23745 1515 23770
rect 1570 23761 1600 23949
rect 1544 23755 1600 23761
rect 1286 23695 1544 23715
rect 1596 23695 1600 23755
rect 1230 23685 1600 23695
rect 1630 24015 2000 24025
rect 1630 23955 1634 24015
rect 1686 23995 1944 24015
rect 1630 23949 1686 23955
rect 1630 23761 1660 23949
rect 1715 23940 1915 23965
rect 1996 23955 2000 24015
rect 1944 23949 2000 23955
rect 1715 23920 1785 23940
rect 1690 23880 1785 23920
rect 1845 23920 1915 23940
rect 1845 23880 1940 23920
rect 1690 23830 1940 23880
rect 1690 23790 1785 23830
rect 1715 23770 1785 23790
rect 1845 23790 1940 23830
rect 1845 23770 1915 23790
rect 1630 23755 1686 23761
rect 1630 23695 1634 23755
rect 1715 23745 1915 23770
rect 1970 23761 2000 23949
rect 1944 23755 2000 23761
rect 1686 23695 1944 23715
rect 1996 23695 2000 23755
rect 1630 23685 2000 23695
rect 2030 24015 2400 24025
rect 2030 23955 2034 24015
rect 2086 23995 2344 24015
rect 2030 23949 2086 23955
rect 2030 23761 2060 23949
rect 2115 23940 2315 23965
rect 2396 23955 2400 24015
rect 2344 23949 2400 23955
rect 2115 23920 2185 23940
rect 2090 23880 2185 23920
rect 2245 23920 2315 23940
rect 2245 23880 2340 23920
rect 2090 23830 2340 23880
rect 2090 23790 2185 23830
rect 2115 23770 2185 23790
rect 2245 23790 2340 23830
rect 2245 23770 2315 23790
rect 2030 23755 2086 23761
rect 2030 23695 2034 23755
rect 2115 23745 2315 23770
rect 2370 23761 2400 23949
rect 2344 23755 2400 23761
rect 2086 23695 2344 23715
rect 2396 23695 2400 23755
rect 2030 23685 2400 23695
rect 2430 24015 2800 24025
rect 2430 23955 2434 24015
rect 2486 23995 2744 24015
rect 2430 23949 2486 23955
rect 2430 23761 2460 23949
rect 2515 23940 2715 23965
rect 2796 23955 2800 24015
rect 2744 23949 2800 23955
rect 2515 23920 2585 23940
rect 2490 23880 2585 23920
rect 2645 23920 2715 23940
rect 2645 23880 2740 23920
rect 2490 23830 2740 23880
rect 2490 23790 2585 23830
rect 2515 23770 2585 23790
rect 2645 23790 2740 23830
rect 2645 23770 2715 23790
rect 2430 23755 2486 23761
rect 2430 23695 2434 23755
rect 2515 23745 2715 23770
rect 2770 23761 2800 23949
rect 2744 23755 2800 23761
rect 2486 23695 2744 23715
rect 2796 23695 2800 23755
rect 2430 23685 2800 23695
rect 2830 24015 3200 24025
rect 2830 23955 2834 24015
rect 2886 23995 3144 24015
rect 2830 23949 2886 23955
rect 2830 23761 2860 23949
rect 2915 23940 3115 23965
rect 3196 23955 3200 24015
rect 3144 23949 3200 23955
rect 2915 23920 2985 23940
rect 2890 23880 2985 23920
rect 3045 23920 3115 23940
rect 3045 23880 3140 23920
rect 2890 23830 3140 23880
rect 2890 23790 2985 23830
rect 2915 23770 2985 23790
rect 3045 23790 3140 23830
rect 3045 23770 3115 23790
rect 2830 23755 2886 23761
rect 2830 23695 2834 23755
rect 2915 23745 3115 23770
rect 3170 23761 3200 23949
rect 3144 23755 3200 23761
rect 2886 23695 3144 23715
rect 3196 23695 3200 23755
rect 2830 23685 3200 23695
rect 3230 24015 3600 24025
rect 3230 23955 3234 24015
rect 3286 23995 3544 24015
rect 3230 23949 3286 23955
rect 3230 23761 3260 23949
rect 3315 23940 3515 23965
rect 3596 23955 3600 24015
rect 3544 23949 3600 23955
rect 3315 23920 3385 23940
rect 3290 23880 3385 23920
rect 3445 23920 3515 23940
rect 3445 23880 3540 23920
rect 3290 23830 3540 23880
rect 3290 23790 3385 23830
rect 3315 23770 3385 23790
rect 3445 23790 3540 23830
rect 3445 23770 3515 23790
rect 3230 23755 3286 23761
rect 3230 23695 3234 23755
rect 3315 23745 3515 23770
rect 3570 23761 3600 23949
rect 3544 23755 3600 23761
rect 3286 23695 3544 23715
rect 3596 23695 3600 23755
rect 3230 23685 3600 23695
rect 3630 24015 4000 24025
rect 3630 23955 3634 24015
rect 3686 23995 3944 24015
rect 3630 23949 3686 23955
rect 3630 23761 3660 23949
rect 3715 23940 3915 23965
rect 3996 23955 4000 24015
rect 3944 23949 4000 23955
rect 3715 23920 3785 23940
rect 3690 23880 3785 23920
rect 3845 23920 3915 23940
rect 3845 23880 3940 23920
rect 3690 23830 3940 23880
rect 3690 23790 3785 23830
rect 3715 23770 3785 23790
rect 3845 23790 3940 23830
rect 3845 23770 3915 23790
rect 3630 23755 3686 23761
rect 3630 23695 3634 23755
rect 3715 23745 3915 23770
rect 3970 23761 4000 23949
rect 3944 23755 4000 23761
rect 3686 23695 3944 23715
rect 3996 23695 4000 23755
rect 3630 23685 4000 23695
rect 4030 24015 4400 24025
rect 4030 23955 4034 24015
rect 4086 23995 4344 24015
rect 4030 23949 4086 23955
rect 4030 23761 4060 23949
rect 4115 23940 4315 23965
rect 4396 23955 4400 24015
rect 4344 23949 4400 23955
rect 4115 23920 4185 23940
rect 4090 23880 4185 23920
rect 4245 23920 4315 23940
rect 4245 23880 4340 23920
rect 4090 23830 4340 23880
rect 4090 23790 4185 23830
rect 4115 23770 4185 23790
rect 4245 23790 4340 23830
rect 4245 23770 4315 23790
rect 4030 23755 4086 23761
rect 4030 23695 4034 23755
rect 4115 23745 4315 23770
rect 4370 23761 4400 23949
rect 4344 23755 4400 23761
rect 4086 23695 4344 23715
rect 4396 23695 4400 23755
rect 4030 23685 4400 23695
rect 4430 24015 4800 24025
rect 4430 23955 4434 24015
rect 4486 23995 4744 24015
rect 4430 23949 4486 23955
rect 4430 23761 4460 23949
rect 4515 23940 4715 23965
rect 4796 23955 4800 24015
rect 4744 23949 4800 23955
rect 4515 23920 4585 23940
rect 4490 23880 4585 23920
rect 4645 23920 4715 23940
rect 4645 23880 4740 23920
rect 4490 23830 4740 23880
rect 4490 23790 4585 23830
rect 4515 23770 4585 23790
rect 4645 23790 4740 23830
rect 4645 23770 4715 23790
rect 4430 23755 4486 23761
rect 4430 23695 4434 23755
rect 4515 23745 4715 23770
rect 4770 23761 4800 23949
rect 4744 23755 4800 23761
rect 4486 23695 4744 23715
rect 4796 23695 4800 23755
rect 4430 23685 4800 23695
rect 4830 24015 5200 24025
rect 4830 23955 4834 24015
rect 4886 23995 5144 24015
rect 4830 23949 4886 23955
rect 4830 23761 4860 23949
rect 4915 23940 5115 23965
rect 5196 23955 5200 24015
rect 5144 23949 5200 23955
rect 4915 23920 4985 23940
rect 4890 23880 4985 23920
rect 5045 23920 5115 23940
rect 5045 23880 5140 23920
rect 4890 23830 5140 23880
rect 4890 23790 4985 23830
rect 4915 23770 4985 23790
rect 5045 23790 5140 23830
rect 5045 23770 5115 23790
rect 4830 23755 4886 23761
rect 4830 23695 4834 23755
rect 4915 23745 5115 23770
rect 5170 23761 5200 23949
rect 5144 23755 5200 23761
rect 4886 23695 5144 23715
rect 5196 23695 5200 23755
rect 4830 23685 5200 23695
rect 5230 24015 5600 24025
rect 5230 23955 5234 24015
rect 5286 23995 5544 24015
rect 5230 23949 5286 23955
rect 5230 23761 5260 23949
rect 5315 23940 5515 23965
rect 5596 23955 5600 24015
rect 5544 23949 5600 23955
rect 5315 23920 5385 23940
rect 5290 23880 5385 23920
rect 5445 23920 5515 23940
rect 5445 23880 5540 23920
rect 5290 23830 5540 23880
rect 5290 23790 5385 23830
rect 5315 23770 5385 23790
rect 5445 23790 5540 23830
rect 5445 23770 5515 23790
rect 5230 23755 5286 23761
rect 5230 23695 5234 23755
rect 5315 23745 5515 23770
rect 5570 23761 5600 23949
rect 5544 23755 5600 23761
rect 5286 23695 5544 23715
rect 5596 23695 5600 23755
rect 5230 23685 5600 23695
rect 5630 24015 6000 24025
rect 5630 23955 5634 24015
rect 5686 23995 5944 24015
rect 5630 23949 5686 23955
rect 5630 23761 5660 23949
rect 5715 23940 5915 23965
rect 5996 23955 6000 24015
rect 5944 23949 6000 23955
rect 5715 23920 5785 23940
rect 5690 23880 5785 23920
rect 5845 23920 5915 23940
rect 5845 23880 5940 23920
rect 5690 23830 5940 23880
rect 5690 23790 5785 23830
rect 5715 23770 5785 23790
rect 5845 23790 5940 23830
rect 5845 23770 5915 23790
rect 5630 23755 5686 23761
rect 5630 23695 5634 23755
rect 5715 23745 5915 23770
rect 5970 23761 6000 23949
rect 5944 23755 6000 23761
rect 5686 23695 5944 23715
rect 5996 23695 6000 23755
rect 5630 23685 6000 23695
rect 6030 24015 6400 24025
rect 6030 23955 6034 24015
rect 6086 23995 6344 24015
rect 6030 23949 6086 23955
rect 6030 23761 6060 23949
rect 6115 23940 6315 23965
rect 6396 23955 6400 24015
rect 6344 23949 6400 23955
rect 6115 23920 6185 23940
rect 6090 23880 6185 23920
rect 6245 23920 6315 23940
rect 6245 23880 6340 23920
rect 6090 23830 6340 23880
rect 6090 23790 6185 23830
rect 6115 23770 6185 23790
rect 6245 23790 6340 23830
rect 6245 23770 6315 23790
rect 6030 23755 6086 23761
rect 6030 23695 6034 23755
rect 6115 23745 6315 23770
rect 6370 23761 6400 23949
rect 6344 23755 6400 23761
rect 6086 23695 6344 23715
rect 6396 23695 6400 23755
rect 6030 23685 6400 23695
rect 6430 24015 6800 24025
rect 6430 23955 6434 24015
rect 6486 23995 6744 24015
rect 6430 23949 6486 23955
rect 6430 23761 6460 23949
rect 6515 23940 6715 23965
rect 6796 23955 6800 24015
rect 6744 23949 6800 23955
rect 6515 23920 6585 23940
rect 6490 23880 6585 23920
rect 6645 23920 6715 23940
rect 6645 23880 6740 23920
rect 6490 23830 6740 23880
rect 6490 23790 6585 23830
rect 6515 23770 6585 23790
rect 6645 23790 6740 23830
rect 6645 23770 6715 23790
rect 6430 23755 6486 23761
rect 6430 23695 6434 23755
rect 6515 23745 6715 23770
rect 6770 23761 6800 23949
rect 6744 23755 6800 23761
rect 6486 23695 6744 23715
rect 6796 23695 6800 23755
rect 6430 23685 6800 23695
rect 6830 24015 7200 24025
rect 6830 23955 6834 24015
rect 6886 23995 7144 24015
rect 6830 23949 6886 23955
rect 6830 23761 6860 23949
rect 6915 23940 7115 23965
rect 7196 23955 7200 24015
rect 7144 23949 7200 23955
rect 6915 23920 6985 23940
rect 6890 23880 6985 23920
rect 7045 23920 7115 23940
rect 7045 23880 7140 23920
rect 6890 23830 7140 23880
rect 6890 23790 6985 23830
rect 6915 23770 6985 23790
rect 7045 23790 7140 23830
rect 7045 23770 7115 23790
rect 6830 23755 6886 23761
rect 6830 23695 6834 23755
rect 6915 23745 7115 23770
rect 7170 23761 7200 23949
rect 7144 23755 7200 23761
rect 6886 23695 7144 23715
rect 7196 23695 7200 23755
rect 6830 23685 7200 23695
rect 7230 24015 7600 24025
rect 7230 23955 7234 24015
rect 7286 23995 7544 24015
rect 7230 23949 7286 23955
rect 7230 23761 7260 23949
rect 7315 23940 7515 23965
rect 7596 23955 7600 24015
rect 7544 23949 7600 23955
rect 7315 23920 7385 23940
rect 7290 23880 7385 23920
rect 7445 23920 7515 23940
rect 7445 23880 7540 23920
rect 7290 23830 7540 23880
rect 7290 23790 7385 23830
rect 7315 23770 7385 23790
rect 7445 23790 7540 23830
rect 7445 23770 7515 23790
rect 7230 23755 7286 23761
rect 7230 23695 7234 23755
rect 7315 23745 7515 23770
rect 7570 23761 7600 23949
rect 7544 23755 7600 23761
rect 7286 23695 7544 23715
rect 7596 23695 7600 23755
rect 7230 23685 7600 23695
rect 7630 24015 8000 24025
rect 7630 23955 7634 24015
rect 7686 23995 7944 24015
rect 7630 23949 7686 23955
rect 7630 23761 7660 23949
rect 7715 23940 7915 23965
rect 7996 23955 8000 24015
rect 7944 23949 8000 23955
rect 7715 23920 7785 23940
rect 7690 23880 7785 23920
rect 7845 23920 7915 23940
rect 7845 23880 7940 23920
rect 7690 23830 7940 23880
rect 7690 23790 7785 23830
rect 7715 23770 7785 23790
rect 7845 23790 7940 23830
rect 7845 23770 7915 23790
rect 7630 23755 7686 23761
rect 7630 23695 7634 23755
rect 7715 23745 7915 23770
rect 7970 23761 8000 23949
rect 7944 23755 8000 23761
rect 7686 23695 7944 23715
rect 7996 23695 8000 23755
rect 7630 23685 8000 23695
rect 8030 24015 8400 24025
rect 8030 23955 8034 24015
rect 8086 23995 8344 24015
rect 8030 23949 8086 23955
rect 8030 23761 8060 23949
rect 8115 23940 8315 23965
rect 8396 23955 8400 24015
rect 8344 23949 8400 23955
rect 8115 23920 8185 23940
rect 8090 23880 8185 23920
rect 8245 23920 8315 23940
rect 8245 23880 8340 23920
rect 8090 23830 8340 23880
rect 8090 23790 8185 23830
rect 8115 23770 8185 23790
rect 8245 23790 8340 23830
rect 8245 23770 8315 23790
rect 8030 23755 8086 23761
rect 8030 23695 8034 23755
rect 8115 23745 8315 23770
rect 8370 23761 8400 23949
rect 8344 23755 8400 23761
rect 8086 23695 8344 23715
rect 8396 23695 8400 23755
rect 8030 23685 8400 23695
rect 8430 24015 8800 24025
rect 8430 23955 8434 24015
rect 8486 23995 8744 24015
rect 8430 23949 8486 23955
rect 8430 23761 8460 23949
rect 8515 23940 8715 23965
rect 8796 23955 8800 24015
rect 8744 23949 8800 23955
rect 8515 23920 8585 23940
rect 8490 23880 8585 23920
rect 8645 23920 8715 23940
rect 8645 23880 8740 23920
rect 8490 23830 8740 23880
rect 8490 23790 8585 23830
rect 8515 23770 8585 23790
rect 8645 23790 8740 23830
rect 8645 23770 8715 23790
rect 8430 23755 8486 23761
rect 8430 23695 8434 23755
rect 8515 23745 8715 23770
rect 8770 23761 8800 23949
rect 8744 23755 8800 23761
rect 8486 23695 8744 23715
rect 8796 23695 8800 23755
rect 8430 23685 8800 23695
rect 8830 24015 9200 24025
rect 8830 23955 8834 24015
rect 8886 23995 9144 24015
rect 8830 23949 8886 23955
rect 8830 23761 8860 23949
rect 8915 23940 9115 23965
rect 9196 23955 9200 24015
rect 9144 23949 9200 23955
rect 8915 23920 8985 23940
rect 8890 23880 8985 23920
rect 9045 23920 9115 23940
rect 9045 23880 9140 23920
rect 8890 23830 9140 23880
rect 8890 23790 8985 23830
rect 8915 23770 8985 23790
rect 9045 23790 9140 23830
rect 9045 23770 9115 23790
rect 8830 23755 8886 23761
rect 8830 23695 8834 23755
rect 8915 23745 9115 23770
rect 9170 23761 9200 23949
rect 9144 23755 9200 23761
rect 8886 23695 9144 23715
rect 9196 23695 9200 23755
rect 8830 23685 9200 23695
rect 9230 24015 9600 24025
rect 9230 23955 9234 24015
rect 9286 23995 9544 24015
rect 9230 23949 9286 23955
rect 9230 23761 9260 23949
rect 9315 23940 9515 23965
rect 9596 23955 9600 24015
rect 9544 23949 9600 23955
rect 9315 23920 9385 23940
rect 9290 23880 9385 23920
rect 9445 23920 9515 23940
rect 9445 23880 9540 23920
rect 9290 23830 9540 23880
rect 9290 23790 9385 23830
rect 9315 23770 9385 23790
rect 9445 23790 9540 23830
rect 9445 23770 9515 23790
rect 9230 23755 9286 23761
rect 9230 23695 9234 23755
rect 9315 23745 9515 23770
rect 9570 23761 9600 23949
rect 9544 23755 9600 23761
rect 9286 23695 9544 23715
rect 9596 23695 9600 23755
rect 9230 23685 9600 23695
rect 9630 24015 10000 24025
rect 9630 23955 9634 24015
rect 9686 23995 9944 24015
rect 9630 23949 9686 23955
rect 9630 23761 9660 23949
rect 9715 23940 9915 23965
rect 9996 23955 10000 24015
rect 9944 23949 10000 23955
rect 9715 23920 9785 23940
rect 9690 23880 9785 23920
rect 9845 23920 9915 23940
rect 9845 23880 9940 23920
rect 9690 23830 9940 23880
rect 9690 23790 9785 23830
rect 9715 23770 9785 23790
rect 9845 23790 9940 23830
rect 9845 23770 9915 23790
rect 9630 23755 9686 23761
rect 9630 23695 9634 23755
rect 9715 23745 9915 23770
rect 9970 23761 10000 23949
rect 9944 23755 10000 23761
rect 9686 23695 9944 23715
rect 9996 23695 10000 23755
rect 9630 23685 10000 23695
rect 10030 24015 10400 24025
rect 10030 23955 10034 24015
rect 10086 23995 10344 24015
rect 10030 23949 10086 23955
rect 10030 23761 10060 23949
rect 10115 23940 10315 23965
rect 10396 23955 10400 24015
rect 10344 23949 10400 23955
rect 10115 23920 10185 23940
rect 10090 23880 10185 23920
rect 10245 23920 10315 23940
rect 10245 23880 10340 23920
rect 10090 23830 10340 23880
rect 10090 23790 10185 23830
rect 10115 23770 10185 23790
rect 10245 23790 10340 23830
rect 10245 23770 10315 23790
rect 10030 23755 10086 23761
rect 10030 23695 10034 23755
rect 10115 23745 10315 23770
rect 10370 23761 10400 23949
rect 10344 23755 10400 23761
rect 10086 23695 10344 23715
rect 10396 23695 10400 23755
rect 10030 23685 10400 23695
rect 10430 24015 10800 24025
rect 10430 23955 10434 24015
rect 10486 23995 10744 24015
rect 10430 23949 10486 23955
rect 10430 23761 10460 23949
rect 10515 23940 10715 23965
rect 10796 23955 10800 24015
rect 10744 23949 10800 23955
rect 10515 23920 10585 23940
rect 10490 23880 10585 23920
rect 10645 23920 10715 23940
rect 10645 23880 10740 23920
rect 10490 23830 10740 23880
rect 10490 23790 10585 23830
rect 10515 23770 10585 23790
rect 10645 23790 10740 23830
rect 10645 23770 10715 23790
rect 10430 23755 10486 23761
rect 10430 23695 10434 23755
rect 10515 23745 10715 23770
rect 10770 23761 10800 23949
rect 10744 23755 10800 23761
rect 10486 23695 10744 23715
rect 10796 23695 10800 23755
rect 10430 23685 10800 23695
rect 10830 24015 11200 24025
rect 10830 23955 10834 24015
rect 10886 23995 11144 24015
rect 10830 23949 10886 23955
rect 10830 23761 10860 23949
rect 10915 23940 11115 23965
rect 11196 23955 11200 24015
rect 11144 23949 11200 23955
rect 10915 23920 10985 23940
rect 10890 23880 10985 23920
rect 11045 23920 11115 23940
rect 11045 23880 11140 23920
rect 10890 23830 11140 23880
rect 10890 23790 10985 23830
rect 10915 23770 10985 23790
rect 11045 23790 11140 23830
rect 11045 23770 11115 23790
rect 10830 23755 10886 23761
rect 10830 23695 10834 23755
rect 10915 23745 11115 23770
rect 11170 23761 11200 23949
rect 11144 23755 11200 23761
rect 10886 23695 11144 23715
rect 11196 23695 11200 23755
rect 10830 23685 11200 23695
rect 11230 24015 11600 24025
rect 11230 23955 11234 24015
rect 11286 23995 11544 24015
rect 11230 23949 11286 23955
rect 11230 23761 11260 23949
rect 11315 23940 11515 23965
rect 11596 23955 11600 24015
rect 11544 23949 11600 23955
rect 11315 23920 11385 23940
rect 11290 23880 11385 23920
rect 11445 23920 11515 23940
rect 11445 23880 11540 23920
rect 11290 23830 11540 23880
rect 11290 23790 11385 23830
rect 11315 23770 11385 23790
rect 11445 23790 11540 23830
rect 11445 23770 11515 23790
rect 11230 23755 11286 23761
rect 11230 23695 11234 23755
rect 11315 23745 11515 23770
rect 11570 23761 11600 23949
rect 11544 23755 11600 23761
rect 11286 23695 11544 23715
rect 11596 23695 11600 23755
rect 11230 23685 11600 23695
rect 11630 24015 12000 24025
rect 11630 23955 11634 24015
rect 11686 23995 11944 24015
rect 11630 23949 11686 23955
rect 11630 23761 11660 23949
rect 11715 23940 11915 23965
rect 11996 23955 12000 24015
rect 11944 23949 12000 23955
rect 11715 23920 11785 23940
rect 11690 23880 11785 23920
rect 11845 23920 11915 23940
rect 11845 23880 11940 23920
rect 11690 23830 11940 23880
rect 11690 23790 11785 23830
rect 11715 23770 11785 23790
rect 11845 23790 11940 23830
rect 11845 23770 11915 23790
rect 11630 23755 11686 23761
rect 11630 23695 11634 23755
rect 11715 23745 11915 23770
rect 11970 23761 12000 23949
rect 11944 23755 12000 23761
rect 11686 23695 11944 23715
rect 11996 23695 12000 23755
rect 11630 23685 12000 23695
rect 12030 24015 12400 24025
rect 12030 23955 12034 24015
rect 12086 23995 12344 24015
rect 12030 23949 12086 23955
rect 12030 23761 12060 23949
rect 12115 23940 12315 23965
rect 12396 23955 12400 24015
rect 12344 23949 12400 23955
rect 12115 23920 12185 23940
rect 12090 23880 12185 23920
rect 12245 23920 12315 23940
rect 12245 23880 12340 23920
rect 12090 23830 12340 23880
rect 12090 23790 12185 23830
rect 12115 23770 12185 23790
rect 12245 23790 12340 23830
rect 12245 23770 12315 23790
rect 12030 23755 12086 23761
rect 12030 23695 12034 23755
rect 12115 23745 12315 23770
rect 12370 23761 12400 23949
rect 12344 23755 12400 23761
rect 12086 23695 12344 23715
rect 12396 23695 12400 23755
rect 12030 23685 12400 23695
rect 12430 24015 12800 24025
rect 12430 23955 12434 24015
rect 12486 23995 12744 24015
rect 12430 23949 12486 23955
rect 12430 23761 12460 23949
rect 12515 23940 12715 23965
rect 12796 23955 12800 24015
rect 12744 23949 12800 23955
rect 12515 23920 12585 23940
rect 12490 23880 12585 23920
rect 12645 23920 12715 23940
rect 12645 23880 12740 23920
rect 12490 23830 12740 23880
rect 12490 23790 12585 23830
rect 12515 23770 12585 23790
rect 12645 23790 12740 23830
rect 12645 23770 12715 23790
rect 12430 23755 12486 23761
rect 12430 23695 12434 23755
rect 12515 23745 12715 23770
rect 12770 23761 12800 23949
rect 12744 23755 12800 23761
rect 12486 23695 12744 23715
rect 12796 23695 12800 23755
rect 12430 23685 12800 23695
rect 12830 24015 13200 24025
rect 12830 23955 12834 24015
rect 12886 23995 13144 24015
rect 12830 23949 12886 23955
rect 12830 23761 12860 23949
rect 12915 23940 13115 23965
rect 13196 23955 13200 24015
rect 13144 23949 13200 23955
rect 12915 23920 12985 23940
rect 12890 23880 12985 23920
rect 13045 23920 13115 23940
rect 13045 23880 13140 23920
rect 12890 23830 13140 23880
rect 12890 23790 12985 23830
rect 12915 23770 12985 23790
rect 13045 23790 13140 23830
rect 13045 23770 13115 23790
rect 12830 23755 12886 23761
rect 12830 23695 12834 23755
rect 12915 23745 13115 23770
rect 13170 23761 13200 23949
rect 13144 23755 13200 23761
rect 12886 23695 13144 23715
rect 13196 23695 13200 23755
rect 12830 23685 13200 23695
rect -370 23645 0 23655
rect -370 23585 -366 23645
rect -314 23625 -56 23645
rect -370 23579 -314 23585
rect -370 23391 -340 23579
rect -285 23570 -85 23595
rect -4 23585 0 23645
rect -56 23579 0 23585
rect -285 23550 -215 23570
rect -310 23510 -215 23550
rect -155 23550 -85 23570
rect -155 23510 -60 23550
rect -310 23460 -60 23510
rect -310 23420 -215 23460
rect -285 23400 -215 23420
rect -155 23420 -60 23460
rect -155 23400 -85 23420
rect -370 23385 -314 23391
rect -370 23325 -366 23385
rect -285 23375 -85 23400
rect -30 23391 0 23579
rect -56 23385 0 23391
rect -314 23325 -56 23345
rect -4 23325 0 23385
rect -370 23315 0 23325
rect 30 23645 400 23655
rect 30 23585 34 23645
rect 86 23625 344 23645
rect 30 23579 86 23585
rect 30 23391 60 23579
rect 115 23570 315 23595
rect 396 23585 400 23645
rect 344 23579 400 23585
rect 115 23550 185 23570
rect 90 23510 185 23550
rect 245 23550 315 23570
rect 245 23510 340 23550
rect 90 23460 340 23510
rect 90 23420 185 23460
rect 115 23400 185 23420
rect 245 23420 340 23460
rect 245 23400 315 23420
rect 30 23385 86 23391
rect 30 23325 34 23385
rect 115 23375 315 23400
rect 370 23391 400 23579
rect 344 23385 400 23391
rect 86 23325 344 23345
rect 396 23325 400 23385
rect 30 23315 400 23325
rect 430 23645 800 23655
rect 430 23585 434 23645
rect 486 23625 744 23645
rect 430 23579 486 23585
rect 430 23391 460 23579
rect 515 23570 715 23595
rect 796 23585 800 23645
rect 744 23579 800 23585
rect 515 23550 585 23570
rect 490 23510 585 23550
rect 645 23550 715 23570
rect 645 23510 740 23550
rect 490 23460 740 23510
rect 490 23420 585 23460
rect 515 23400 585 23420
rect 645 23420 740 23460
rect 645 23400 715 23420
rect 430 23385 486 23391
rect 430 23325 434 23385
rect 515 23375 715 23400
rect 770 23391 800 23579
rect 744 23385 800 23391
rect 486 23325 744 23345
rect 796 23325 800 23385
rect 430 23315 800 23325
rect 830 23645 1200 23655
rect 830 23585 834 23645
rect 886 23625 1144 23645
rect 830 23579 886 23585
rect 830 23391 860 23579
rect 915 23570 1115 23595
rect 1196 23585 1200 23645
rect 1144 23579 1200 23585
rect 915 23550 985 23570
rect 890 23510 985 23550
rect 1045 23550 1115 23570
rect 1045 23510 1140 23550
rect 890 23460 1140 23510
rect 890 23420 985 23460
rect 915 23400 985 23420
rect 1045 23420 1140 23460
rect 1045 23400 1115 23420
rect 830 23385 886 23391
rect 830 23325 834 23385
rect 915 23375 1115 23400
rect 1170 23391 1200 23579
rect 1144 23385 1200 23391
rect 886 23325 1144 23345
rect 1196 23325 1200 23385
rect 830 23315 1200 23325
rect 1230 23645 1600 23655
rect 1230 23585 1234 23645
rect 1286 23625 1544 23645
rect 1230 23579 1286 23585
rect 1230 23391 1260 23579
rect 1315 23570 1515 23595
rect 1596 23585 1600 23645
rect 1544 23579 1600 23585
rect 1315 23550 1385 23570
rect 1290 23510 1385 23550
rect 1445 23550 1515 23570
rect 1445 23510 1540 23550
rect 1290 23460 1540 23510
rect 1290 23420 1385 23460
rect 1315 23400 1385 23420
rect 1445 23420 1540 23460
rect 1445 23400 1515 23420
rect 1230 23385 1286 23391
rect 1230 23325 1234 23385
rect 1315 23375 1515 23400
rect 1570 23391 1600 23579
rect 1544 23385 1600 23391
rect 1286 23325 1544 23345
rect 1596 23325 1600 23385
rect 1230 23315 1600 23325
rect 1630 23645 2000 23655
rect 1630 23585 1634 23645
rect 1686 23625 1944 23645
rect 1630 23579 1686 23585
rect 1630 23391 1660 23579
rect 1715 23570 1915 23595
rect 1996 23585 2000 23645
rect 1944 23579 2000 23585
rect 1715 23550 1785 23570
rect 1690 23510 1785 23550
rect 1845 23550 1915 23570
rect 1845 23510 1940 23550
rect 1690 23460 1940 23510
rect 1690 23420 1785 23460
rect 1715 23400 1785 23420
rect 1845 23420 1940 23460
rect 1845 23400 1915 23420
rect 1630 23385 1686 23391
rect 1630 23325 1634 23385
rect 1715 23375 1915 23400
rect 1970 23391 2000 23579
rect 1944 23385 2000 23391
rect 1686 23325 1944 23345
rect 1996 23325 2000 23385
rect 1630 23315 2000 23325
rect 2030 23645 2400 23655
rect 2030 23585 2034 23645
rect 2086 23625 2344 23645
rect 2030 23579 2086 23585
rect 2030 23391 2060 23579
rect 2115 23570 2315 23595
rect 2396 23585 2400 23645
rect 2344 23579 2400 23585
rect 2115 23550 2185 23570
rect 2090 23510 2185 23550
rect 2245 23550 2315 23570
rect 2245 23510 2340 23550
rect 2090 23460 2340 23510
rect 2090 23420 2185 23460
rect 2115 23400 2185 23420
rect 2245 23420 2340 23460
rect 2245 23400 2315 23420
rect 2030 23385 2086 23391
rect 2030 23325 2034 23385
rect 2115 23375 2315 23400
rect 2370 23391 2400 23579
rect 2344 23385 2400 23391
rect 2086 23325 2344 23345
rect 2396 23325 2400 23385
rect 2030 23315 2400 23325
rect 2430 23645 2800 23655
rect 2430 23585 2434 23645
rect 2486 23625 2744 23645
rect 2430 23579 2486 23585
rect 2430 23391 2460 23579
rect 2515 23570 2715 23595
rect 2796 23585 2800 23645
rect 2744 23579 2800 23585
rect 2515 23550 2585 23570
rect 2490 23510 2585 23550
rect 2645 23550 2715 23570
rect 2645 23510 2740 23550
rect 2490 23460 2740 23510
rect 2490 23420 2585 23460
rect 2515 23400 2585 23420
rect 2645 23420 2740 23460
rect 2645 23400 2715 23420
rect 2430 23385 2486 23391
rect 2430 23325 2434 23385
rect 2515 23375 2715 23400
rect 2770 23391 2800 23579
rect 2744 23385 2800 23391
rect 2486 23325 2744 23345
rect 2796 23325 2800 23385
rect 2430 23315 2800 23325
rect 2830 23645 3200 23655
rect 2830 23585 2834 23645
rect 2886 23625 3144 23645
rect 2830 23579 2886 23585
rect 2830 23391 2860 23579
rect 2915 23570 3115 23595
rect 3196 23585 3200 23645
rect 3144 23579 3200 23585
rect 2915 23550 2985 23570
rect 2890 23510 2985 23550
rect 3045 23550 3115 23570
rect 3045 23510 3140 23550
rect 2890 23460 3140 23510
rect 2890 23420 2985 23460
rect 2915 23400 2985 23420
rect 3045 23420 3140 23460
rect 3045 23400 3115 23420
rect 2830 23385 2886 23391
rect 2830 23325 2834 23385
rect 2915 23375 3115 23400
rect 3170 23391 3200 23579
rect 3144 23385 3200 23391
rect 2886 23325 3144 23345
rect 3196 23325 3200 23385
rect 2830 23315 3200 23325
rect 3230 23645 3600 23655
rect 3230 23585 3234 23645
rect 3286 23625 3544 23645
rect 3230 23579 3286 23585
rect 3230 23391 3260 23579
rect 3315 23570 3515 23595
rect 3596 23585 3600 23645
rect 3544 23579 3600 23585
rect 3315 23550 3385 23570
rect 3290 23510 3385 23550
rect 3445 23550 3515 23570
rect 3445 23510 3540 23550
rect 3290 23460 3540 23510
rect 3290 23420 3385 23460
rect 3315 23400 3385 23420
rect 3445 23420 3540 23460
rect 3445 23400 3515 23420
rect 3230 23385 3286 23391
rect 3230 23325 3234 23385
rect 3315 23375 3515 23400
rect 3570 23391 3600 23579
rect 3544 23385 3600 23391
rect 3286 23325 3544 23345
rect 3596 23325 3600 23385
rect 3230 23315 3600 23325
rect 3630 23645 4000 23655
rect 3630 23585 3634 23645
rect 3686 23625 3944 23645
rect 3630 23579 3686 23585
rect 3630 23391 3660 23579
rect 3715 23570 3915 23595
rect 3996 23585 4000 23645
rect 3944 23579 4000 23585
rect 3715 23550 3785 23570
rect 3690 23510 3785 23550
rect 3845 23550 3915 23570
rect 3845 23510 3940 23550
rect 3690 23460 3940 23510
rect 3690 23420 3785 23460
rect 3715 23400 3785 23420
rect 3845 23420 3940 23460
rect 3845 23400 3915 23420
rect 3630 23385 3686 23391
rect 3630 23325 3634 23385
rect 3715 23375 3915 23400
rect 3970 23391 4000 23579
rect 3944 23385 4000 23391
rect 3686 23325 3944 23345
rect 3996 23325 4000 23385
rect 3630 23315 4000 23325
rect 4030 23645 4400 23655
rect 4030 23585 4034 23645
rect 4086 23625 4344 23645
rect 4030 23579 4086 23585
rect 4030 23391 4060 23579
rect 4115 23570 4315 23595
rect 4396 23585 4400 23645
rect 4344 23579 4400 23585
rect 4115 23550 4185 23570
rect 4090 23510 4185 23550
rect 4245 23550 4315 23570
rect 4245 23510 4340 23550
rect 4090 23460 4340 23510
rect 4090 23420 4185 23460
rect 4115 23400 4185 23420
rect 4245 23420 4340 23460
rect 4245 23400 4315 23420
rect 4030 23385 4086 23391
rect 4030 23325 4034 23385
rect 4115 23375 4315 23400
rect 4370 23391 4400 23579
rect 4344 23385 4400 23391
rect 4086 23325 4344 23345
rect 4396 23325 4400 23385
rect 4030 23315 4400 23325
rect 4430 23645 4800 23655
rect 4430 23585 4434 23645
rect 4486 23625 4744 23645
rect 4430 23579 4486 23585
rect 4430 23391 4460 23579
rect 4515 23570 4715 23595
rect 4796 23585 4800 23645
rect 4744 23579 4800 23585
rect 4515 23550 4585 23570
rect 4490 23510 4585 23550
rect 4645 23550 4715 23570
rect 4645 23510 4740 23550
rect 4490 23460 4740 23510
rect 4490 23420 4585 23460
rect 4515 23400 4585 23420
rect 4645 23420 4740 23460
rect 4645 23400 4715 23420
rect 4430 23385 4486 23391
rect 4430 23325 4434 23385
rect 4515 23375 4715 23400
rect 4770 23391 4800 23579
rect 4744 23385 4800 23391
rect 4486 23325 4744 23345
rect 4796 23325 4800 23385
rect 4430 23315 4800 23325
rect 4830 23645 5200 23655
rect 4830 23585 4834 23645
rect 4886 23625 5144 23645
rect 4830 23579 4886 23585
rect 4830 23391 4860 23579
rect 4915 23570 5115 23595
rect 5196 23585 5200 23645
rect 5144 23579 5200 23585
rect 4915 23550 4985 23570
rect 4890 23510 4985 23550
rect 5045 23550 5115 23570
rect 5045 23510 5140 23550
rect 4890 23460 5140 23510
rect 4890 23420 4985 23460
rect 4915 23400 4985 23420
rect 5045 23420 5140 23460
rect 5045 23400 5115 23420
rect 4830 23385 4886 23391
rect 4830 23325 4834 23385
rect 4915 23375 5115 23400
rect 5170 23391 5200 23579
rect 5144 23385 5200 23391
rect 4886 23325 5144 23345
rect 5196 23325 5200 23385
rect 4830 23315 5200 23325
rect 5230 23645 5600 23655
rect 5230 23585 5234 23645
rect 5286 23625 5544 23645
rect 5230 23579 5286 23585
rect 5230 23391 5260 23579
rect 5315 23570 5515 23595
rect 5596 23585 5600 23645
rect 5544 23579 5600 23585
rect 5315 23550 5385 23570
rect 5290 23510 5385 23550
rect 5445 23550 5515 23570
rect 5445 23510 5540 23550
rect 5290 23460 5540 23510
rect 5290 23420 5385 23460
rect 5315 23400 5385 23420
rect 5445 23420 5540 23460
rect 5445 23400 5515 23420
rect 5230 23385 5286 23391
rect 5230 23325 5234 23385
rect 5315 23375 5515 23400
rect 5570 23391 5600 23579
rect 5544 23385 5600 23391
rect 5286 23325 5544 23345
rect 5596 23325 5600 23385
rect 5230 23315 5600 23325
rect 5630 23645 6000 23655
rect 5630 23585 5634 23645
rect 5686 23625 5944 23645
rect 5630 23579 5686 23585
rect 5630 23391 5660 23579
rect 5715 23570 5915 23595
rect 5996 23585 6000 23645
rect 5944 23579 6000 23585
rect 5715 23550 5785 23570
rect 5690 23510 5785 23550
rect 5845 23550 5915 23570
rect 5845 23510 5940 23550
rect 5690 23460 5940 23510
rect 5690 23420 5785 23460
rect 5715 23400 5785 23420
rect 5845 23420 5940 23460
rect 5845 23400 5915 23420
rect 5630 23385 5686 23391
rect 5630 23325 5634 23385
rect 5715 23375 5915 23400
rect 5970 23391 6000 23579
rect 5944 23385 6000 23391
rect 5686 23325 5944 23345
rect 5996 23325 6000 23385
rect 5630 23315 6000 23325
rect 6030 23645 6400 23655
rect 6030 23585 6034 23645
rect 6086 23625 6344 23645
rect 6030 23579 6086 23585
rect 6030 23391 6060 23579
rect 6115 23570 6315 23595
rect 6396 23585 6400 23645
rect 6344 23579 6400 23585
rect 6115 23550 6185 23570
rect 6090 23510 6185 23550
rect 6245 23550 6315 23570
rect 6245 23510 6340 23550
rect 6090 23460 6340 23510
rect 6090 23420 6185 23460
rect 6115 23400 6185 23420
rect 6245 23420 6340 23460
rect 6245 23400 6315 23420
rect 6030 23385 6086 23391
rect 6030 23325 6034 23385
rect 6115 23375 6315 23400
rect 6370 23391 6400 23579
rect 6344 23385 6400 23391
rect 6086 23325 6344 23345
rect 6396 23325 6400 23385
rect 6030 23315 6400 23325
rect 6430 23645 6800 23655
rect 6430 23585 6434 23645
rect 6486 23625 6744 23645
rect 6430 23579 6486 23585
rect 6430 23391 6460 23579
rect 6515 23570 6715 23595
rect 6796 23585 6800 23645
rect 6744 23579 6800 23585
rect 6515 23550 6585 23570
rect 6490 23510 6585 23550
rect 6645 23550 6715 23570
rect 6645 23510 6740 23550
rect 6490 23460 6740 23510
rect 6490 23420 6585 23460
rect 6515 23400 6585 23420
rect 6645 23420 6740 23460
rect 6645 23400 6715 23420
rect 6430 23385 6486 23391
rect 6430 23325 6434 23385
rect 6515 23375 6715 23400
rect 6770 23391 6800 23579
rect 6744 23385 6800 23391
rect 6486 23325 6744 23345
rect 6796 23325 6800 23385
rect 6430 23315 6800 23325
rect 6830 23645 7200 23655
rect 6830 23585 6834 23645
rect 6886 23625 7144 23645
rect 6830 23579 6886 23585
rect 6830 23391 6860 23579
rect 6915 23570 7115 23595
rect 7196 23585 7200 23645
rect 7144 23579 7200 23585
rect 6915 23550 6985 23570
rect 6890 23510 6985 23550
rect 7045 23550 7115 23570
rect 7045 23510 7140 23550
rect 6890 23460 7140 23510
rect 6890 23420 6985 23460
rect 6915 23400 6985 23420
rect 7045 23420 7140 23460
rect 7045 23400 7115 23420
rect 6830 23385 6886 23391
rect 6830 23325 6834 23385
rect 6915 23375 7115 23400
rect 7170 23391 7200 23579
rect 7144 23385 7200 23391
rect 6886 23325 7144 23345
rect 7196 23325 7200 23385
rect 6830 23315 7200 23325
rect 7230 23645 7600 23655
rect 7230 23585 7234 23645
rect 7286 23625 7544 23645
rect 7230 23579 7286 23585
rect 7230 23391 7260 23579
rect 7315 23570 7515 23595
rect 7596 23585 7600 23645
rect 7544 23579 7600 23585
rect 7315 23550 7385 23570
rect 7290 23510 7385 23550
rect 7445 23550 7515 23570
rect 7445 23510 7540 23550
rect 7290 23460 7540 23510
rect 7290 23420 7385 23460
rect 7315 23400 7385 23420
rect 7445 23420 7540 23460
rect 7445 23400 7515 23420
rect 7230 23385 7286 23391
rect 7230 23325 7234 23385
rect 7315 23375 7515 23400
rect 7570 23391 7600 23579
rect 7544 23385 7600 23391
rect 7286 23325 7544 23345
rect 7596 23325 7600 23385
rect 7230 23315 7600 23325
rect 7630 23645 8000 23655
rect 7630 23585 7634 23645
rect 7686 23625 7944 23645
rect 7630 23579 7686 23585
rect 7630 23391 7660 23579
rect 7715 23570 7915 23595
rect 7996 23585 8000 23645
rect 7944 23579 8000 23585
rect 7715 23550 7785 23570
rect 7690 23510 7785 23550
rect 7845 23550 7915 23570
rect 7845 23510 7940 23550
rect 7690 23460 7940 23510
rect 7690 23420 7785 23460
rect 7715 23400 7785 23420
rect 7845 23420 7940 23460
rect 7845 23400 7915 23420
rect 7630 23385 7686 23391
rect 7630 23325 7634 23385
rect 7715 23375 7915 23400
rect 7970 23391 8000 23579
rect 7944 23385 8000 23391
rect 7686 23325 7944 23345
rect 7996 23325 8000 23385
rect 7630 23315 8000 23325
rect 8030 23645 8400 23655
rect 8030 23585 8034 23645
rect 8086 23625 8344 23645
rect 8030 23579 8086 23585
rect 8030 23391 8060 23579
rect 8115 23570 8315 23595
rect 8396 23585 8400 23645
rect 8344 23579 8400 23585
rect 8115 23550 8185 23570
rect 8090 23510 8185 23550
rect 8245 23550 8315 23570
rect 8245 23510 8340 23550
rect 8090 23460 8340 23510
rect 8090 23420 8185 23460
rect 8115 23400 8185 23420
rect 8245 23420 8340 23460
rect 8245 23400 8315 23420
rect 8030 23385 8086 23391
rect 8030 23325 8034 23385
rect 8115 23375 8315 23400
rect 8370 23391 8400 23579
rect 8344 23385 8400 23391
rect 8086 23325 8344 23345
rect 8396 23325 8400 23385
rect 8030 23315 8400 23325
rect 8430 23645 8800 23655
rect 8430 23585 8434 23645
rect 8486 23625 8744 23645
rect 8430 23579 8486 23585
rect 8430 23391 8460 23579
rect 8515 23570 8715 23595
rect 8796 23585 8800 23645
rect 8744 23579 8800 23585
rect 8515 23550 8585 23570
rect 8490 23510 8585 23550
rect 8645 23550 8715 23570
rect 8645 23510 8740 23550
rect 8490 23460 8740 23510
rect 8490 23420 8585 23460
rect 8515 23400 8585 23420
rect 8645 23420 8740 23460
rect 8645 23400 8715 23420
rect 8430 23385 8486 23391
rect 8430 23325 8434 23385
rect 8515 23375 8715 23400
rect 8770 23391 8800 23579
rect 8744 23385 8800 23391
rect 8486 23325 8744 23345
rect 8796 23325 8800 23385
rect 8430 23315 8800 23325
rect 8830 23645 9200 23655
rect 8830 23585 8834 23645
rect 8886 23625 9144 23645
rect 8830 23579 8886 23585
rect 8830 23391 8860 23579
rect 8915 23570 9115 23595
rect 9196 23585 9200 23645
rect 9144 23579 9200 23585
rect 8915 23550 8985 23570
rect 8890 23510 8985 23550
rect 9045 23550 9115 23570
rect 9045 23510 9140 23550
rect 8890 23460 9140 23510
rect 8890 23420 8985 23460
rect 8915 23400 8985 23420
rect 9045 23420 9140 23460
rect 9045 23400 9115 23420
rect 8830 23385 8886 23391
rect 8830 23325 8834 23385
rect 8915 23375 9115 23400
rect 9170 23391 9200 23579
rect 9144 23385 9200 23391
rect 8886 23325 9144 23345
rect 9196 23325 9200 23385
rect 8830 23315 9200 23325
rect 9230 23645 9600 23655
rect 9230 23585 9234 23645
rect 9286 23625 9544 23645
rect 9230 23579 9286 23585
rect 9230 23391 9260 23579
rect 9315 23570 9515 23595
rect 9596 23585 9600 23645
rect 9544 23579 9600 23585
rect 9315 23550 9385 23570
rect 9290 23510 9385 23550
rect 9445 23550 9515 23570
rect 9445 23510 9540 23550
rect 9290 23460 9540 23510
rect 9290 23420 9385 23460
rect 9315 23400 9385 23420
rect 9445 23420 9540 23460
rect 9445 23400 9515 23420
rect 9230 23385 9286 23391
rect 9230 23325 9234 23385
rect 9315 23375 9515 23400
rect 9570 23391 9600 23579
rect 9544 23385 9600 23391
rect 9286 23325 9544 23345
rect 9596 23325 9600 23385
rect 9230 23315 9600 23325
rect 9630 23645 10000 23655
rect 9630 23585 9634 23645
rect 9686 23625 9944 23645
rect 9630 23579 9686 23585
rect 9630 23391 9660 23579
rect 9715 23570 9915 23595
rect 9996 23585 10000 23645
rect 9944 23579 10000 23585
rect 9715 23550 9785 23570
rect 9690 23510 9785 23550
rect 9845 23550 9915 23570
rect 9845 23510 9940 23550
rect 9690 23460 9940 23510
rect 9690 23420 9785 23460
rect 9715 23400 9785 23420
rect 9845 23420 9940 23460
rect 9845 23400 9915 23420
rect 9630 23385 9686 23391
rect 9630 23325 9634 23385
rect 9715 23375 9915 23400
rect 9970 23391 10000 23579
rect 9944 23385 10000 23391
rect 9686 23325 9944 23345
rect 9996 23325 10000 23385
rect 9630 23315 10000 23325
rect 10030 23645 10400 23655
rect 10030 23585 10034 23645
rect 10086 23625 10344 23645
rect 10030 23579 10086 23585
rect 10030 23391 10060 23579
rect 10115 23570 10315 23595
rect 10396 23585 10400 23645
rect 10344 23579 10400 23585
rect 10115 23550 10185 23570
rect 10090 23510 10185 23550
rect 10245 23550 10315 23570
rect 10245 23510 10340 23550
rect 10090 23460 10340 23510
rect 10090 23420 10185 23460
rect 10115 23400 10185 23420
rect 10245 23420 10340 23460
rect 10245 23400 10315 23420
rect 10030 23385 10086 23391
rect 10030 23325 10034 23385
rect 10115 23375 10315 23400
rect 10370 23391 10400 23579
rect 10344 23385 10400 23391
rect 10086 23325 10344 23345
rect 10396 23325 10400 23385
rect 10030 23315 10400 23325
rect 10430 23645 10800 23655
rect 10430 23585 10434 23645
rect 10486 23625 10744 23645
rect 10430 23579 10486 23585
rect 10430 23391 10460 23579
rect 10515 23570 10715 23595
rect 10796 23585 10800 23645
rect 10744 23579 10800 23585
rect 10515 23550 10585 23570
rect 10490 23510 10585 23550
rect 10645 23550 10715 23570
rect 10645 23510 10740 23550
rect 10490 23460 10740 23510
rect 10490 23420 10585 23460
rect 10515 23400 10585 23420
rect 10645 23420 10740 23460
rect 10645 23400 10715 23420
rect 10430 23385 10486 23391
rect 10430 23325 10434 23385
rect 10515 23375 10715 23400
rect 10770 23391 10800 23579
rect 10744 23385 10800 23391
rect 10486 23325 10744 23345
rect 10796 23325 10800 23385
rect 10430 23315 10800 23325
rect 10830 23645 11200 23655
rect 10830 23585 10834 23645
rect 10886 23625 11144 23645
rect 10830 23579 10886 23585
rect 10830 23391 10860 23579
rect 10915 23570 11115 23595
rect 11196 23585 11200 23645
rect 11144 23579 11200 23585
rect 10915 23550 10985 23570
rect 10890 23510 10985 23550
rect 11045 23550 11115 23570
rect 11045 23510 11140 23550
rect 10890 23460 11140 23510
rect 10890 23420 10985 23460
rect 10915 23400 10985 23420
rect 11045 23420 11140 23460
rect 11045 23400 11115 23420
rect 10830 23385 10886 23391
rect 10830 23325 10834 23385
rect 10915 23375 11115 23400
rect 11170 23391 11200 23579
rect 11144 23385 11200 23391
rect 10886 23325 11144 23345
rect 11196 23325 11200 23385
rect 10830 23315 11200 23325
rect 11230 23645 11600 23655
rect 11230 23585 11234 23645
rect 11286 23625 11544 23645
rect 11230 23579 11286 23585
rect 11230 23391 11260 23579
rect 11315 23570 11515 23595
rect 11596 23585 11600 23645
rect 11544 23579 11600 23585
rect 11315 23550 11385 23570
rect 11290 23510 11385 23550
rect 11445 23550 11515 23570
rect 11445 23510 11540 23550
rect 11290 23460 11540 23510
rect 11290 23420 11385 23460
rect 11315 23400 11385 23420
rect 11445 23420 11540 23460
rect 11445 23400 11515 23420
rect 11230 23385 11286 23391
rect 11230 23325 11234 23385
rect 11315 23375 11515 23400
rect 11570 23391 11600 23579
rect 11544 23385 11600 23391
rect 11286 23325 11544 23345
rect 11596 23325 11600 23385
rect 11230 23315 11600 23325
rect 11630 23645 12000 23655
rect 11630 23585 11634 23645
rect 11686 23625 11944 23645
rect 11630 23579 11686 23585
rect 11630 23391 11660 23579
rect 11715 23570 11915 23595
rect 11996 23585 12000 23645
rect 11944 23579 12000 23585
rect 11715 23550 11785 23570
rect 11690 23510 11785 23550
rect 11845 23550 11915 23570
rect 11845 23510 11940 23550
rect 11690 23460 11940 23510
rect 11690 23420 11785 23460
rect 11715 23400 11785 23420
rect 11845 23420 11940 23460
rect 11845 23400 11915 23420
rect 11630 23385 11686 23391
rect 11630 23325 11634 23385
rect 11715 23375 11915 23400
rect 11970 23391 12000 23579
rect 11944 23385 12000 23391
rect 11686 23325 11944 23345
rect 11996 23325 12000 23385
rect 11630 23315 12000 23325
rect 12030 23645 12400 23655
rect 12030 23585 12034 23645
rect 12086 23625 12344 23645
rect 12030 23579 12086 23585
rect 12030 23391 12060 23579
rect 12115 23570 12315 23595
rect 12396 23585 12400 23645
rect 12344 23579 12400 23585
rect 12115 23550 12185 23570
rect 12090 23510 12185 23550
rect 12245 23550 12315 23570
rect 12245 23510 12340 23550
rect 12090 23460 12340 23510
rect 12090 23420 12185 23460
rect 12115 23400 12185 23420
rect 12245 23420 12340 23460
rect 12245 23400 12315 23420
rect 12030 23385 12086 23391
rect 12030 23325 12034 23385
rect 12115 23375 12315 23400
rect 12370 23391 12400 23579
rect 12344 23385 12400 23391
rect 12086 23325 12344 23345
rect 12396 23325 12400 23385
rect 12030 23315 12400 23325
rect 12430 23645 12800 23655
rect 12430 23585 12434 23645
rect 12486 23625 12744 23645
rect 12430 23579 12486 23585
rect 12430 23391 12460 23579
rect 12515 23570 12715 23595
rect 12796 23585 12800 23645
rect 12744 23579 12800 23585
rect 12515 23550 12585 23570
rect 12490 23510 12585 23550
rect 12645 23550 12715 23570
rect 12645 23510 12740 23550
rect 12490 23460 12740 23510
rect 12490 23420 12585 23460
rect 12515 23400 12585 23420
rect 12645 23420 12740 23460
rect 12645 23400 12715 23420
rect 12430 23385 12486 23391
rect 12430 23325 12434 23385
rect 12515 23375 12715 23400
rect 12770 23391 12800 23579
rect 12744 23385 12800 23391
rect 12486 23325 12744 23345
rect 12796 23325 12800 23385
rect 12430 23315 12800 23325
rect 12830 23645 13200 23655
rect 12830 23585 12834 23645
rect 12886 23625 13144 23645
rect 12830 23579 12886 23585
rect 12830 23391 12860 23579
rect 12915 23570 13115 23595
rect 13196 23585 13200 23645
rect 13144 23579 13200 23585
rect 12915 23550 12985 23570
rect 12890 23510 12985 23550
rect 13045 23550 13115 23570
rect 13045 23510 13140 23550
rect 12890 23460 13140 23510
rect 12890 23420 12985 23460
rect 12915 23400 12985 23420
rect 13045 23420 13140 23460
rect 13045 23400 13115 23420
rect 12830 23385 12886 23391
rect 12830 23325 12834 23385
rect 12915 23375 13115 23400
rect 13170 23391 13200 23579
rect 13144 23385 13200 23391
rect 12886 23325 13144 23345
rect 13196 23325 13200 23385
rect 12830 23315 13200 23325
rect -370 23275 0 23285
rect -370 23215 -366 23275
rect -314 23255 -56 23275
rect -370 23209 -314 23215
rect -370 23021 -340 23209
rect -285 23200 -85 23225
rect -4 23215 0 23275
rect -56 23209 0 23215
rect -285 23180 -215 23200
rect -310 23140 -215 23180
rect -155 23180 -85 23200
rect -155 23140 -60 23180
rect -310 23090 -60 23140
rect -310 23050 -215 23090
rect -285 23030 -215 23050
rect -155 23050 -60 23090
rect -155 23030 -85 23050
rect -370 23015 -314 23021
rect -370 22955 -366 23015
rect -285 23005 -85 23030
rect -30 23021 0 23209
rect -56 23015 0 23021
rect -314 22955 -56 22975
rect -4 22955 0 23015
rect -370 22945 0 22955
rect 30 23275 400 23285
rect 30 23215 34 23275
rect 86 23255 344 23275
rect 30 23209 86 23215
rect 30 23021 60 23209
rect 115 23200 315 23225
rect 396 23215 400 23275
rect 344 23209 400 23215
rect 115 23180 185 23200
rect 90 23140 185 23180
rect 245 23180 315 23200
rect 245 23140 340 23180
rect 90 23090 340 23140
rect 90 23050 185 23090
rect 115 23030 185 23050
rect 245 23050 340 23090
rect 245 23030 315 23050
rect 30 23015 86 23021
rect 30 22955 34 23015
rect 115 23005 315 23030
rect 370 23021 400 23209
rect 344 23015 400 23021
rect 86 22955 344 22975
rect 396 22955 400 23015
rect 30 22945 400 22955
rect 430 23275 800 23285
rect 430 23215 434 23275
rect 486 23255 744 23275
rect 430 23209 486 23215
rect 430 23021 460 23209
rect 515 23200 715 23225
rect 796 23215 800 23275
rect 744 23209 800 23215
rect 515 23180 585 23200
rect 490 23140 585 23180
rect 645 23180 715 23200
rect 645 23140 740 23180
rect 490 23090 740 23140
rect 490 23050 585 23090
rect 515 23030 585 23050
rect 645 23050 740 23090
rect 645 23030 715 23050
rect 430 23015 486 23021
rect 430 22955 434 23015
rect 515 23005 715 23030
rect 770 23021 800 23209
rect 744 23015 800 23021
rect 486 22955 744 22975
rect 796 22955 800 23015
rect 430 22945 800 22955
rect 830 23275 1200 23285
rect 830 23215 834 23275
rect 886 23255 1144 23275
rect 830 23209 886 23215
rect 830 23021 860 23209
rect 915 23200 1115 23225
rect 1196 23215 1200 23275
rect 1144 23209 1200 23215
rect 915 23180 985 23200
rect 890 23140 985 23180
rect 1045 23180 1115 23200
rect 1045 23140 1140 23180
rect 890 23090 1140 23140
rect 890 23050 985 23090
rect 915 23030 985 23050
rect 1045 23050 1140 23090
rect 1045 23030 1115 23050
rect 830 23015 886 23021
rect 830 22955 834 23015
rect 915 23005 1115 23030
rect 1170 23021 1200 23209
rect 1144 23015 1200 23021
rect 886 22955 1144 22975
rect 1196 22955 1200 23015
rect 830 22945 1200 22955
rect 1230 23275 1600 23285
rect 1230 23215 1234 23275
rect 1286 23255 1544 23275
rect 1230 23209 1286 23215
rect 1230 23021 1260 23209
rect 1315 23200 1515 23225
rect 1596 23215 1600 23275
rect 1544 23209 1600 23215
rect 1315 23180 1385 23200
rect 1290 23140 1385 23180
rect 1445 23180 1515 23200
rect 1445 23140 1540 23180
rect 1290 23090 1540 23140
rect 1290 23050 1385 23090
rect 1315 23030 1385 23050
rect 1445 23050 1540 23090
rect 1445 23030 1515 23050
rect 1230 23015 1286 23021
rect 1230 22955 1234 23015
rect 1315 23005 1515 23030
rect 1570 23021 1600 23209
rect 1544 23015 1600 23021
rect 1286 22955 1544 22975
rect 1596 22955 1600 23015
rect 1230 22945 1600 22955
rect 1630 23275 2000 23285
rect 1630 23215 1634 23275
rect 1686 23255 1944 23275
rect 1630 23209 1686 23215
rect 1630 23021 1660 23209
rect 1715 23200 1915 23225
rect 1996 23215 2000 23275
rect 1944 23209 2000 23215
rect 1715 23180 1785 23200
rect 1690 23140 1785 23180
rect 1845 23180 1915 23200
rect 1845 23140 1940 23180
rect 1690 23090 1940 23140
rect 1690 23050 1785 23090
rect 1715 23030 1785 23050
rect 1845 23050 1940 23090
rect 1845 23030 1915 23050
rect 1630 23015 1686 23021
rect 1630 22955 1634 23015
rect 1715 23005 1915 23030
rect 1970 23021 2000 23209
rect 1944 23015 2000 23021
rect 1686 22955 1944 22975
rect 1996 22955 2000 23015
rect 1630 22945 2000 22955
rect 2030 23275 2400 23285
rect 2030 23215 2034 23275
rect 2086 23255 2344 23275
rect 2030 23209 2086 23215
rect 2030 23021 2060 23209
rect 2115 23200 2315 23225
rect 2396 23215 2400 23275
rect 2344 23209 2400 23215
rect 2115 23180 2185 23200
rect 2090 23140 2185 23180
rect 2245 23180 2315 23200
rect 2245 23140 2340 23180
rect 2090 23090 2340 23140
rect 2090 23050 2185 23090
rect 2115 23030 2185 23050
rect 2245 23050 2340 23090
rect 2245 23030 2315 23050
rect 2030 23015 2086 23021
rect 2030 22955 2034 23015
rect 2115 23005 2315 23030
rect 2370 23021 2400 23209
rect 2344 23015 2400 23021
rect 2086 22955 2344 22975
rect 2396 22955 2400 23015
rect 2030 22945 2400 22955
rect 2430 23275 2800 23285
rect 2430 23215 2434 23275
rect 2486 23255 2744 23275
rect 2430 23209 2486 23215
rect 2430 23021 2460 23209
rect 2515 23200 2715 23225
rect 2796 23215 2800 23275
rect 2744 23209 2800 23215
rect 2515 23180 2585 23200
rect 2490 23140 2585 23180
rect 2645 23180 2715 23200
rect 2645 23140 2740 23180
rect 2490 23090 2740 23140
rect 2490 23050 2585 23090
rect 2515 23030 2585 23050
rect 2645 23050 2740 23090
rect 2645 23030 2715 23050
rect 2430 23015 2486 23021
rect 2430 22955 2434 23015
rect 2515 23005 2715 23030
rect 2770 23021 2800 23209
rect 2744 23015 2800 23021
rect 2486 22955 2744 22975
rect 2796 22955 2800 23015
rect 2430 22945 2800 22955
rect 2830 23275 3200 23285
rect 2830 23215 2834 23275
rect 2886 23255 3144 23275
rect 2830 23209 2886 23215
rect 2830 23021 2860 23209
rect 2915 23200 3115 23225
rect 3196 23215 3200 23275
rect 3144 23209 3200 23215
rect 2915 23180 2985 23200
rect 2890 23140 2985 23180
rect 3045 23180 3115 23200
rect 3045 23140 3140 23180
rect 2890 23090 3140 23140
rect 2890 23050 2985 23090
rect 2915 23030 2985 23050
rect 3045 23050 3140 23090
rect 3045 23030 3115 23050
rect 2830 23015 2886 23021
rect 2830 22955 2834 23015
rect 2915 23005 3115 23030
rect 3170 23021 3200 23209
rect 3144 23015 3200 23021
rect 2886 22955 3144 22975
rect 3196 22955 3200 23015
rect 2830 22945 3200 22955
rect 3230 23275 3600 23285
rect 3230 23215 3234 23275
rect 3286 23255 3544 23275
rect 3230 23209 3286 23215
rect 3230 23021 3260 23209
rect 3315 23200 3515 23225
rect 3596 23215 3600 23275
rect 3544 23209 3600 23215
rect 3315 23180 3385 23200
rect 3290 23140 3385 23180
rect 3445 23180 3515 23200
rect 3445 23140 3540 23180
rect 3290 23090 3540 23140
rect 3290 23050 3385 23090
rect 3315 23030 3385 23050
rect 3445 23050 3540 23090
rect 3445 23030 3515 23050
rect 3230 23015 3286 23021
rect 3230 22955 3234 23015
rect 3315 23005 3515 23030
rect 3570 23021 3600 23209
rect 3544 23015 3600 23021
rect 3286 22955 3544 22975
rect 3596 22955 3600 23015
rect 3230 22945 3600 22955
rect 3630 23275 4000 23285
rect 3630 23215 3634 23275
rect 3686 23255 3944 23275
rect 3630 23209 3686 23215
rect 3630 23021 3660 23209
rect 3715 23200 3915 23225
rect 3996 23215 4000 23275
rect 3944 23209 4000 23215
rect 3715 23180 3785 23200
rect 3690 23140 3785 23180
rect 3845 23180 3915 23200
rect 3845 23140 3940 23180
rect 3690 23090 3940 23140
rect 3690 23050 3785 23090
rect 3715 23030 3785 23050
rect 3845 23050 3940 23090
rect 3845 23030 3915 23050
rect 3630 23015 3686 23021
rect 3630 22955 3634 23015
rect 3715 23005 3915 23030
rect 3970 23021 4000 23209
rect 3944 23015 4000 23021
rect 3686 22955 3944 22975
rect 3996 22955 4000 23015
rect 3630 22945 4000 22955
rect 4030 23275 4400 23285
rect 4030 23215 4034 23275
rect 4086 23255 4344 23275
rect 4030 23209 4086 23215
rect 4030 23021 4060 23209
rect 4115 23200 4315 23225
rect 4396 23215 4400 23275
rect 4344 23209 4400 23215
rect 4115 23180 4185 23200
rect 4090 23140 4185 23180
rect 4245 23180 4315 23200
rect 4245 23140 4340 23180
rect 4090 23090 4340 23140
rect 4090 23050 4185 23090
rect 4115 23030 4185 23050
rect 4245 23050 4340 23090
rect 4245 23030 4315 23050
rect 4030 23015 4086 23021
rect 4030 22955 4034 23015
rect 4115 23005 4315 23030
rect 4370 23021 4400 23209
rect 4344 23015 4400 23021
rect 4086 22955 4344 22975
rect 4396 22955 4400 23015
rect 4030 22945 4400 22955
rect 4430 23275 4800 23285
rect 4430 23215 4434 23275
rect 4486 23255 4744 23275
rect 4430 23209 4486 23215
rect 4430 23021 4460 23209
rect 4515 23200 4715 23225
rect 4796 23215 4800 23275
rect 4744 23209 4800 23215
rect 4515 23180 4585 23200
rect 4490 23140 4585 23180
rect 4645 23180 4715 23200
rect 4645 23140 4740 23180
rect 4490 23090 4740 23140
rect 4490 23050 4585 23090
rect 4515 23030 4585 23050
rect 4645 23050 4740 23090
rect 4645 23030 4715 23050
rect 4430 23015 4486 23021
rect 4430 22955 4434 23015
rect 4515 23005 4715 23030
rect 4770 23021 4800 23209
rect 4744 23015 4800 23021
rect 4486 22955 4744 22975
rect 4796 22955 4800 23015
rect 4430 22945 4800 22955
rect 4830 23275 5200 23285
rect 4830 23215 4834 23275
rect 4886 23255 5144 23275
rect 4830 23209 4886 23215
rect 4830 23021 4860 23209
rect 4915 23200 5115 23225
rect 5196 23215 5200 23275
rect 5144 23209 5200 23215
rect 4915 23180 4985 23200
rect 4890 23140 4985 23180
rect 5045 23180 5115 23200
rect 5045 23140 5140 23180
rect 4890 23090 5140 23140
rect 4890 23050 4985 23090
rect 4915 23030 4985 23050
rect 5045 23050 5140 23090
rect 5045 23030 5115 23050
rect 4830 23015 4886 23021
rect 4830 22955 4834 23015
rect 4915 23005 5115 23030
rect 5170 23021 5200 23209
rect 5144 23015 5200 23021
rect 4886 22955 5144 22975
rect 5196 22955 5200 23015
rect 4830 22945 5200 22955
rect 5230 23275 5600 23285
rect 5230 23215 5234 23275
rect 5286 23255 5544 23275
rect 5230 23209 5286 23215
rect 5230 23021 5260 23209
rect 5315 23200 5515 23225
rect 5596 23215 5600 23275
rect 5544 23209 5600 23215
rect 5315 23180 5385 23200
rect 5290 23140 5385 23180
rect 5445 23180 5515 23200
rect 5445 23140 5540 23180
rect 5290 23090 5540 23140
rect 5290 23050 5385 23090
rect 5315 23030 5385 23050
rect 5445 23050 5540 23090
rect 5445 23030 5515 23050
rect 5230 23015 5286 23021
rect 5230 22955 5234 23015
rect 5315 23005 5515 23030
rect 5570 23021 5600 23209
rect 5544 23015 5600 23021
rect 5286 22955 5544 22975
rect 5596 22955 5600 23015
rect 5230 22945 5600 22955
rect 5630 23275 6000 23285
rect 5630 23215 5634 23275
rect 5686 23255 5944 23275
rect 5630 23209 5686 23215
rect 5630 23021 5660 23209
rect 5715 23200 5915 23225
rect 5996 23215 6000 23275
rect 5944 23209 6000 23215
rect 5715 23180 5785 23200
rect 5690 23140 5785 23180
rect 5845 23180 5915 23200
rect 5845 23140 5940 23180
rect 5690 23090 5940 23140
rect 5690 23050 5785 23090
rect 5715 23030 5785 23050
rect 5845 23050 5940 23090
rect 5845 23030 5915 23050
rect 5630 23015 5686 23021
rect 5630 22955 5634 23015
rect 5715 23005 5915 23030
rect 5970 23021 6000 23209
rect 5944 23015 6000 23021
rect 5686 22955 5944 22975
rect 5996 22955 6000 23015
rect 5630 22945 6000 22955
rect 6030 23275 6400 23285
rect 6030 23215 6034 23275
rect 6086 23255 6344 23275
rect 6030 23209 6086 23215
rect 6030 23021 6060 23209
rect 6115 23200 6315 23225
rect 6396 23215 6400 23275
rect 6344 23209 6400 23215
rect 6115 23180 6185 23200
rect 6090 23140 6185 23180
rect 6245 23180 6315 23200
rect 6245 23140 6340 23180
rect 6090 23090 6340 23140
rect 6090 23050 6185 23090
rect 6115 23030 6185 23050
rect 6245 23050 6340 23090
rect 6245 23030 6315 23050
rect 6030 23015 6086 23021
rect 6030 22955 6034 23015
rect 6115 23005 6315 23030
rect 6370 23021 6400 23209
rect 6344 23015 6400 23021
rect 6086 22955 6344 22975
rect 6396 22955 6400 23015
rect 6030 22945 6400 22955
rect 6430 23275 6800 23285
rect 6430 23215 6434 23275
rect 6486 23255 6744 23275
rect 6430 23209 6486 23215
rect 6430 23021 6460 23209
rect 6515 23200 6715 23225
rect 6796 23215 6800 23275
rect 6744 23209 6800 23215
rect 6515 23180 6585 23200
rect 6490 23140 6585 23180
rect 6645 23180 6715 23200
rect 6645 23140 6740 23180
rect 6490 23090 6740 23140
rect 6490 23050 6585 23090
rect 6515 23030 6585 23050
rect 6645 23050 6740 23090
rect 6645 23030 6715 23050
rect 6430 23015 6486 23021
rect 6430 22955 6434 23015
rect 6515 23005 6715 23030
rect 6770 23021 6800 23209
rect 6744 23015 6800 23021
rect 6486 22955 6744 22975
rect 6796 22955 6800 23015
rect 6430 22945 6800 22955
rect 6830 23275 7200 23285
rect 6830 23215 6834 23275
rect 6886 23255 7144 23275
rect 6830 23209 6886 23215
rect 6830 23021 6860 23209
rect 6915 23200 7115 23225
rect 7196 23215 7200 23275
rect 7144 23209 7200 23215
rect 6915 23180 6985 23200
rect 6890 23140 6985 23180
rect 7045 23180 7115 23200
rect 7045 23140 7140 23180
rect 6890 23090 7140 23140
rect 6890 23050 6985 23090
rect 6915 23030 6985 23050
rect 7045 23050 7140 23090
rect 7045 23030 7115 23050
rect 6830 23015 6886 23021
rect 6830 22955 6834 23015
rect 6915 23005 7115 23030
rect 7170 23021 7200 23209
rect 7144 23015 7200 23021
rect 6886 22955 7144 22975
rect 7196 22955 7200 23015
rect 6830 22945 7200 22955
rect 7230 23275 7600 23285
rect 7230 23215 7234 23275
rect 7286 23255 7544 23275
rect 7230 23209 7286 23215
rect 7230 23021 7260 23209
rect 7315 23200 7515 23225
rect 7596 23215 7600 23275
rect 7544 23209 7600 23215
rect 7315 23180 7385 23200
rect 7290 23140 7385 23180
rect 7445 23180 7515 23200
rect 7445 23140 7540 23180
rect 7290 23090 7540 23140
rect 7290 23050 7385 23090
rect 7315 23030 7385 23050
rect 7445 23050 7540 23090
rect 7445 23030 7515 23050
rect 7230 23015 7286 23021
rect 7230 22955 7234 23015
rect 7315 23005 7515 23030
rect 7570 23021 7600 23209
rect 7544 23015 7600 23021
rect 7286 22955 7544 22975
rect 7596 22955 7600 23015
rect 7230 22945 7600 22955
rect 7630 23275 8000 23285
rect 7630 23215 7634 23275
rect 7686 23255 7944 23275
rect 7630 23209 7686 23215
rect 7630 23021 7660 23209
rect 7715 23200 7915 23225
rect 7996 23215 8000 23275
rect 7944 23209 8000 23215
rect 7715 23180 7785 23200
rect 7690 23140 7785 23180
rect 7845 23180 7915 23200
rect 7845 23140 7940 23180
rect 7690 23090 7940 23140
rect 7690 23050 7785 23090
rect 7715 23030 7785 23050
rect 7845 23050 7940 23090
rect 7845 23030 7915 23050
rect 7630 23015 7686 23021
rect 7630 22955 7634 23015
rect 7715 23005 7915 23030
rect 7970 23021 8000 23209
rect 7944 23015 8000 23021
rect 7686 22955 7944 22975
rect 7996 22955 8000 23015
rect 7630 22945 8000 22955
rect 8030 23275 8400 23285
rect 8030 23215 8034 23275
rect 8086 23255 8344 23275
rect 8030 23209 8086 23215
rect 8030 23021 8060 23209
rect 8115 23200 8315 23225
rect 8396 23215 8400 23275
rect 8344 23209 8400 23215
rect 8115 23180 8185 23200
rect 8090 23140 8185 23180
rect 8245 23180 8315 23200
rect 8245 23140 8340 23180
rect 8090 23090 8340 23140
rect 8090 23050 8185 23090
rect 8115 23030 8185 23050
rect 8245 23050 8340 23090
rect 8245 23030 8315 23050
rect 8030 23015 8086 23021
rect 8030 22955 8034 23015
rect 8115 23005 8315 23030
rect 8370 23021 8400 23209
rect 8344 23015 8400 23021
rect 8086 22955 8344 22975
rect 8396 22955 8400 23015
rect 8030 22945 8400 22955
rect 8430 23275 8800 23285
rect 8430 23215 8434 23275
rect 8486 23255 8744 23275
rect 8430 23209 8486 23215
rect 8430 23021 8460 23209
rect 8515 23200 8715 23225
rect 8796 23215 8800 23275
rect 8744 23209 8800 23215
rect 8515 23180 8585 23200
rect 8490 23140 8585 23180
rect 8645 23180 8715 23200
rect 8645 23140 8740 23180
rect 8490 23090 8740 23140
rect 8490 23050 8585 23090
rect 8515 23030 8585 23050
rect 8645 23050 8740 23090
rect 8645 23030 8715 23050
rect 8430 23015 8486 23021
rect 8430 22955 8434 23015
rect 8515 23005 8715 23030
rect 8770 23021 8800 23209
rect 8744 23015 8800 23021
rect 8486 22955 8744 22975
rect 8796 22955 8800 23015
rect 8430 22945 8800 22955
rect 8830 23275 9200 23285
rect 8830 23215 8834 23275
rect 8886 23255 9144 23275
rect 8830 23209 8886 23215
rect 8830 23021 8860 23209
rect 8915 23200 9115 23225
rect 9196 23215 9200 23275
rect 9144 23209 9200 23215
rect 8915 23180 8985 23200
rect 8890 23140 8985 23180
rect 9045 23180 9115 23200
rect 9045 23140 9140 23180
rect 8890 23090 9140 23140
rect 8890 23050 8985 23090
rect 8915 23030 8985 23050
rect 9045 23050 9140 23090
rect 9045 23030 9115 23050
rect 8830 23015 8886 23021
rect 8830 22955 8834 23015
rect 8915 23005 9115 23030
rect 9170 23021 9200 23209
rect 9144 23015 9200 23021
rect 8886 22955 9144 22975
rect 9196 22955 9200 23015
rect 8830 22945 9200 22955
rect 9230 23275 9600 23285
rect 9230 23215 9234 23275
rect 9286 23255 9544 23275
rect 9230 23209 9286 23215
rect 9230 23021 9260 23209
rect 9315 23200 9515 23225
rect 9596 23215 9600 23275
rect 9544 23209 9600 23215
rect 9315 23180 9385 23200
rect 9290 23140 9385 23180
rect 9445 23180 9515 23200
rect 9445 23140 9540 23180
rect 9290 23090 9540 23140
rect 9290 23050 9385 23090
rect 9315 23030 9385 23050
rect 9445 23050 9540 23090
rect 9445 23030 9515 23050
rect 9230 23015 9286 23021
rect 9230 22955 9234 23015
rect 9315 23005 9515 23030
rect 9570 23021 9600 23209
rect 9544 23015 9600 23021
rect 9286 22955 9544 22975
rect 9596 22955 9600 23015
rect 9230 22945 9600 22955
rect 9630 23275 10000 23285
rect 9630 23215 9634 23275
rect 9686 23255 9944 23275
rect 9630 23209 9686 23215
rect 9630 23021 9660 23209
rect 9715 23200 9915 23225
rect 9996 23215 10000 23275
rect 9944 23209 10000 23215
rect 9715 23180 9785 23200
rect 9690 23140 9785 23180
rect 9845 23180 9915 23200
rect 9845 23140 9940 23180
rect 9690 23090 9940 23140
rect 9690 23050 9785 23090
rect 9715 23030 9785 23050
rect 9845 23050 9940 23090
rect 9845 23030 9915 23050
rect 9630 23015 9686 23021
rect 9630 22955 9634 23015
rect 9715 23005 9915 23030
rect 9970 23021 10000 23209
rect 9944 23015 10000 23021
rect 9686 22955 9944 22975
rect 9996 22955 10000 23015
rect 9630 22945 10000 22955
rect 10030 23275 10400 23285
rect 10030 23215 10034 23275
rect 10086 23255 10344 23275
rect 10030 23209 10086 23215
rect 10030 23021 10060 23209
rect 10115 23200 10315 23225
rect 10396 23215 10400 23275
rect 10344 23209 10400 23215
rect 10115 23180 10185 23200
rect 10090 23140 10185 23180
rect 10245 23180 10315 23200
rect 10245 23140 10340 23180
rect 10090 23090 10340 23140
rect 10090 23050 10185 23090
rect 10115 23030 10185 23050
rect 10245 23050 10340 23090
rect 10245 23030 10315 23050
rect 10030 23015 10086 23021
rect 10030 22955 10034 23015
rect 10115 23005 10315 23030
rect 10370 23021 10400 23209
rect 10344 23015 10400 23021
rect 10086 22955 10344 22975
rect 10396 22955 10400 23015
rect 10030 22945 10400 22955
rect 10430 23275 10800 23285
rect 10430 23215 10434 23275
rect 10486 23255 10744 23275
rect 10430 23209 10486 23215
rect 10430 23021 10460 23209
rect 10515 23200 10715 23225
rect 10796 23215 10800 23275
rect 10744 23209 10800 23215
rect 10515 23180 10585 23200
rect 10490 23140 10585 23180
rect 10645 23180 10715 23200
rect 10645 23140 10740 23180
rect 10490 23090 10740 23140
rect 10490 23050 10585 23090
rect 10515 23030 10585 23050
rect 10645 23050 10740 23090
rect 10645 23030 10715 23050
rect 10430 23015 10486 23021
rect 10430 22955 10434 23015
rect 10515 23005 10715 23030
rect 10770 23021 10800 23209
rect 10744 23015 10800 23021
rect 10486 22955 10744 22975
rect 10796 22955 10800 23015
rect 10430 22945 10800 22955
rect 10830 23275 11200 23285
rect 10830 23215 10834 23275
rect 10886 23255 11144 23275
rect 10830 23209 10886 23215
rect 10830 23021 10860 23209
rect 10915 23200 11115 23225
rect 11196 23215 11200 23275
rect 11144 23209 11200 23215
rect 10915 23180 10985 23200
rect 10890 23140 10985 23180
rect 11045 23180 11115 23200
rect 11045 23140 11140 23180
rect 10890 23090 11140 23140
rect 10890 23050 10985 23090
rect 10915 23030 10985 23050
rect 11045 23050 11140 23090
rect 11045 23030 11115 23050
rect 10830 23015 10886 23021
rect 10830 22955 10834 23015
rect 10915 23005 11115 23030
rect 11170 23021 11200 23209
rect 11144 23015 11200 23021
rect 10886 22955 11144 22975
rect 11196 22955 11200 23015
rect 10830 22945 11200 22955
rect 11230 23275 11600 23285
rect 11230 23215 11234 23275
rect 11286 23255 11544 23275
rect 11230 23209 11286 23215
rect 11230 23021 11260 23209
rect 11315 23200 11515 23225
rect 11596 23215 11600 23275
rect 11544 23209 11600 23215
rect 11315 23180 11385 23200
rect 11290 23140 11385 23180
rect 11445 23180 11515 23200
rect 11445 23140 11540 23180
rect 11290 23090 11540 23140
rect 11290 23050 11385 23090
rect 11315 23030 11385 23050
rect 11445 23050 11540 23090
rect 11445 23030 11515 23050
rect 11230 23015 11286 23021
rect 11230 22955 11234 23015
rect 11315 23005 11515 23030
rect 11570 23021 11600 23209
rect 11544 23015 11600 23021
rect 11286 22955 11544 22975
rect 11596 22955 11600 23015
rect 11230 22945 11600 22955
rect 11630 23275 12000 23285
rect 11630 23215 11634 23275
rect 11686 23255 11944 23275
rect 11630 23209 11686 23215
rect 11630 23021 11660 23209
rect 11715 23200 11915 23225
rect 11996 23215 12000 23275
rect 11944 23209 12000 23215
rect 11715 23180 11785 23200
rect 11690 23140 11785 23180
rect 11845 23180 11915 23200
rect 11845 23140 11940 23180
rect 11690 23090 11940 23140
rect 11690 23050 11785 23090
rect 11715 23030 11785 23050
rect 11845 23050 11940 23090
rect 11845 23030 11915 23050
rect 11630 23015 11686 23021
rect 11630 22955 11634 23015
rect 11715 23005 11915 23030
rect 11970 23021 12000 23209
rect 11944 23015 12000 23021
rect 11686 22955 11944 22975
rect 11996 22955 12000 23015
rect 11630 22945 12000 22955
rect 12030 23275 12400 23285
rect 12030 23215 12034 23275
rect 12086 23255 12344 23275
rect 12030 23209 12086 23215
rect 12030 23021 12060 23209
rect 12115 23200 12315 23225
rect 12396 23215 12400 23275
rect 12344 23209 12400 23215
rect 12115 23180 12185 23200
rect 12090 23140 12185 23180
rect 12245 23180 12315 23200
rect 12245 23140 12340 23180
rect 12090 23090 12340 23140
rect 12090 23050 12185 23090
rect 12115 23030 12185 23050
rect 12245 23050 12340 23090
rect 12245 23030 12315 23050
rect 12030 23015 12086 23021
rect 12030 22955 12034 23015
rect 12115 23005 12315 23030
rect 12370 23021 12400 23209
rect 12344 23015 12400 23021
rect 12086 22955 12344 22975
rect 12396 22955 12400 23015
rect 12030 22945 12400 22955
rect 12430 23275 12800 23285
rect 12430 23215 12434 23275
rect 12486 23255 12744 23275
rect 12430 23209 12486 23215
rect 12430 23021 12460 23209
rect 12515 23200 12715 23225
rect 12796 23215 12800 23275
rect 12744 23209 12800 23215
rect 12515 23180 12585 23200
rect 12490 23140 12585 23180
rect 12645 23180 12715 23200
rect 12645 23140 12740 23180
rect 12490 23090 12740 23140
rect 12490 23050 12585 23090
rect 12515 23030 12585 23050
rect 12645 23050 12740 23090
rect 12645 23030 12715 23050
rect 12430 23015 12486 23021
rect 12430 22955 12434 23015
rect 12515 23005 12715 23030
rect 12770 23021 12800 23209
rect 12744 23015 12800 23021
rect 12486 22955 12744 22975
rect 12796 22955 12800 23015
rect 12430 22945 12800 22955
rect 12830 23275 13200 23285
rect 12830 23215 12834 23275
rect 12886 23255 13144 23275
rect 12830 23209 12886 23215
rect 12830 23021 12860 23209
rect 12915 23200 13115 23225
rect 13196 23215 13200 23275
rect 13144 23209 13200 23215
rect 12915 23180 12985 23200
rect 12890 23140 12985 23180
rect 13045 23180 13115 23200
rect 13045 23140 13140 23180
rect 12890 23090 13140 23140
rect 12890 23050 12985 23090
rect 12915 23030 12985 23050
rect 13045 23050 13140 23090
rect 13045 23030 13115 23050
rect 12830 23015 12886 23021
rect 12830 22955 12834 23015
rect 12915 23005 13115 23030
rect 13170 23021 13200 23209
rect 13144 23015 13200 23021
rect 12886 22955 13144 22975
rect 13196 22955 13200 23015
rect 12830 22945 13200 22955
rect -370 22905 0 22915
rect -370 22845 -366 22905
rect -314 22885 -56 22905
rect -370 22839 -314 22845
rect -370 22651 -340 22839
rect -285 22830 -85 22855
rect -4 22845 0 22905
rect -56 22839 0 22845
rect -285 22810 -215 22830
rect -310 22770 -215 22810
rect -155 22810 -85 22830
rect -155 22770 -60 22810
rect -310 22720 -60 22770
rect -310 22680 -215 22720
rect -285 22660 -215 22680
rect -155 22680 -60 22720
rect -155 22660 -85 22680
rect -370 22645 -314 22651
rect -370 22585 -366 22645
rect -285 22635 -85 22660
rect -30 22651 0 22839
rect -56 22645 0 22651
rect -314 22585 -56 22605
rect -4 22585 0 22645
rect -370 22575 0 22585
rect 30 22905 400 22915
rect 30 22845 34 22905
rect 86 22885 344 22905
rect 30 22839 86 22845
rect 30 22651 60 22839
rect 115 22830 315 22855
rect 396 22845 400 22905
rect 344 22839 400 22845
rect 115 22810 185 22830
rect 90 22770 185 22810
rect 245 22810 315 22830
rect 245 22770 340 22810
rect 90 22720 340 22770
rect 90 22680 185 22720
rect 115 22660 185 22680
rect 245 22680 340 22720
rect 245 22660 315 22680
rect 30 22645 86 22651
rect 30 22585 34 22645
rect 115 22635 315 22660
rect 370 22651 400 22839
rect 344 22645 400 22651
rect 86 22585 344 22605
rect 396 22585 400 22645
rect 30 22575 400 22585
rect 430 22905 800 22915
rect 430 22845 434 22905
rect 486 22885 744 22905
rect 430 22839 486 22845
rect 430 22651 460 22839
rect 515 22830 715 22855
rect 796 22845 800 22905
rect 744 22839 800 22845
rect 515 22810 585 22830
rect 490 22770 585 22810
rect 645 22810 715 22830
rect 645 22770 740 22810
rect 490 22720 740 22770
rect 490 22680 585 22720
rect 515 22660 585 22680
rect 645 22680 740 22720
rect 645 22660 715 22680
rect 430 22645 486 22651
rect 430 22585 434 22645
rect 515 22635 715 22660
rect 770 22651 800 22839
rect 744 22645 800 22651
rect 486 22585 744 22605
rect 796 22585 800 22645
rect 430 22575 800 22585
rect 830 22905 1200 22915
rect 830 22845 834 22905
rect 886 22885 1144 22905
rect 830 22839 886 22845
rect 830 22651 860 22839
rect 915 22830 1115 22855
rect 1196 22845 1200 22905
rect 1144 22839 1200 22845
rect 915 22810 985 22830
rect 890 22770 985 22810
rect 1045 22810 1115 22830
rect 1045 22770 1140 22810
rect 890 22720 1140 22770
rect 890 22680 985 22720
rect 915 22660 985 22680
rect 1045 22680 1140 22720
rect 1045 22660 1115 22680
rect 830 22645 886 22651
rect 830 22585 834 22645
rect 915 22635 1115 22660
rect 1170 22651 1200 22839
rect 1144 22645 1200 22651
rect 886 22585 1144 22605
rect 1196 22585 1200 22645
rect 830 22575 1200 22585
rect 1230 22905 1600 22915
rect 1230 22845 1234 22905
rect 1286 22885 1544 22905
rect 1230 22839 1286 22845
rect 1230 22651 1260 22839
rect 1315 22830 1515 22855
rect 1596 22845 1600 22905
rect 1544 22839 1600 22845
rect 1315 22810 1385 22830
rect 1290 22770 1385 22810
rect 1445 22810 1515 22830
rect 1445 22770 1540 22810
rect 1290 22720 1540 22770
rect 1290 22680 1385 22720
rect 1315 22660 1385 22680
rect 1445 22680 1540 22720
rect 1445 22660 1515 22680
rect 1230 22645 1286 22651
rect 1230 22585 1234 22645
rect 1315 22635 1515 22660
rect 1570 22651 1600 22839
rect 1544 22645 1600 22651
rect 1286 22585 1544 22605
rect 1596 22585 1600 22645
rect 1230 22575 1600 22585
rect 1630 22905 2000 22915
rect 1630 22845 1634 22905
rect 1686 22885 1944 22905
rect 1630 22839 1686 22845
rect 1630 22651 1660 22839
rect 1715 22830 1915 22855
rect 1996 22845 2000 22905
rect 1944 22839 2000 22845
rect 1715 22810 1785 22830
rect 1690 22770 1785 22810
rect 1845 22810 1915 22830
rect 1845 22770 1940 22810
rect 1690 22720 1940 22770
rect 1690 22680 1785 22720
rect 1715 22660 1785 22680
rect 1845 22680 1940 22720
rect 1845 22660 1915 22680
rect 1630 22645 1686 22651
rect 1630 22585 1634 22645
rect 1715 22635 1915 22660
rect 1970 22651 2000 22839
rect 1944 22645 2000 22651
rect 1686 22585 1944 22605
rect 1996 22585 2000 22645
rect 1630 22575 2000 22585
rect 2030 22905 2400 22915
rect 2030 22845 2034 22905
rect 2086 22885 2344 22905
rect 2030 22839 2086 22845
rect 2030 22651 2060 22839
rect 2115 22830 2315 22855
rect 2396 22845 2400 22905
rect 2344 22839 2400 22845
rect 2115 22810 2185 22830
rect 2090 22770 2185 22810
rect 2245 22810 2315 22830
rect 2245 22770 2340 22810
rect 2090 22720 2340 22770
rect 2090 22680 2185 22720
rect 2115 22660 2185 22680
rect 2245 22680 2340 22720
rect 2245 22660 2315 22680
rect 2030 22645 2086 22651
rect 2030 22585 2034 22645
rect 2115 22635 2315 22660
rect 2370 22651 2400 22839
rect 2344 22645 2400 22651
rect 2086 22585 2344 22605
rect 2396 22585 2400 22645
rect 2030 22575 2400 22585
rect 2430 22905 2800 22915
rect 2430 22845 2434 22905
rect 2486 22885 2744 22905
rect 2430 22839 2486 22845
rect 2430 22651 2460 22839
rect 2515 22830 2715 22855
rect 2796 22845 2800 22905
rect 2744 22839 2800 22845
rect 2515 22810 2585 22830
rect 2490 22770 2585 22810
rect 2645 22810 2715 22830
rect 2645 22770 2740 22810
rect 2490 22720 2740 22770
rect 2490 22680 2585 22720
rect 2515 22660 2585 22680
rect 2645 22680 2740 22720
rect 2645 22660 2715 22680
rect 2430 22645 2486 22651
rect 2430 22585 2434 22645
rect 2515 22635 2715 22660
rect 2770 22651 2800 22839
rect 2744 22645 2800 22651
rect 2486 22585 2744 22605
rect 2796 22585 2800 22645
rect 2430 22575 2800 22585
rect 2830 22905 3200 22915
rect 2830 22845 2834 22905
rect 2886 22885 3144 22905
rect 2830 22839 2886 22845
rect 2830 22651 2860 22839
rect 2915 22830 3115 22855
rect 3196 22845 3200 22905
rect 3144 22839 3200 22845
rect 2915 22810 2985 22830
rect 2890 22770 2985 22810
rect 3045 22810 3115 22830
rect 3045 22770 3140 22810
rect 2890 22720 3140 22770
rect 2890 22680 2985 22720
rect 2915 22660 2985 22680
rect 3045 22680 3140 22720
rect 3045 22660 3115 22680
rect 2830 22645 2886 22651
rect 2830 22585 2834 22645
rect 2915 22635 3115 22660
rect 3170 22651 3200 22839
rect 3144 22645 3200 22651
rect 2886 22585 3144 22605
rect 3196 22585 3200 22645
rect 2830 22575 3200 22585
rect 3230 22905 3600 22915
rect 3230 22845 3234 22905
rect 3286 22885 3544 22905
rect 3230 22839 3286 22845
rect 3230 22651 3260 22839
rect 3315 22830 3515 22855
rect 3596 22845 3600 22905
rect 3544 22839 3600 22845
rect 3315 22810 3385 22830
rect 3290 22770 3385 22810
rect 3445 22810 3515 22830
rect 3445 22770 3540 22810
rect 3290 22720 3540 22770
rect 3290 22680 3385 22720
rect 3315 22660 3385 22680
rect 3445 22680 3540 22720
rect 3445 22660 3515 22680
rect 3230 22645 3286 22651
rect 3230 22585 3234 22645
rect 3315 22635 3515 22660
rect 3570 22651 3600 22839
rect 3544 22645 3600 22651
rect 3286 22585 3544 22605
rect 3596 22585 3600 22645
rect 3230 22575 3600 22585
rect 3630 22905 4000 22915
rect 3630 22845 3634 22905
rect 3686 22885 3944 22905
rect 3630 22839 3686 22845
rect 3630 22651 3660 22839
rect 3715 22830 3915 22855
rect 3996 22845 4000 22905
rect 3944 22839 4000 22845
rect 3715 22810 3785 22830
rect 3690 22770 3785 22810
rect 3845 22810 3915 22830
rect 3845 22770 3940 22810
rect 3690 22720 3940 22770
rect 3690 22680 3785 22720
rect 3715 22660 3785 22680
rect 3845 22680 3940 22720
rect 3845 22660 3915 22680
rect 3630 22645 3686 22651
rect 3630 22585 3634 22645
rect 3715 22635 3915 22660
rect 3970 22651 4000 22839
rect 3944 22645 4000 22651
rect 3686 22585 3944 22605
rect 3996 22585 4000 22645
rect 3630 22575 4000 22585
rect 4030 22905 4400 22915
rect 4030 22845 4034 22905
rect 4086 22885 4344 22905
rect 4030 22839 4086 22845
rect 4030 22651 4060 22839
rect 4115 22830 4315 22855
rect 4396 22845 4400 22905
rect 4344 22839 4400 22845
rect 4115 22810 4185 22830
rect 4090 22770 4185 22810
rect 4245 22810 4315 22830
rect 4245 22770 4340 22810
rect 4090 22720 4340 22770
rect 4090 22680 4185 22720
rect 4115 22660 4185 22680
rect 4245 22680 4340 22720
rect 4245 22660 4315 22680
rect 4030 22645 4086 22651
rect 4030 22585 4034 22645
rect 4115 22635 4315 22660
rect 4370 22651 4400 22839
rect 4344 22645 4400 22651
rect 4086 22585 4344 22605
rect 4396 22585 4400 22645
rect 4030 22575 4400 22585
rect 4430 22905 4800 22915
rect 4430 22845 4434 22905
rect 4486 22885 4744 22905
rect 4430 22839 4486 22845
rect 4430 22651 4460 22839
rect 4515 22830 4715 22855
rect 4796 22845 4800 22905
rect 4744 22839 4800 22845
rect 4515 22810 4585 22830
rect 4490 22770 4585 22810
rect 4645 22810 4715 22830
rect 4645 22770 4740 22810
rect 4490 22720 4740 22770
rect 4490 22680 4585 22720
rect 4515 22660 4585 22680
rect 4645 22680 4740 22720
rect 4645 22660 4715 22680
rect 4430 22645 4486 22651
rect 4430 22585 4434 22645
rect 4515 22635 4715 22660
rect 4770 22651 4800 22839
rect 4744 22645 4800 22651
rect 4486 22585 4744 22605
rect 4796 22585 4800 22645
rect 4430 22575 4800 22585
rect 4830 22905 5200 22915
rect 4830 22845 4834 22905
rect 4886 22885 5144 22905
rect 4830 22839 4886 22845
rect 4830 22651 4860 22839
rect 4915 22830 5115 22855
rect 5196 22845 5200 22905
rect 5144 22839 5200 22845
rect 4915 22810 4985 22830
rect 4890 22770 4985 22810
rect 5045 22810 5115 22830
rect 5045 22770 5140 22810
rect 4890 22720 5140 22770
rect 4890 22680 4985 22720
rect 4915 22660 4985 22680
rect 5045 22680 5140 22720
rect 5045 22660 5115 22680
rect 4830 22645 4886 22651
rect 4830 22585 4834 22645
rect 4915 22635 5115 22660
rect 5170 22651 5200 22839
rect 5144 22645 5200 22651
rect 4886 22585 5144 22605
rect 5196 22585 5200 22645
rect 4830 22575 5200 22585
rect 5230 22905 5600 22915
rect 5230 22845 5234 22905
rect 5286 22885 5544 22905
rect 5230 22839 5286 22845
rect 5230 22651 5260 22839
rect 5315 22830 5515 22855
rect 5596 22845 5600 22905
rect 5544 22839 5600 22845
rect 5315 22810 5385 22830
rect 5290 22770 5385 22810
rect 5445 22810 5515 22830
rect 5445 22770 5540 22810
rect 5290 22720 5540 22770
rect 5290 22680 5385 22720
rect 5315 22660 5385 22680
rect 5445 22680 5540 22720
rect 5445 22660 5515 22680
rect 5230 22645 5286 22651
rect 5230 22585 5234 22645
rect 5315 22635 5515 22660
rect 5570 22651 5600 22839
rect 5544 22645 5600 22651
rect 5286 22585 5544 22605
rect 5596 22585 5600 22645
rect 5230 22575 5600 22585
rect 5630 22905 6000 22915
rect 5630 22845 5634 22905
rect 5686 22885 5944 22905
rect 5630 22839 5686 22845
rect 5630 22651 5660 22839
rect 5715 22830 5915 22855
rect 5996 22845 6000 22905
rect 5944 22839 6000 22845
rect 5715 22810 5785 22830
rect 5690 22770 5785 22810
rect 5845 22810 5915 22830
rect 5845 22770 5940 22810
rect 5690 22720 5940 22770
rect 5690 22680 5785 22720
rect 5715 22660 5785 22680
rect 5845 22680 5940 22720
rect 5845 22660 5915 22680
rect 5630 22645 5686 22651
rect 5630 22585 5634 22645
rect 5715 22635 5915 22660
rect 5970 22651 6000 22839
rect 5944 22645 6000 22651
rect 5686 22585 5944 22605
rect 5996 22585 6000 22645
rect 5630 22575 6000 22585
rect 6030 22905 6400 22915
rect 6030 22845 6034 22905
rect 6086 22885 6344 22905
rect 6030 22839 6086 22845
rect 6030 22651 6060 22839
rect 6115 22830 6315 22855
rect 6396 22845 6400 22905
rect 6344 22839 6400 22845
rect 6115 22810 6185 22830
rect 6090 22770 6185 22810
rect 6245 22810 6315 22830
rect 6245 22770 6340 22810
rect 6090 22720 6340 22770
rect 6090 22680 6185 22720
rect 6115 22660 6185 22680
rect 6245 22680 6340 22720
rect 6245 22660 6315 22680
rect 6030 22645 6086 22651
rect 6030 22585 6034 22645
rect 6115 22635 6315 22660
rect 6370 22651 6400 22839
rect 6344 22645 6400 22651
rect 6086 22585 6344 22605
rect 6396 22585 6400 22645
rect 6030 22575 6400 22585
rect 6430 22905 6800 22915
rect 6430 22845 6434 22905
rect 6486 22885 6744 22905
rect 6430 22839 6486 22845
rect 6430 22651 6460 22839
rect 6515 22830 6715 22855
rect 6796 22845 6800 22905
rect 6744 22839 6800 22845
rect 6515 22810 6585 22830
rect 6490 22770 6585 22810
rect 6645 22810 6715 22830
rect 6645 22770 6740 22810
rect 6490 22720 6740 22770
rect 6490 22680 6585 22720
rect 6515 22660 6585 22680
rect 6645 22680 6740 22720
rect 6645 22660 6715 22680
rect 6430 22645 6486 22651
rect 6430 22585 6434 22645
rect 6515 22635 6715 22660
rect 6770 22651 6800 22839
rect 6744 22645 6800 22651
rect 6486 22585 6744 22605
rect 6796 22585 6800 22645
rect 6430 22575 6800 22585
rect 6830 22905 7200 22915
rect 6830 22845 6834 22905
rect 6886 22885 7144 22905
rect 6830 22839 6886 22845
rect 6830 22651 6860 22839
rect 6915 22830 7115 22855
rect 7196 22845 7200 22905
rect 7144 22839 7200 22845
rect 6915 22810 6985 22830
rect 6890 22770 6985 22810
rect 7045 22810 7115 22830
rect 7045 22770 7140 22810
rect 6890 22720 7140 22770
rect 6890 22680 6985 22720
rect 6915 22660 6985 22680
rect 7045 22680 7140 22720
rect 7045 22660 7115 22680
rect 6830 22645 6886 22651
rect 6830 22585 6834 22645
rect 6915 22635 7115 22660
rect 7170 22651 7200 22839
rect 7144 22645 7200 22651
rect 6886 22585 7144 22605
rect 7196 22585 7200 22645
rect 6830 22575 7200 22585
rect 7230 22905 7600 22915
rect 7230 22845 7234 22905
rect 7286 22885 7544 22905
rect 7230 22839 7286 22845
rect 7230 22651 7260 22839
rect 7315 22830 7515 22855
rect 7596 22845 7600 22905
rect 7544 22839 7600 22845
rect 7315 22810 7385 22830
rect 7290 22770 7385 22810
rect 7445 22810 7515 22830
rect 7445 22770 7540 22810
rect 7290 22720 7540 22770
rect 7290 22680 7385 22720
rect 7315 22660 7385 22680
rect 7445 22680 7540 22720
rect 7445 22660 7515 22680
rect 7230 22645 7286 22651
rect 7230 22585 7234 22645
rect 7315 22635 7515 22660
rect 7570 22651 7600 22839
rect 7544 22645 7600 22651
rect 7286 22585 7544 22605
rect 7596 22585 7600 22645
rect 7230 22575 7600 22585
rect 7630 22905 8000 22915
rect 7630 22845 7634 22905
rect 7686 22885 7944 22905
rect 7630 22839 7686 22845
rect 7630 22651 7660 22839
rect 7715 22830 7915 22855
rect 7996 22845 8000 22905
rect 7944 22839 8000 22845
rect 7715 22810 7785 22830
rect 7690 22770 7785 22810
rect 7845 22810 7915 22830
rect 7845 22770 7940 22810
rect 7690 22720 7940 22770
rect 7690 22680 7785 22720
rect 7715 22660 7785 22680
rect 7845 22680 7940 22720
rect 7845 22660 7915 22680
rect 7630 22645 7686 22651
rect 7630 22585 7634 22645
rect 7715 22635 7915 22660
rect 7970 22651 8000 22839
rect 7944 22645 8000 22651
rect 7686 22585 7944 22605
rect 7996 22585 8000 22645
rect 7630 22575 8000 22585
rect 8030 22905 8400 22915
rect 8030 22845 8034 22905
rect 8086 22885 8344 22905
rect 8030 22839 8086 22845
rect 8030 22651 8060 22839
rect 8115 22830 8315 22855
rect 8396 22845 8400 22905
rect 8344 22839 8400 22845
rect 8115 22810 8185 22830
rect 8090 22770 8185 22810
rect 8245 22810 8315 22830
rect 8245 22770 8340 22810
rect 8090 22720 8340 22770
rect 8090 22680 8185 22720
rect 8115 22660 8185 22680
rect 8245 22680 8340 22720
rect 8245 22660 8315 22680
rect 8030 22645 8086 22651
rect 8030 22585 8034 22645
rect 8115 22635 8315 22660
rect 8370 22651 8400 22839
rect 8344 22645 8400 22651
rect 8086 22585 8344 22605
rect 8396 22585 8400 22645
rect 8030 22575 8400 22585
rect 8430 22905 8800 22915
rect 8430 22845 8434 22905
rect 8486 22885 8744 22905
rect 8430 22839 8486 22845
rect 8430 22651 8460 22839
rect 8515 22830 8715 22855
rect 8796 22845 8800 22905
rect 8744 22839 8800 22845
rect 8515 22810 8585 22830
rect 8490 22770 8585 22810
rect 8645 22810 8715 22830
rect 8645 22770 8740 22810
rect 8490 22720 8740 22770
rect 8490 22680 8585 22720
rect 8515 22660 8585 22680
rect 8645 22680 8740 22720
rect 8645 22660 8715 22680
rect 8430 22645 8486 22651
rect 8430 22585 8434 22645
rect 8515 22635 8715 22660
rect 8770 22651 8800 22839
rect 8744 22645 8800 22651
rect 8486 22585 8744 22605
rect 8796 22585 8800 22645
rect 8430 22575 8800 22585
rect 8830 22905 9200 22915
rect 8830 22845 8834 22905
rect 8886 22885 9144 22905
rect 8830 22839 8886 22845
rect 8830 22651 8860 22839
rect 8915 22830 9115 22855
rect 9196 22845 9200 22905
rect 9144 22839 9200 22845
rect 8915 22810 8985 22830
rect 8890 22770 8985 22810
rect 9045 22810 9115 22830
rect 9045 22770 9140 22810
rect 8890 22720 9140 22770
rect 8890 22680 8985 22720
rect 8915 22660 8985 22680
rect 9045 22680 9140 22720
rect 9045 22660 9115 22680
rect 8830 22645 8886 22651
rect 8830 22585 8834 22645
rect 8915 22635 9115 22660
rect 9170 22651 9200 22839
rect 9144 22645 9200 22651
rect 8886 22585 9144 22605
rect 9196 22585 9200 22645
rect 8830 22575 9200 22585
rect 9230 22905 9600 22915
rect 9230 22845 9234 22905
rect 9286 22885 9544 22905
rect 9230 22839 9286 22845
rect 9230 22651 9260 22839
rect 9315 22830 9515 22855
rect 9596 22845 9600 22905
rect 9544 22839 9600 22845
rect 9315 22810 9385 22830
rect 9290 22770 9385 22810
rect 9445 22810 9515 22830
rect 9445 22770 9540 22810
rect 9290 22720 9540 22770
rect 9290 22680 9385 22720
rect 9315 22660 9385 22680
rect 9445 22680 9540 22720
rect 9445 22660 9515 22680
rect 9230 22645 9286 22651
rect 9230 22585 9234 22645
rect 9315 22635 9515 22660
rect 9570 22651 9600 22839
rect 9544 22645 9600 22651
rect 9286 22585 9544 22605
rect 9596 22585 9600 22645
rect 9230 22575 9600 22585
rect 9630 22905 10000 22915
rect 9630 22845 9634 22905
rect 9686 22885 9944 22905
rect 9630 22839 9686 22845
rect 9630 22651 9660 22839
rect 9715 22830 9915 22855
rect 9996 22845 10000 22905
rect 9944 22839 10000 22845
rect 9715 22810 9785 22830
rect 9690 22770 9785 22810
rect 9845 22810 9915 22830
rect 9845 22770 9940 22810
rect 9690 22720 9940 22770
rect 9690 22680 9785 22720
rect 9715 22660 9785 22680
rect 9845 22680 9940 22720
rect 9845 22660 9915 22680
rect 9630 22645 9686 22651
rect 9630 22585 9634 22645
rect 9715 22635 9915 22660
rect 9970 22651 10000 22839
rect 9944 22645 10000 22651
rect 9686 22585 9944 22605
rect 9996 22585 10000 22645
rect 9630 22575 10000 22585
rect 10030 22905 10400 22915
rect 10030 22845 10034 22905
rect 10086 22885 10344 22905
rect 10030 22839 10086 22845
rect 10030 22651 10060 22839
rect 10115 22830 10315 22855
rect 10396 22845 10400 22905
rect 10344 22839 10400 22845
rect 10115 22810 10185 22830
rect 10090 22770 10185 22810
rect 10245 22810 10315 22830
rect 10245 22770 10340 22810
rect 10090 22720 10340 22770
rect 10090 22680 10185 22720
rect 10115 22660 10185 22680
rect 10245 22680 10340 22720
rect 10245 22660 10315 22680
rect 10030 22645 10086 22651
rect 10030 22585 10034 22645
rect 10115 22635 10315 22660
rect 10370 22651 10400 22839
rect 10344 22645 10400 22651
rect 10086 22585 10344 22605
rect 10396 22585 10400 22645
rect 10030 22575 10400 22585
rect 10430 22905 10800 22915
rect 10430 22845 10434 22905
rect 10486 22885 10744 22905
rect 10430 22839 10486 22845
rect 10430 22651 10460 22839
rect 10515 22830 10715 22855
rect 10796 22845 10800 22905
rect 10744 22839 10800 22845
rect 10515 22810 10585 22830
rect 10490 22770 10585 22810
rect 10645 22810 10715 22830
rect 10645 22770 10740 22810
rect 10490 22720 10740 22770
rect 10490 22680 10585 22720
rect 10515 22660 10585 22680
rect 10645 22680 10740 22720
rect 10645 22660 10715 22680
rect 10430 22645 10486 22651
rect 10430 22585 10434 22645
rect 10515 22635 10715 22660
rect 10770 22651 10800 22839
rect 10744 22645 10800 22651
rect 10486 22585 10744 22605
rect 10796 22585 10800 22645
rect 10430 22575 10800 22585
rect 10830 22905 11200 22915
rect 10830 22845 10834 22905
rect 10886 22885 11144 22905
rect 10830 22839 10886 22845
rect 10830 22651 10860 22839
rect 10915 22830 11115 22855
rect 11196 22845 11200 22905
rect 11144 22839 11200 22845
rect 10915 22810 10985 22830
rect 10890 22770 10985 22810
rect 11045 22810 11115 22830
rect 11045 22770 11140 22810
rect 10890 22720 11140 22770
rect 10890 22680 10985 22720
rect 10915 22660 10985 22680
rect 11045 22680 11140 22720
rect 11045 22660 11115 22680
rect 10830 22645 10886 22651
rect 10830 22585 10834 22645
rect 10915 22635 11115 22660
rect 11170 22651 11200 22839
rect 11144 22645 11200 22651
rect 10886 22585 11144 22605
rect 11196 22585 11200 22645
rect 10830 22575 11200 22585
rect 11230 22905 11600 22915
rect 11230 22845 11234 22905
rect 11286 22885 11544 22905
rect 11230 22839 11286 22845
rect 11230 22651 11260 22839
rect 11315 22830 11515 22855
rect 11596 22845 11600 22905
rect 11544 22839 11600 22845
rect 11315 22810 11385 22830
rect 11290 22770 11385 22810
rect 11445 22810 11515 22830
rect 11445 22770 11540 22810
rect 11290 22720 11540 22770
rect 11290 22680 11385 22720
rect 11315 22660 11385 22680
rect 11445 22680 11540 22720
rect 11445 22660 11515 22680
rect 11230 22645 11286 22651
rect 11230 22585 11234 22645
rect 11315 22635 11515 22660
rect 11570 22651 11600 22839
rect 11544 22645 11600 22651
rect 11286 22585 11544 22605
rect 11596 22585 11600 22645
rect 11230 22575 11600 22585
rect 11630 22905 12000 22915
rect 11630 22845 11634 22905
rect 11686 22885 11944 22905
rect 11630 22839 11686 22845
rect 11630 22651 11660 22839
rect 11715 22830 11915 22855
rect 11996 22845 12000 22905
rect 11944 22839 12000 22845
rect 11715 22810 11785 22830
rect 11690 22770 11785 22810
rect 11845 22810 11915 22830
rect 11845 22770 11940 22810
rect 11690 22720 11940 22770
rect 11690 22680 11785 22720
rect 11715 22660 11785 22680
rect 11845 22680 11940 22720
rect 11845 22660 11915 22680
rect 11630 22645 11686 22651
rect 11630 22585 11634 22645
rect 11715 22635 11915 22660
rect 11970 22651 12000 22839
rect 11944 22645 12000 22651
rect 11686 22585 11944 22605
rect 11996 22585 12000 22645
rect 11630 22575 12000 22585
rect 12030 22905 12400 22915
rect 12030 22845 12034 22905
rect 12086 22885 12344 22905
rect 12030 22839 12086 22845
rect 12030 22651 12060 22839
rect 12115 22830 12315 22855
rect 12396 22845 12400 22905
rect 12344 22839 12400 22845
rect 12115 22810 12185 22830
rect 12090 22770 12185 22810
rect 12245 22810 12315 22830
rect 12245 22770 12340 22810
rect 12090 22720 12340 22770
rect 12090 22680 12185 22720
rect 12115 22660 12185 22680
rect 12245 22680 12340 22720
rect 12245 22660 12315 22680
rect 12030 22645 12086 22651
rect 12030 22585 12034 22645
rect 12115 22635 12315 22660
rect 12370 22651 12400 22839
rect 12344 22645 12400 22651
rect 12086 22585 12344 22605
rect 12396 22585 12400 22645
rect 12030 22575 12400 22585
rect 12430 22905 12800 22915
rect 12430 22845 12434 22905
rect 12486 22885 12744 22905
rect 12430 22839 12486 22845
rect 12430 22651 12460 22839
rect 12515 22830 12715 22855
rect 12796 22845 12800 22905
rect 12744 22839 12800 22845
rect 12515 22810 12585 22830
rect 12490 22770 12585 22810
rect 12645 22810 12715 22830
rect 12645 22770 12740 22810
rect 12490 22720 12740 22770
rect 12490 22680 12585 22720
rect 12515 22660 12585 22680
rect 12645 22680 12740 22720
rect 12645 22660 12715 22680
rect 12430 22645 12486 22651
rect 12430 22585 12434 22645
rect 12515 22635 12715 22660
rect 12770 22651 12800 22839
rect 12744 22645 12800 22651
rect 12486 22585 12744 22605
rect 12796 22585 12800 22645
rect 12430 22575 12800 22585
rect 12830 22905 13200 22915
rect 12830 22845 12834 22905
rect 12886 22885 13144 22905
rect 12830 22839 12886 22845
rect 12830 22651 12860 22839
rect 12915 22830 13115 22855
rect 13196 22845 13200 22905
rect 13144 22839 13200 22845
rect 12915 22810 12985 22830
rect 12890 22770 12985 22810
rect 13045 22810 13115 22830
rect 13045 22770 13140 22810
rect 12890 22720 13140 22770
rect 12890 22680 12985 22720
rect 12915 22660 12985 22680
rect 13045 22680 13140 22720
rect 13045 22660 13115 22680
rect 12830 22645 12886 22651
rect 12830 22585 12834 22645
rect 12915 22635 13115 22660
rect 13170 22651 13200 22839
rect 13144 22645 13200 22651
rect 12886 22585 13144 22605
rect 13196 22585 13200 22645
rect 12830 22575 13200 22585
rect -370 22535 0 22545
rect -370 22475 -366 22535
rect -314 22515 -56 22535
rect -370 22469 -314 22475
rect -370 22281 -340 22469
rect -285 22460 -85 22485
rect -4 22475 0 22535
rect -56 22469 0 22475
rect -285 22440 -215 22460
rect -310 22400 -215 22440
rect -155 22440 -85 22460
rect -155 22400 -60 22440
rect -310 22350 -60 22400
rect -310 22310 -215 22350
rect -285 22290 -215 22310
rect -155 22310 -60 22350
rect -155 22290 -85 22310
rect -370 22275 -314 22281
rect -370 22215 -366 22275
rect -285 22265 -85 22290
rect -30 22281 0 22469
rect -56 22275 0 22281
rect -314 22215 -56 22235
rect -4 22215 0 22275
rect -370 22205 0 22215
rect 30 22535 400 22545
rect 30 22475 34 22535
rect 86 22515 344 22535
rect 30 22469 86 22475
rect 30 22281 60 22469
rect 115 22460 315 22485
rect 396 22475 400 22535
rect 344 22469 400 22475
rect 115 22440 185 22460
rect 90 22400 185 22440
rect 245 22440 315 22460
rect 245 22400 340 22440
rect 90 22350 340 22400
rect 90 22310 185 22350
rect 115 22290 185 22310
rect 245 22310 340 22350
rect 245 22290 315 22310
rect 30 22275 86 22281
rect 30 22215 34 22275
rect 115 22265 315 22290
rect 370 22281 400 22469
rect 344 22275 400 22281
rect 86 22215 344 22235
rect 396 22215 400 22275
rect 30 22205 400 22215
rect 430 22535 800 22545
rect 430 22475 434 22535
rect 486 22515 744 22535
rect 430 22469 486 22475
rect 430 22281 460 22469
rect 515 22460 715 22485
rect 796 22475 800 22535
rect 744 22469 800 22475
rect 515 22440 585 22460
rect 490 22400 585 22440
rect 645 22440 715 22460
rect 645 22400 740 22440
rect 490 22350 740 22400
rect 490 22310 585 22350
rect 515 22290 585 22310
rect 645 22310 740 22350
rect 645 22290 715 22310
rect 430 22275 486 22281
rect 430 22215 434 22275
rect 515 22265 715 22290
rect 770 22281 800 22469
rect 744 22275 800 22281
rect 486 22215 744 22235
rect 796 22215 800 22275
rect 430 22205 800 22215
rect 830 22535 1200 22545
rect 830 22475 834 22535
rect 886 22515 1144 22535
rect 830 22469 886 22475
rect 830 22281 860 22469
rect 915 22460 1115 22485
rect 1196 22475 1200 22535
rect 1144 22469 1200 22475
rect 915 22440 985 22460
rect 890 22400 985 22440
rect 1045 22440 1115 22460
rect 1045 22400 1140 22440
rect 890 22350 1140 22400
rect 890 22310 985 22350
rect 915 22290 985 22310
rect 1045 22310 1140 22350
rect 1045 22290 1115 22310
rect 830 22275 886 22281
rect 830 22215 834 22275
rect 915 22265 1115 22290
rect 1170 22281 1200 22469
rect 1144 22275 1200 22281
rect 886 22215 1144 22235
rect 1196 22215 1200 22275
rect 830 22205 1200 22215
rect 1230 22535 1600 22545
rect 1230 22475 1234 22535
rect 1286 22515 1544 22535
rect 1230 22469 1286 22475
rect 1230 22281 1260 22469
rect 1315 22460 1515 22485
rect 1596 22475 1600 22535
rect 1544 22469 1600 22475
rect 1315 22440 1385 22460
rect 1290 22400 1385 22440
rect 1445 22440 1515 22460
rect 1445 22400 1540 22440
rect 1290 22350 1540 22400
rect 1290 22310 1385 22350
rect 1315 22290 1385 22310
rect 1445 22310 1540 22350
rect 1445 22290 1515 22310
rect 1230 22275 1286 22281
rect 1230 22215 1234 22275
rect 1315 22265 1515 22290
rect 1570 22281 1600 22469
rect 1544 22275 1600 22281
rect 1286 22215 1544 22235
rect 1596 22215 1600 22275
rect 1230 22205 1600 22215
rect 1630 22535 2000 22545
rect 1630 22475 1634 22535
rect 1686 22515 1944 22535
rect 1630 22469 1686 22475
rect 1630 22281 1660 22469
rect 1715 22460 1915 22485
rect 1996 22475 2000 22535
rect 1944 22469 2000 22475
rect 1715 22440 1785 22460
rect 1690 22400 1785 22440
rect 1845 22440 1915 22460
rect 1845 22400 1940 22440
rect 1690 22350 1940 22400
rect 1690 22310 1785 22350
rect 1715 22290 1785 22310
rect 1845 22310 1940 22350
rect 1845 22290 1915 22310
rect 1630 22275 1686 22281
rect 1630 22215 1634 22275
rect 1715 22265 1915 22290
rect 1970 22281 2000 22469
rect 1944 22275 2000 22281
rect 1686 22215 1944 22235
rect 1996 22215 2000 22275
rect 1630 22205 2000 22215
rect 2030 22535 2400 22545
rect 2030 22475 2034 22535
rect 2086 22515 2344 22535
rect 2030 22469 2086 22475
rect 2030 22281 2060 22469
rect 2115 22460 2315 22485
rect 2396 22475 2400 22535
rect 2344 22469 2400 22475
rect 2115 22440 2185 22460
rect 2090 22400 2185 22440
rect 2245 22440 2315 22460
rect 2245 22400 2340 22440
rect 2090 22350 2340 22400
rect 2090 22310 2185 22350
rect 2115 22290 2185 22310
rect 2245 22310 2340 22350
rect 2245 22290 2315 22310
rect 2030 22275 2086 22281
rect 2030 22215 2034 22275
rect 2115 22265 2315 22290
rect 2370 22281 2400 22469
rect 2344 22275 2400 22281
rect 2086 22215 2344 22235
rect 2396 22215 2400 22275
rect 2030 22205 2400 22215
rect 2430 22535 2800 22545
rect 2430 22475 2434 22535
rect 2486 22515 2744 22535
rect 2430 22469 2486 22475
rect 2430 22281 2460 22469
rect 2515 22460 2715 22485
rect 2796 22475 2800 22535
rect 2744 22469 2800 22475
rect 2515 22440 2585 22460
rect 2490 22400 2585 22440
rect 2645 22440 2715 22460
rect 2645 22400 2740 22440
rect 2490 22350 2740 22400
rect 2490 22310 2585 22350
rect 2515 22290 2585 22310
rect 2645 22310 2740 22350
rect 2645 22290 2715 22310
rect 2430 22275 2486 22281
rect 2430 22215 2434 22275
rect 2515 22265 2715 22290
rect 2770 22281 2800 22469
rect 2744 22275 2800 22281
rect 2486 22215 2744 22235
rect 2796 22215 2800 22275
rect 2430 22205 2800 22215
rect 2830 22535 3200 22545
rect 2830 22475 2834 22535
rect 2886 22515 3144 22535
rect 2830 22469 2886 22475
rect 2830 22281 2860 22469
rect 2915 22460 3115 22485
rect 3196 22475 3200 22535
rect 3144 22469 3200 22475
rect 2915 22440 2985 22460
rect 2890 22400 2985 22440
rect 3045 22440 3115 22460
rect 3045 22400 3140 22440
rect 2890 22350 3140 22400
rect 2890 22310 2985 22350
rect 2915 22290 2985 22310
rect 3045 22310 3140 22350
rect 3045 22290 3115 22310
rect 2830 22275 2886 22281
rect 2830 22215 2834 22275
rect 2915 22265 3115 22290
rect 3170 22281 3200 22469
rect 3144 22275 3200 22281
rect 2886 22215 3144 22235
rect 3196 22215 3200 22275
rect 2830 22205 3200 22215
rect 3230 22535 3600 22545
rect 3230 22475 3234 22535
rect 3286 22515 3544 22535
rect 3230 22469 3286 22475
rect 3230 22281 3260 22469
rect 3315 22460 3515 22485
rect 3596 22475 3600 22535
rect 3544 22469 3600 22475
rect 3315 22440 3385 22460
rect 3290 22400 3385 22440
rect 3445 22440 3515 22460
rect 3445 22400 3540 22440
rect 3290 22350 3540 22400
rect 3290 22310 3385 22350
rect 3315 22290 3385 22310
rect 3445 22310 3540 22350
rect 3445 22290 3515 22310
rect 3230 22275 3286 22281
rect 3230 22215 3234 22275
rect 3315 22265 3515 22290
rect 3570 22281 3600 22469
rect 3544 22275 3600 22281
rect 3286 22215 3544 22235
rect 3596 22215 3600 22275
rect 3230 22205 3600 22215
rect 3630 22535 4000 22545
rect 3630 22475 3634 22535
rect 3686 22515 3944 22535
rect 3630 22469 3686 22475
rect 3630 22281 3660 22469
rect 3715 22460 3915 22485
rect 3996 22475 4000 22535
rect 3944 22469 4000 22475
rect 3715 22440 3785 22460
rect 3690 22400 3785 22440
rect 3845 22440 3915 22460
rect 3845 22400 3940 22440
rect 3690 22350 3940 22400
rect 3690 22310 3785 22350
rect 3715 22290 3785 22310
rect 3845 22310 3940 22350
rect 3845 22290 3915 22310
rect 3630 22275 3686 22281
rect 3630 22215 3634 22275
rect 3715 22265 3915 22290
rect 3970 22281 4000 22469
rect 3944 22275 4000 22281
rect 3686 22215 3944 22235
rect 3996 22215 4000 22275
rect 3630 22205 4000 22215
rect 4030 22535 4400 22545
rect 4030 22475 4034 22535
rect 4086 22515 4344 22535
rect 4030 22469 4086 22475
rect 4030 22281 4060 22469
rect 4115 22460 4315 22485
rect 4396 22475 4400 22535
rect 4344 22469 4400 22475
rect 4115 22440 4185 22460
rect 4090 22400 4185 22440
rect 4245 22440 4315 22460
rect 4245 22400 4340 22440
rect 4090 22350 4340 22400
rect 4090 22310 4185 22350
rect 4115 22290 4185 22310
rect 4245 22310 4340 22350
rect 4245 22290 4315 22310
rect 4030 22275 4086 22281
rect 4030 22215 4034 22275
rect 4115 22265 4315 22290
rect 4370 22281 4400 22469
rect 4344 22275 4400 22281
rect 4086 22215 4344 22235
rect 4396 22215 4400 22275
rect 4030 22205 4400 22215
rect 4430 22535 4800 22545
rect 4430 22475 4434 22535
rect 4486 22515 4744 22535
rect 4430 22469 4486 22475
rect 4430 22281 4460 22469
rect 4515 22460 4715 22485
rect 4796 22475 4800 22535
rect 4744 22469 4800 22475
rect 4515 22440 4585 22460
rect 4490 22400 4585 22440
rect 4645 22440 4715 22460
rect 4645 22400 4740 22440
rect 4490 22350 4740 22400
rect 4490 22310 4585 22350
rect 4515 22290 4585 22310
rect 4645 22310 4740 22350
rect 4645 22290 4715 22310
rect 4430 22275 4486 22281
rect 4430 22215 4434 22275
rect 4515 22265 4715 22290
rect 4770 22281 4800 22469
rect 4744 22275 4800 22281
rect 4486 22215 4744 22235
rect 4796 22215 4800 22275
rect 4430 22205 4800 22215
rect 4830 22535 5200 22545
rect 4830 22475 4834 22535
rect 4886 22515 5144 22535
rect 4830 22469 4886 22475
rect 4830 22281 4860 22469
rect 4915 22460 5115 22485
rect 5196 22475 5200 22535
rect 5144 22469 5200 22475
rect 4915 22440 4985 22460
rect 4890 22400 4985 22440
rect 5045 22440 5115 22460
rect 5045 22400 5140 22440
rect 4890 22350 5140 22400
rect 4890 22310 4985 22350
rect 4915 22290 4985 22310
rect 5045 22310 5140 22350
rect 5045 22290 5115 22310
rect 4830 22275 4886 22281
rect 4830 22215 4834 22275
rect 4915 22265 5115 22290
rect 5170 22281 5200 22469
rect 5144 22275 5200 22281
rect 4886 22215 5144 22235
rect 5196 22215 5200 22275
rect 4830 22205 5200 22215
rect 5230 22535 5600 22545
rect 5230 22475 5234 22535
rect 5286 22515 5544 22535
rect 5230 22469 5286 22475
rect 5230 22281 5260 22469
rect 5315 22460 5515 22485
rect 5596 22475 5600 22535
rect 5544 22469 5600 22475
rect 5315 22440 5385 22460
rect 5290 22400 5385 22440
rect 5445 22440 5515 22460
rect 5445 22400 5540 22440
rect 5290 22350 5540 22400
rect 5290 22310 5385 22350
rect 5315 22290 5385 22310
rect 5445 22310 5540 22350
rect 5445 22290 5515 22310
rect 5230 22275 5286 22281
rect 5230 22215 5234 22275
rect 5315 22265 5515 22290
rect 5570 22281 5600 22469
rect 5544 22275 5600 22281
rect 5286 22215 5544 22235
rect 5596 22215 5600 22275
rect 5230 22205 5600 22215
rect 5630 22535 6000 22545
rect 5630 22475 5634 22535
rect 5686 22515 5944 22535
rect 5630 22469 5686 22475
rect 5630 22281 5660 22469
rect 5715 22460 5915 22485
rect 5996 22475 6000 22535
rect 5944 22469 6000 22475
rect 5715 22440 5785 22460
rect 5690 22400 5785 22440
rect 5845 22440 5915 22460
rect 5845 22400 5940 22440
rect 5690 22350 5940 22400
rect 5690 22310 5785 22350
rect 5715 22290 5785 22310
rect 5845 22310 5940 22350
rect 5845 22290 5915 22310
rect 5630 22275 5686 22281
rect 5630 22215 5634 22275
rect 5715 22265 5915 22290
rect 5970 22281 6000 22469
rect 5944 22275 6000 22281
rect 5686 22215 5944 22235
rect 5996 22215 6000 22275
rect 5630 22205 6000 22215
rect 6030 22535 6400 22545
rect 6030 22475 6034 22535
rect 6086 22515 6344 22535
rect 6030 22469 6086 22475
rect 6030 22281 6060 22469
rect 6115 22460 6315 22485
rect 6396 22475 6400 22535
rect 6344 22469 6400 22475
rect 6115 22440 6185 22460
rect 6090 22400 6185 22440
rect 6245 22440 6315 22460
rect 6245 22400 6340 22440
rect 6090 22350 6340 22400
rect 6090 22310 6185 22350
rect 6115 22290 6185 22310
rect 6245 22310 6340 22350
rect 6245 22290 6315 22310
rect 6030 22275 6086 22281
rect 6030 22215 6034 22275
rect 6115 22265 6315 22290
rect 6370 22281 6400 22469
rect 6344 22275 6400 22281
rect 6086 22215 6344 22235
rect 6396 22215 6400 22275
rect 6030 22205 6400 22215
rect 6430 22535 6800 22545
rect 6430 22475 6434 22535
rect 6486 22515 6744 22535
rect 6430 22469 6486 22475
rect 6430 22281 6460 22469
rect 6515 22460 6715 22485
rect 6796 22475 6800 22535
rect 6744 22469 6800 22475
rect 6515 22440 6585 22460
rect 6490 22400 6585 22440
rect 6645 22440 6715 22460
rect 6645 22400 6740 22440
rect 6490 22350 6740 22400
rect 6490 22310 6585 22350
rect 6515 22290 6585 22310
rect 6645 22310 6740 22350
rect 6645 22290 6715 22310
rect 6430 22275 6486 22281
rect 6430 22215 6434 22275
rect 6515 22265 6715 22290
rect 6770 22281 6800 22469
rect 6744 22275 6800 22281
rect 6486 22215 6744 22235
rect 6796 22215 6800 22275
rect 6430 22205 6800 22215
rect 6830 22535 7200 22545
rect 6830 22475 6834 22535
rect 6886 22515 7144 22535
rect 6830 22469 6886 22475
rect 6830 22281 6860 22469
rect 6915 22460 7115 22485
rect 7196 22475 7200 22535
rect 7144 22469 7200 22475
rect 6915 22440 6985 22460
rect 6890 22400 6985 22440
rect 7045 22440 7115 22460
rect 7045 22400 7140 22440
rect 6890 22350 7140 22400
rect 6890 22310 6985 22350
rect 6915 22290 6985 22310
rect 7045 22310 7140 22350
rect 7045 22290 7115 22310
rect 6830 22275 6886 22281
rect 6830 22215 6834 22275
rect 6915 22265 7115 22290
rect 7170 22281 7200 22469
rect 7144 22275 7200 22281
rect 6886 22215 7144 22235
rect 7196 22215 7200 22275
rect 6830 22205 7200 22215
rect 7230 22535 7600 22545
rect 7230 22475 7234 22535
rect 7286 22515 7544 22535
rect 7230 22469 7286 22475
rect 7230 22281 7260 22469
rect 7315 22460 7515 22485
rect 7596 22475 7600 22535
rect 7544 22469 7600 22475
rect 7315 22440 7385 22460
rect 7290 22400 7385 22440
rect 7445 22440 7515 22460
rect 7445 22400 7540 22440
rect 7290 22350 7540 22400
rect 7290 22310 7385 22350
rect 7315 22290 7385 22310
rect 7445 22310 7540 22350
rect 7445 22290 7515 22310
rect 7230 22275 7286 22281
rect 7230 22215 7234 22275
rect 7315 22265 7515 22290
rect 7570 22281 7600 22469
rect 7544 22275 7600 22281
rect 7286 22215 7544 22235
rect 7596 22215 7600 22275
rect 7230 22205 7600 22215
rect 7630 22535 8000 22545
rect 7630 22475 7634 22535
rect 7686 22515 7944 22535
rect 7630 22469 7686 22475
rect 7630 22281 7660 22469
rect 7715 22460 7915 22485
rect 7996 22475 8000 22535
rect 7944 22469 8000 22475
rect 7715 22440 7785 22460
rect 7690 22400 7785 22440
rect 7845 22440 7915 22460
rect 7845 22400 7940 22440
rect 7690 22350 7940 22400
rect 7690 22310 7785 22350
rect 7715 22290 7785 22310
rect 7845 22310 7940 22350
rect 7845 22290 7915 22310
rect 7630 22275 7686 22281
rect 7630 22215 7634 22275
rect 7715 22265 7915 22290
rect 7970 22281 8000 22469
rect 7944 22275 8000 22281
rect 7686 22215 7944 22235
rect 7996 22215 8000 22275
rect 7630 22205 8000 22215
rect 8030 22535 8400 22545
rect 8030 22475 8034 22535
rect 8086 22515 8344 22535
rect 8030 22469 8086 22475
rect 8030 22281 8060 22469
rect 8115 22460 8315 22485
rect 8396 22475 8400 22535
rect 8344 22469 8400 22475
rect 8115 22440 8185 22460
rect 8090 22400 8185 22440
rect 8245 22440 8315 22460
rect 8245 22400 8340 22440
rect 8090 22350 8340 22400
rect 8090 22310 8185 22350
rect 8115 22290 8185 22310
rect 8245 22310 8340 22350
rect 8245 22290 8315 22310
rect 8030 22275 8086 22281
rect 8030 22215 8034 22275
rect 8115 22265 8315 22290
rect 8370 22281 8400 22469
rect 8344 22275 8400 22281
rect 8086 22215 8344 22235
rect 8396 22215 8400 22275
rect 8030 22205 8400 22215
rect 8430 22535 8800 22545
rect 8430 22475 8434 22535
rect 8486 22515 8744 22535
rect 8430 22469 8486 22475
rect 8430 22281 8460 22469
rect 8515 22460 8715 22485
rect 8796 22475 8800 22535
rect 8744 22469 8800 22475
rect 8515 22440 8585 22460
rect 8490 22400 8585 22440
rect 8645 22440 8715 22460
rect 8645 22400 8740 22440
rect 8490 22350 8740 22400
rect 8490 22310 8585 22350
rect 8515 22290 8585 22310
rect 8645 22310 8740 22350
rect 8645 22290 8715 22310
rect 8430 22275 8486 22281
rect 8430 22215 8434 22275
rect 8515 22265 8715 22290
rect 8770 22281 8800 22469
rect 8744 22275 8800 22281
rect 8486 22215 8744 22235
rect 8796 22215 8800 22275
rect 8430 22205 8800 22215
rect 8830 22535 9200 22545
rect 8830 22475 8834 22535
rect 8886 22515 9144 22535
rect 8830 22469 8886 22475
rect 8830 22281 8860 22469
rect 8915 22460 9115 22485
rect 9196 22475 9200 22535
rect 9144 22469 9200 22475
rect 8915 22440 8985 22460
rect 8890 22400 8985 22440
rect 9045 22440 9115 22460
rect 9045 22400 9140 22440
rect 8890 22350 9140 22400
rect 8890 22310 8985 22350
rect 8915 22290 8985 22310
rect 9045 22310 9140 22350
rect 9045 22290 9115 22310
rect 8830 22275 8886 22281
rect 8830 22215 8834 22275
rect 8915 22265 9115 22290
rect 9170 22281 9200 22469
rect 9144 22275 9200 22281
rect 8886 22215 9144 22235
rect 9196 22215 9200 22275
rect 8830 22205 9200 22215
rect 9230 22535 9600 22545
rect 9230 22475 9234 22535
rect 9286 22515 9544 22535
rect 9230 22469 9286 22475
rect 9230 22281 9260 22469
rect 9315 22460 9515 22485
rect 9596 22475 9600 22535
rect 9544 22469 9600 22475
rect 9315 22440 9385 22460
rect 9290 22400 9385 22440
rect 9445 22440 9515 22460
rect 9445 22400 9540 22440
rect 9290 22350 9540 22400
rect 9290 22310 9385 22350
rect 9315 22290 9385 22310
rect 9445 22310 9540 22350
rect 9445 22290 9515 22310
rect 9230 22275 9286 22281
rect 9230 22215 9234 22275
rect 9315 22265 9515 22290
rect 9570 22281 9600 22469
rect 9544 22275 9600 22281
rect 9286 22215 9544 22235
rect 9596 22215 9600 22275
rect 9230 22205 9600 22215
rect 9630 22535 10000 22545
rect 9630 22475 9634 22535
rect 9686 22515 9944 22535
rect 9630 22469 9686 22475
rect 9630 22281 9660 22469
rect 9715 22460 9915 22485
rect 9996 22475 10000 22535
rect 9944 22469 10000 22475
rect 9715 22440 9785 22460
rect 9690 22400 9785 22440
rect 9845 22440 9915 22460
rect 9845 22400 9940 22440
rect 9690 22350 9940 22400
rect 9690 22310 9785 22350
rect 9715 22290 9785 22310
rect 9845 22310 9940 22350
rect 9845 22290 9915 22310
rect 9630 22275 9686 22281
rect 9630 22215 9634 22275
rect 9715 22265 9915 22290
rect 9970 22281 10000 22469
rect 9944 22275 10000 22281
rect 9686 22215 9944 22235
rect 9996 22215 10000 22275
rect 9630 22205 10000 22215
rect 10030 22535 10400 22545
rect 10030 22475 10034 22535
rect 10086 22515 10344 22535
rect 10030 22469 10086 22475
rect 10030 22281 10060 22469
rect 10115 22460 10315 22485
rect 10396 22475 10400 22535
rect 10344 22469 10400 22475
rect 10115 22440 10185 22460
rect 10090 22400 10185 22440
rect 10245 22440 10315 22460
rect 10245 22400 10340 22440
rect 10090 22350 10340 22400
rect 10090 22310 10185 22350
rect 10115 22290 10185 22310
rect 10245 22310 10340 22350
rect 10245 22290 10315 22310
rect 10030 22275 10086 22281
rect 10030 22215 10034 22275
rect 10115 22265 10315 22290
rect 10370 22281 10400 22469
rect 10344 22275 10400 22281
rect 10086 22215 10344 22235
rect 10396 22215 10400 22275
rect 10030 22205 10400 22215
rect 10430 22535 10800 22545
rect 10430 22475 10434 22535
rect 10486 22515 10744 22535
rect 10430 22469 10486 22475
rect 10430 22281 10460 22469
rect 10515 22460 10715 22485
rect 10796 22475 10800 22535
rect 10744 22469 10800 22475
rect 10515 22440 10585 22460
rect 10490 22400 10585 22440
rect 10645 22440 10715 22460
rect 10645 22400 10740 22440
rect 10490 22350 10740 22400
rect 10490 22310 10585 22350
rect 10515 22290 10585 22310
rect 10645 22310 10740 22350
rect 10645 22290 10715 22310
rect 10430 22275 10486 22281
rect 10430 22215 10434 22275
rect 10515 22265 10715 22290
rect 10770 22281 10800 22469
rect 10744 22275 10800 22281
rect 10486 22215 10744 22235
rect 10796 22215 10800 22275
rect 10430 22205 10800 22215
rect 10830 22535 11200 22545
rect 10830 22475 10834 22535
rect 10886 22515 11144 22535
rect 10830 22469 10886 22475
rect 10830 22281 10860 22469
rect 10915 22460 11115 22485
rect 11196 22475 11200 22535
rect 11144 22469 11200 22475
rect 10915 22440 10985 22460
rect 10890 22400 10985 22440
rect 11045 22440 11115 22460
rect 11045 22400 11140 22440
rect 10890 22350 11140 22400
rect 10890 22310 10985 22350
rect 10915 22290 10985 22310
rect 11045 22310 11140 22350
rect 11045 22290 11115 22310
rect 10830 22275 10886 22281
rect 10830 22215 10834 22275
rect 10915 22265 11115 22290
rect 11170 22281 11200 22469
rect 11144 22275 11200 22281
rect 10886 22215 11144 22235
rect 11196 22215 11200 22275
rect 10830 22205 11200 22215
rect 11230 22535 11600 22545
rect 11230 22475 11234 22535
rect 11286 22515 11544 22535
rect 11230 22469 11286 22475
rect 11230 22281 11260 22469
rect 11315 22460 11515 22485
rect 11596 22475 11600 22535
rect 11544 22469 11600 22475
rect 11315 22440 11385 22460
rect 11290 22400 11385 22440
rect 11445 22440 11515 22460
rect 11445 22400 11540 22440
rect 11290 22350 11540 22400
rect 11290 22310 11385 22350
rect 11315 22290 11385 22310
rect 11445 22310 11540 22350
rect 11445 22290 11515 22310
rect 11230 22275 11286 22281
rect 11230 22215 11234 22275
rect 11315 22265 11515 22290
rect 11570 22281 11600 22469
rect 11544 22275 11600 22281
rect 11286 22215 11544 22235
rect 11596 22215 11600 22275
rect 11230 22205 11600 22215
rect 11630 22535 12000 22545
rect 11630 22475 11634 22535
rect 11686 22515 11944 22535
rect 11630 22469 11686 22475
rect 11630 22281 11660 22469
rect 11715 22460 11915 22485
rect 11996 22475 12000 22535
rect 11944 22469 12000 22475
rect 11715 22440 11785 22460
rect 11690 22400 11785 22440
rect 11845 22440 11915 22460
rect 11845 22400 11940 22440
rect 11690 22350 11940 22400
rect 11690 22310 11785 22350
rect 11715 22290 11785 22310
rect 11845 22310 11940 22350
rect 11845 22290 11915 22310
rect 11630 22275 11686 22281
rect 11630 22215 11634 22275
rect 11715 22265 11915 22290
rect 11970 22281 12000 22469
rect 11944 22275 12000 22281
rect 11686 22215 11944 22235
rect 11996 22215 12000 22275
rect 11630 22205 12000 22215
rect 12030 22535 12400 22545
rect 12030 22475 12034 22535
rect 12086 22515 12344 22535
rect 12030 22469 12086 22475
rect 12030 22281 12060 22469
rect 12115 22460 12315 22485
rect 12396 22475 12400 22535
rect 12344 22469 12400 22475
rect 12115 22440 12185 22460
rect 12090 22400 12185 22440
rect 12245 22440 12315 22460
rect 12245 22400 12340 22440
rect 12090 22350 12340 22400
rect 12090 22310 12185 22350
rect 12115 22290 12185 22310
rect 12245 22310 12340 22350
rect 12245 22290 12315 22310
rect 12030 22275 12086 22281
rect 12030 22215 12034 22275
rect 12115 22265 12315 22290
rect 12370 22281 12400 22469
rect 12344 22275 12400 22281
rect 12086 22215 12344 22235
rect 12396 22215 12400 22275
rect 12030 22205 12400 22215
rect 12430 22535 12800 22545
rect 12430 22475 12434 22535
rect 12486 22515 12744 22535
rect 12430 22469 12486 22475
rect 12430 22281 12460 22469
rect 12515 22460 12715 22485
rect 12796 22475 12800 22535
rect 12744 22469 12800 22475
rect 12515 22440 12585 22460
rect 12490 22400 12585 22440
rect 12645 22440 12715 22460
rect 12645 22400 12740 22440
rect 12490 22350 12740 22400
rect 12490 22310 12585 22350
rect 12515 22290 12585 22310
rect 12645 22310 12740 22350
rect 12645 22290 12715 22310
rect 12430 22275 12486 22281
rect 12430 22215 12434 22275
rect 12515 22265 12715 22290
rect 12770 22281 12800 22469
rect 12744 22275 12800 22281
rect 12486 22215 12744 22235
rect 12796 22215 12800 22275
rect 12430 22205 12800 22215
rect 12830 22535 13200 22545
rect 12830 22475 12834 22535
rect 12886 22515 13144 22535
rect 12830 22469 12886 22475
rect 12830 22281 12860 22469
rect 12915 22460 13115 22485
rect 13196 22475 13200 22535
rect 13144 22469 13200 22475
rect 12915 22440 12985 22460
rect 12890 22400 12985 22440
rect 13045 22440 13115 22460
rect 13045 22400 13140 22440
rect 12890 22350 13140 22400
rect 12890 22310 12985 22350
rect 12915 22290 12985 22310
rect 13045 22310 13140 22350
rect 13045 22290 13115 22310
rect 12830 22275 12886 22281
rect 12830 22215 12834 22275
rect 12915 22265 13115 22290
rect 13170 22281 13200 22469
rect 13144 22275 13200 22281
rect 12886 22215 13144 22235
rect 13196 22215 13200 22275
rect 12830 22205 13200 22215
rect -370 22165 0 22175
rect -370 22105 -366 22165
rect -314 22145 -56 22165
rect -370 22099 -314 22105
rect -370 21911 -340 22099
rect -285 22090 -85 22115
rect -4 22105 0 22165
rect -56 22099 0 22105
rect -285 22070 -215 22090
rect -310 22030 -215 22070
rect -155 22070 -85 22090
rect -155 22030 -60 22070
rect -310 21980 -60 22030
rect -310 21940 -215 21980
rect -285 21920 -215 21940
rect -155 21940 -60 21980
rect -155 21920 -85 21940
rect -370 21905 -314 21911
rect -370 21845 -366 21905
rect -285 21895 -85 21920
rect -30 21911 0 22099
rect -56 21905 0 21911
rect -314 21845 -56 21865
rect -4 21845 0 21905
rect -370 21835 0 21845
rect 30 22165 400 22175
rect 30 22105 34 22165
rect 86 22145 344 22165
rect 30 22099 86 22105
rect 30 21911 60 22099
rect 115 22090 315 22115
rect 396 22105 400 22165
rect 344 22099 400 22105
rect 115 22070 185 22090
rect 90 22030 185 22070
rect 245 22070 315 22090
rect 245 22030 340 22070
rect 90 21980 340 22030
rect 90 21940 185 21980
rect 115 21920 185 21940
rect 245 21940 340 21980
rect 245 21920 315 21940
rect 30 21905 86 21911
rect 30 21845 34 21905
rect 115 21895 315 21920
rect 370 21911 400 22099
rect 344 21905 400 21911
rect 86 21845 344 21865
rect 396 21845 400 21905
rect 30 21835 400 21845
rect 430 22165 800 22175
rect 430 22105 434 22165
rect 486 22145 744 22165
rect 430 22099 486 22105
rect 430 21911 460 22099
rect 515 22090 715 22115
rect 796 22105 800 22165
rect 744 22099 800 22105
rect 515 22070 585 22090
rect 490 22030 585 22070
rect 645 22070 715 22090
rect 645 22030 740 22070
rect 490 21980 740 22030
rect 490 21940 585 21980
rect 515 21920 585 21940
rect 645 21940 740 21980
rect 645 21920 715 21940
rect 430 21905 486 21911
rect 430 21845 434 21905
rect 515 21895 715 21920
rect 770 21911 800 22099
rect 744 21905 800 21911
rect 486 21845 744 21865
rect 796 21845 800 21905
rect 430 21835 800 21845
rect 830 22165 1200 22175
rect 830 22105 834 22165
rect 886 22145 1144 22165
rect 830 22099 886 22105
rect 830 21911 860 22099
rect 915 22090 1115 22115
rect 1196 22105 1200 22165
rect 1144 22099 1200 22105
rect 915 22070 985 22090
rect 890 22030 985 22070
rect 1045 22070 1115 22090
rect 1045 22030 1140 22070
rect 890 21980 1140 22030
rect 890 21940 985 21980
rect 915 21920 985 21940
rect 1045 21940 1140 21980
rect 1045 21920 1115 21940
rect 830 21905 886 21911
rect 830 21845 834 21905
rect 915 21895 1115 21920
rect 1170 21911 1200 22099
rect 1144 21905 1200 21911
rect 886 21845 1144 21865
rect 1196 21845 1200 21905
rect 830 21835 1200 21845
rect 1230 22165 1600 22175
rect 1230 22105 1234 22165
rect 1286 22145 1544 22165
rect 1230 22099 1286 22105
rect 1230 21911 1260 22099
rect 1315 22090 1515 22115
rect 1596 22105 1600 22165
rect 1544 22099 1600 22105
rect 1315 22070 1385 22090
rect 1290 22030 1385 22070
rect 1445 22070 1515 22090
rect 1445 22030 1540 22070
rect 1290 21980 1540 22030
rect 1290 21940 1385 21980
rect 1315 21920 1385 21940
rect 1445 21940 1540 21980
rect 1445 21920 1515 21940
rect 1230 21905 1286 21911
rect 1230 21845 1234 21905
rect 1315 21895 1515 21920
rect 1570 21911 1600 22099
rect 1544 21905 1600 21911
rect 1286 21845 1544 21865
rect 1596 21845 1600 21905
rect 1230 21835 1600 21845
rect 1630 22165 2000 22175
rect 1630 22105 1634 22165
rect 1686 22145 1944 22165
rect 1630 22099 1686 22105
rect 1630 21911 1660 22099
rect 1715 22090 1915 22115
rect 1996 22105 2000 22165
rect 1944 22099 2000 22105
rect 1715 22070 1785 22090
rect 1690 22030 1785 22070
rect 1845 22070 1915 22090
rect 1845 22030 1940 22070
rect 1690 21980 1940 22030
rect 1690 21940 1785 21980
rect 1715 21920 1785 21940
rect 1845 21940 1940 21980
rect 1845 21920 1915 21940
rect 1630 21905 1686 21911
rect 1630 21845 1634 21905
rect 1715 21895 1915 21920
rect 1970 21911 2000 22099
rect 1944 21905 2000 21911
rect 1686 21845 1944 21865
rect 1996 21845 2000 21905
rect 1630 21835 2000 21845
rect 2030 22165 2400 22175
rect 2030 22105 2034 22165
rect 2086 22145 2344 22165
rect 2030 22099 2086 22105
rect 2030 21911 2060 22099
rect 2115 22090 2315 22115
rect 2396 22105 2400 22165
rect 2344 22099 2400 22105
rect 2115 22070 2185 22090
rect 2090 22030 2185 22070
rect 2245 22070 2315 22090
rect 2245 22030 2340 22070
rect 2090 21980 2340 22030
rect 2090 21940 2185 21980
rect 2115 21920 2185 21940
rect 2245 21940 2340 21980
rect 2245 21920 2315 21940
rect 2030 21905 2086 21911
rect 2030 21845 2034 21905
rect 2115 21895 2315 21920
rect 2370 21911 2400 22099
rect 2344 21905 2400 21911
rect 2086 21845 2344 21865
rect 2396 21845 2400 21905
rect 2030 21835 2400 21845
rect 2430 22165 2800 22175
rect 2430 22105 2434 22165
rect 2486 22145 2744 22165
rect 2430 22099 2486 22105
rect 2430 21911 2460 22099
rect 2515 22090 2715 22115
rect 2796 22105 2800 22165
rect 2744 22099 2800 22105
rect 2515 22070 2585 22090
rect 2490 22030 2585 22070
rect 2645 22070 2715 22090
rect 2645 22030 2740 22070
rect 2490 21980 2740 22030
rect 2490 21940 2585 21980
rect 2515 21920 2585 21940
rect 2645 21940 2740 21980
rect 2645 21920 2715 21940
rect 2430 21905 2486 21911
rect 2430 21845 2434 21905
rect 2515 21895 2715 21920
rect 2770 21911 2800 22099
rect 2744 21905 2800 21911
rect 2486 21845 2744 21865
rect 2796 21845 2800 21905
rect 2430 21835 2800 21845
rect 2830 22165 3200 22175
rect 2830 22105 2834 22165
rect 2886 22145 3144 22165
rect 2830 22099 2886 22105
rect 2830 21911 2860 22099
rect 2915 22090 3115 22115
rect 3196 22105 3200 22165
rect 3144 22099 3200 22105
rect 2915 22070 2985 22090
rect 2890 22030 2985 22070
rect 3045 22070 3115 22090
rect 3045 22030 3140 22070
rect 2890 21980 3140 22030
rect 2890 21940 2985 21980
rect 2915 21920 2985 21940
rect 3045 21940 3140 21980
rect 3045 21920 3115 21940
rect 2830 21905 2886 21911
rect 2830 21845 2834 21905
rect 2915 21895 3115 21920
rect 3170 21911 3200 22099
rect 3144 21905 3200 21911
rect 2886 21845 3144 21865
rect 3196 21845 3200 21905
rect 2830 21835 3200 21845
rect 3230 22165 3600 22175
rect 3230 22105 3234 22165
rect 3286 22145 3544 22165
rect 3230 22099 3286 22105
rect 3230 21911 3260 22099
rect 3315 22090 3515 22115
rect 3596 22105 3600 22165
rect 3544 22099 3600 22105
rect 3315 22070 3385 22090
rect 3290 22030 3385 22070
rect 3445 22070 3515 22090
rect 3445 22030 3540 22070
rect 3290 21980 3540 22030
rect 3290 21940 3385 21980
rect 3315 21920 3385 21940
rect 3445 21940 3540 21980
rect 3445 21920 3515 21940
rect 3230 21905 3286 21911
rect 3230 21845 3234 21905
rect 3315 21895 3515 21920
rect 3570 21911 3600 22099
rect 3544 21905 3600 21911
rect 3286 21845 3544 21865
rect 3596 21845 3600 21905
rect 3230 21835 3600 21845
rect 3630 22165 4000 22175
rect 3630 22105 3634 22165
rect 3686 22145 3944 22165
rect 3630 22099 3686 22105
rect 3630 21911 3660 22099
rect 3715 22090 3915 22115
rect 3996 22105 4000 22165
rect 3944 22099 4000 22105
rect 3715 22070 3785 22090
rect 3690 22030 3785 22070
rect 3845 22070 3915 22090
rect 3845 22030 3940 22070
rect 3690 21980 3940 22030
rect 3690 21940 3785 21980
rect 3715 21920 3785 21940
rect 3845 21940 3940 21980
rect 3845 21920 3915 21940
rect 3630 21905 3686 21911
rect 3630 21845 3634 21905
rect 3715 21895 3915 21920
rect 3970 21911 4000 22099
rect 3944 21905 4000 21911
rect 3686 21845 3944 21865
rect 3996 21845 4000 21905
rect 3630 21835 4000 21845
rect 4030 22165 4400 22175
rect 4030 22105 4034 22165
rect 4086 22145 4344 22165
rect 4030 22099 4086 22105
rect 4030 21911 4060 22099
rect 4115 22090 4315 22115
rect 4396 22105 4400 22165
rect 4344 22099 4400 22105
rect 4115 22070 4185 22090
rect 4090 22030 4185 22070
rect 4245 22070 4315 22090
rect 4245 22030 4340 22070
rect 4090 21980 4340 22030
rect 4090 21940 4185 21980
rect 4115 21920 4185 21940
rect 4245 21940 4340 21980
rect 4245 21920 4315 21940
rect 4030 21905 4086 21911
rect 4030 21845 4034 21905
rect 4115 21895 4315 21920
rect 4370 21911 4400 22099
rect 4344 21905 4400 21911
rect 4086 21845 4344 21865
rect 4396 21845 4400 21905
rect 4030 21835 4400 21845
rect 4430 22165 4800 22175
rect 4430 22105 4434 22165
rect 4486 22145 4744 22165
rect 4430 22099 4486 22105
rect 4430 21911 4460 22099
rect 4515 22090 4715 22115
rect 4796 22105 4800 22165
rect 4744 22099 4800 22105
rect 4515 22070 4585 22090
rect 4490 22030 4585 22070
rect 4645 22070 4715 22090
rect 4645 22030 4740 22070
rect 4490 21980 4740 22030
rect 4490 21940 4585 21980
rect 4515 21920 4585 21940
rect 4645 21940 4740 21980
rect 4645 21920 4715 21940
rect 4430 21905 4486 21911
rect 4430 21845 4434 21905
rect 4515 21895 4715 21920
rect 4770 21911 4800 22099
rect 4744 21905 4800 21911
rect 4486 21845 4744 21865
rect 4796 21845 4800 21905
rect 4430 21835 4800 21845
rect 4830 22165 5200 22175
rect 4830 22105 4834 22165
rect 4886 22145 5144 22165
rect 4830 22099 4886 22105
rect 4830 21911 4860 22099
rect 4915 22090 5115 22115
rect 5196 22105 5200 22165
rect 5144 22099 5200 22105
rect 4915 22070 4985 22090
rect 4890 22030 4985 22070
rect 5045 22070 5115 22090
rect 5045 22030 5140 22070
rect 4890 21980 5140 22030
rect 4890 21940 4985 21980
rect 4915 21920 4985 21940
rect 5045 21940 5140 21980
rect 5045 21920 5115 21940
rect 4830 21905 4886 21911
rect 4830 21845 4834 21905
rect 4915 21895 5115 21920
rect 5170 21911 5200 22099
rect 5144 21905 5200 21911
rect 4886 21845 5144 21865
rect 5196 21845 5200 21905
rect 4830 21835 5200 21845
rect 5230 22165 5600 22175
rect 5230 22105 5234 22165
rect 5286 22145 5544 22165
rect 5230 22099 5286 22105
rect 5230 21911 5260 22099
rect 5315 22090 5515 22115
rect 5596 22105 5600 22165
rect 5544 22099 5600 22105
rect 5315 22070 5385 22090
rect 5290 22030 5385 22070
rect 5445 22070 5515 22090
rect 5445 22030 5540 22070
rect 5290 21980 5540 22030
rect 5290 21940 5385 21980
rect 5315 21920 5385 21940
rect 5445 21940 5540 21980
rect 5445 21920 5515 21940
rect 5230 21905 5286 21911
rect 5230 21845 5234 21905
rect 5315 21895 5515 21920
rect 5570 21911 5600 22099
rect 5544 21905 5600 21911
rect 5286 21845 5544 21865
rect 5596 21845 5600 21905
rect 5230 21835 5600 21845
rect 5630 22165 6000 22175
rect 5630 22105 5634 22165
rect 5686 22145 5944 22165
rect 5630 22099 5686 22105
rect 5630 21911 5660 22099
rect 5715 22090 5915 22115
rect 5996 22105 6000 22165
rect 5944 22099 6000 22105
rect 5715 22070 5785 22090
rect 5690 22030 5785 22070
rect 5845 22070 5915 22090
rect 5845 22030 5940 22070
rect 5690 21980 5940 22030
rect 5690 21940 5785 21980
rect 5715 21920 5785 21940
rect 5845 21940 5940 21980
rect 5845 21920 5915 21940
rect 5630 21905 5686 21911
rect 5630 21845 5634 21905
rect 5715 21895 5915 21920
rect 5970 21911 6000 22099
rect 5944 21905 6000 21911
rect 5686 21845 5944 21865
rect 5996 21845 6000 21905
rect 5630 21835 6000 21845
rect 6030 22165 6400 22175
rect 6030 22105 6034 22165
rect 6086 22145 6344 22165
rect 6030 22099 6086 22105
rect 6030 21911 6060 22099
rect 6115 22090 6315 22115
rect 6396 22105 6400 22165
rect 6344 22099 6400 22105
rect 6115 22070 6185 22090
rect 6090 22030 6185 22070
rect 6245 22070 6315 22090
rect 6245 22030 6340 22070
rect 6090 21980 6340 22030
rect 6090 21940 6185 21980
rect 6115 21920 6185 21940
rect 6245 21940 6340 21980
rect 6245 21920 6315 21940
rect 6030 21905 6086 21911
rect 6030 21845 6034 21905
rect 6115 21895 6315 21920
rect 6370 21911 6400 22099
rect 6344 21905 6400 21911
rect 6086 21845 6344 21865
rect 6396 21845 6400 21905
rect 6030 21835 6400 21845
rect 6430 22165 6800 22175
rect 6430 22105 6434 22165
rect 6486 22145 6744 22165
rect 6430 22099 6486 22105
rect 6430 21911 6460 22099
rect 6515 22090 6715 22115
rect 6796 22105 6800 22165
rect 6744 22099 6800 22105
rect 6515 22070 6585 22090
rect 6490 22030 6585 22070
rect 6645 22070 6715 22090
rect 6645 22030 6740 22070
rect 6490 21980 6740 22030
rect 6490 21940 6585 21980
rect 6515 21920 6585 21940
rect 6645 21940 6740 21980
rect 6645 21920 6715 21940
rect 6430 21905 6486 21911
rect 6430 21845 6434 21905
rect 6515 21895 6715 21920
rect 6770 21911 6800 22099
rect 6744 21905 6800 21911
rect 6486 21845 6744 21865
rect 6796 21845 6800 21905
rect 6430 21835 6800 21845
rect 6830 22165 7200 22175
rect 6830 22105 6834 22165
rect 6886 22145 7144 22165
rect 6830 22099 6886 22105
rect 6830 21911 6860 22099
rect 6915 22090 7115 22115
rect 7196 22105 7200 22165
rect 7144 22099 7200 22105
rect 6915 22070 6985 22090
rect 6890 22030 6985 22070
rect 7045 22070 7115 22090
rect 7045 22030 7140 22070
rect 6890 21980 7140 22030
rect 6890 21940 6985 21980
rect 6915 21920 6985 21940
rect 7045 21940 7140 21980
rect 7045 21920 7115 21940
rect 6830 21905 6886 21911
rect 6830 21845 6834 21905
rect 6915 21895 7115 21920
rect 7170 21911 7200 22099
rect 7144 21905 7200 21911
rect 6886 21845 7144 21865
rect 7196 21845 7200 21905
rect 6830 21835 7200 21845
rect 7230 22165 7600 22175
rect 7230 22105 7234 22165
rect 7286 22145 7544 22165
rect 7230 22099 7286 22105
rect 7230 21911 7260 22099
rect 7315 22090 7515 22115
rect 7596 22105 7600 22165
rect 7544 22099 7600 22105
rect 7315 22070 7385 22090
rect 7290 22030 7385 22070
rect 7445 22070 7515 22090
rect 7445 22030 7540 22070
rect 7290 21980 7540 22030
rect 7290 21940 7385 21980
rect 7315 21920 7385 21940
rect 7445 21940 7540 21980
rect 7445 21920 7515 21940
rect 7230 21905 7286 21911
rect 7230 21845 7234 21905
rect 7315 21895 7515 21920
rect 7570 21911 7600 22099
rect 7544 21905 7600 21911
rect 7286 21845 7544 21865
rect 7596 21845 7600 21905
rect 7230 21835 7600 21845
rect 7630 22165 8000 22175
rect 7630 22105 7634 22165
rect 7686 22145 7944 22165
rect 7630 22099 7686 22105
rect 7630 21911 7660 22099
rect 7715 22090 7915 22115
rect 7996 22105 8000 22165
rect 7944 22099 8000 22105
rect 7715 22070 7785 22090
rect 7690 22030 7785 22070
rect 7845 22070 7915 22090
rect 7845 22030 7940 22070
rect 7690 21980 7940 22030
rect 7690 21940 7785 21980
rect 7715 21920 7785 21940
rect 7845 21940 7940 21980
rect 7845 21920 7915 21940
rect 7630 21905 7686 21911
rect 7630 21845 7634 21905
rect 7715 21895 7915 21920
rect 7970 21911 8000 22099
rect 7944 21905 8000 21911
rect 7686 21845 7944 21865
rect 7996 21845 8000 21905
rect 7630 21835 8000 21845
rect 8030 22165 8400 22175
rect 8030 22105 8034 22165
rect 8086 22145 8344 22165
rect 8030 22099 8086 22105
rect 8030 21911 8060 22099
rect 8115 22090 8315 22115
rect 8396 22105 8400 22165
rect 8344 22099 8400 22105
rect 8115 22070 8185 22090
rect 8090 22030 8185 22070
rect 8245 22070 8315 22090
rect 8245 22030 8340 22070
rect 8090 21980 8340 22030
rect 8090 21940 8185 21980
rect 8115 21920 8185 21940
rect 8245 21940 8340 21980
rect 8245 21920 8315 21940
rect 8030 21905 8086 21911
rect 8030 21845 8034 21905
rect 8115 21895 8315 21920
rect 8370 21911 8400 22099
rect 8344 21905 8400 21911
rect 8086 21845 8344 21865
rect 8396 21845 8400 21905
rect 8030 21835 8400 21845
rect 8430 22165 8800 22175
rect 8430 22105 8434 22165
rect 8486 22145 8744 22165
rect 8430 22099 8486 22105
rect 8430 21911 8460 22099
rect 8515 22090 8715 22115
rect 8796 22105 8800 22165
rect 8744 22099 8800 22105
rect 8515 22070 8585 22090
rect 8490 22030 8585 22070
rect 8645 22070 8715 22090
rect 8645 22030 8740 22070
rect 8490 21980 8740 22030
rect 8490 21940 8585 21980
rect 8515 21920 8585 21940
rect 8645 21940 8740 21980
rect 8645 21920 8715 21940
rect 8430 21905 8486 21911
rect 8430 21845 8434 21905
rect 8515 21895 8715 21920
rect 8770 21911 8800 22099
rect 8744 21905 8800 21911
rect 8486 21845 8744 21865
rect 8796 21845 8800 21905
rect 8430 21835 8800 21845
rect 8830 22165 9200 22175
rect 8830 22105 8834 22165
rect 8886 22145 9144 22165
rect 8830 22099 8886 22105
rect 8830 21911 8860 22099
rect 8915 22090 9115 22115
rect 9196 22105 9200 22165
rect 9144 22099 9200 22105
rect 8915 22070 8985 22090
rect 8890 22030 8985 22070
rect 9045 22070 9115 22090
rect 9045 22030 9140 22070
rect 8890 21980 9140 22030
rect 8890 21940 8985 21980
rect 8915 21920 8985 21940
rect 9045 21940 9140 21980
rect 9045 21920 9115 21940
rect 8830 21905 8886 21911
rect 8830 21845 8834 21905
rect 8915 21895 9115 21920
rect 9170 21911 9200 22099
rect 9144 21905 9200 21911
rect 8886 21845 9144 21865
rect 9196 21845 9200 21905
rect 8830 21835 9200 21845
rect 9230 22165 9600 22175
rect 9230 22105 9234 22165
rect 9286 22145 9544 22165
rect 9230 22099 9286 22105
rect 9230 21911 9260 22099
rect 9315 22090 9515 22115
rect 9596 22105 9600 22165
rect 9544 22099 9600 22105
rect 9315 22070 9385 22090
rect 9290 22030 9385 22070
rect 9445 22070 9515 22090
rect 9445 22030 9540 22070
rect 9290 21980 9540 22030
rect 9290 21940 9385 21980
rect 9315 21920 9385 21940
rect 9445 21940 9540 21980
rect 9445 21920 9515 21940
rect 9230 21905 9286 21911
rect 9230 21845 9234 21905
rect 9315 21895 9515 21920
rect 9570 21911 9600 22099
rect 9544 21905 9600 21911
rect 9286 21845 9544 21865
rect 9596 21845 9600 21905
rect 9230 21835 9600 21845
rect 9630 22165 10000 22175
rect 9630 22105 9634 22165
rect 9686 22145 9944 22165
rect 9630 22099 9686 22105
rect 9630 21911 9660 22099
rect 9715 22090 9915 22115
rect 9996 22105 10000 22165
rect 9944 22099 10000 22105
rect 9715 22070 9785 22090
rect 9690 22030 9785 22070
rect 9845 22070 9915 22090
rect 9845 22030 9940 22070
rect 9690 21980 9940 22030
rect 9690 21940 9785 21980
rect 9715 21920 9785 21940
rect 9845 21940 9940 21980
rect 9845 21920 9915 21940
rect 9630 21905 9686 21911
rect 9630 21845 9634 21905
rect 9715 21895 9915 21920
rect 9970 21911 10000 22099
rect 9944 21905 10000 21911
rect 9686 21845 9944 21865
rect 9996 21845 10000 21905
rect 9630 21835 10000 21845
rect 10030 22165 10400 22175
rect 10030 22105 10034 22165
rect 10086 22145 10344 22165
rect 10030 22099 10086 22105
rect 10030 21911 10060 22099
rect 10115 22090 10315 22115
rect 10396 22105 10400 22165
rect 10344 22099 10400 22105
rect 10115 22070 10185 22090
rect 10090 22030 10185 22070
rect 10245 22070 10315 22090
rect 10245 22030 10340 22070
rect 10090 21980 10340 22030
rect 10090 21940 10185 21980
rect 10115 21920 10185 21940
rect 10245 21940 10340 21980
rect 10245 21920 10315 21940
rect 10030 21905 10086 21911
rect 10030 21845 10034 21905
rect 10115 21895 10315 21920
rect 10370 21911 10400 22099
rect 10344 21905 10400 21911
rect 10086 21845 10344 21865
rect 10396 21845 10400 21905
rect 10030 21835 10400 21845
rect 10430 22165 10800 22175
rect 10430 22105 10434 22165
rect 10486 22145 10744 22165
rect 10430 22099 10486 22105
rect 10430 21911 10460 22099
rect 10515 22090 10715 22115
rect 10796 22105 10800 22165
rect 10744 22099 10800 22105
rect 10515 22070 10585 22090
rect 10490 22030 10585 22070
rect 10645 22070 10715 22090
rect 10645 22030 10740 22070
rect 10490 21980 10740 22030
rect 10490 21940 10585 21980
rect 10515 21920 10585 21940
rect 10645 21940 10740 21980
rect 10645 21920 10715 21940
rect 10430 21905 10486 21911
rect 10430 21845 10434 21905
rect 10515 21895 10715 21920
rect 10770 21911 10800 22099
rect 10744 21905 10800 21911
rect 10486 21845 10744 21865
rect 10796 21845 10800 21905
rect 10430 21835 10800 21845
rect 10830 22165 11200 22175
rect 10830 22105 10834 22165
rect 10886 22145 11144 22165
rect 10830 22099 10886 22105
rect 10830 21911 10860 22099
rect 10915 22090 11115 22115
rect 11196 22105 11200 22165
rect 11144 22099 11200 22105
rect 10915 22070 10985 22090
rect 10890 22030 10985 22070
rect 11045 22070 11115 22090
rect 11045 22030 11140 22070
rect 10890 21980 11140 22030
rect 10890 21940 10985 21980
rect 10915 21920 10985 21940
rect 11045 21940 11140 21980
rect 11045 21920 11115 21940
rect 10830 21905 10886 21911
rect 10830 21845 10834 21905
rect 10915 21895 11115 21920
rect 11170 21911 11200 22099
rect 11144 21905 11200 21911
rect 10886 21845 11144 21865
rect 11196 21845 11200 21905
rect 10830 21835 11200 21845
rect 11230 22165 11600 22175
rect 11230 22105 11234 22165
rect 11286 22145 11544 22165
rect 11230 22099 11286 22105
rect 11230 21911 11260 22099
rect 11315 22090 11515 22115
rect 11596 22105 11600 22165
rect 11544 22099 11600 22105
rect 11315 22070 11385 22090
rect 11290 22030 11385 22070
rect 11445 22070 11515 22090
rect 11445 22030 11540 22070
rect 11290 21980 11540 22030
rect 11290 21940 11385 21980
rect 11315 21920 11385 21940
rect 11445 21940 11540 21980
rect 11445 21920 11515 21940
rect 11230 21905 11286 21911
rect 11230 21845 11234 21905
rect 11315 21895 11515 21920
rect 11570 21911 11600 22099
rect 11544 21905 11600 21911
rect 11286 21845 11544 21865
rect 11596 21845 11600 21905
rect 11230 21835 11600 21845
rect 11630 22165 12000 22175
rect 11630 22105 11634 22165
rect 11686 22145 11944 22165
rect 11630 22099 11686 22105
rect 11630 21911 11660 22099
rect 11715 22090 11915 22115
rect 11996 22105 12000 22165
rect 11944 22099 12000 22105
rect 11715 22070 11785 22090
rect 11690 22030 11785 22070
rect 11845 22070 11915 22090
rect 11845 22030 11940 22070
rect 11690 21980 11940 22030
rect 11690 21940 11785 21980
rect 11715 21920 11785 21940
rect 11845 21940 11940 21980
rect 11845 21920 11915 21940
rect 11630 21905 11686 21911
rect 11630 21845 11634 21905
rect 11715 21895 11915 21920
rect 11970 21911 12000 22099
rect 11944 21905 12000 21911
rect 11686 21845 11944 21865
rect 11996 21845 12000 21905
rect 11630 21835 12000 21845
rect 12030 22165 12400 22175
rect 12030 22105 12034 22165
rect 12086 22145 12344 22165
rect 12030 22099 12086 22105
rect 12030 21911 12060 22099
rect 12115 22090 12315 22115
rect 12396 22105 12400 22165
rect 12344 22099 12400 22105
rect 12115 22070 12185 22090
rect 12090 22030 12185 22070
rect 12245 22070 12315 22090
rect 12245 22030 12340 22070
rect 12090 21980 12340 22030
rect 12090 21940 12185 21980
rect 12115 21920 12185 21940
rect 12245 21940 12340 21980
rect 12245 21920 12315 21940
rect 12030 21905 12086 21911
rect 12030 21845 12034 21905
rect 12115 21895 12315 21920
rect 12370 21911 12400 22099
rect 12344 21905 12400 21911
rect 12086 21845 12344 21865
rect 12396 21845 12400 21905
rect 12030 21835 12400 21845
rect 12430 22165 12800 22175
rect 12430 22105 12434 22165
rect 12486 22145 12744 22165
rect 12430 22099 12486 22105
rect 12430 21911 12460 22099
rect 12515 22090 12715 22115
rect 12796 22105 12800 22165
rect 12744 22099 12800 22105
rect 12515 22070 12585 22090
rect 12490 22030 12585 22070
rect 12645 22070 12715 22090
rect 12645 22030 12740 22070
rect 12490 21980 12740 22030
rect 12490 21940 12585 21980
rect 12515 21920 12585 21940
rect 12645 21940 12740 21980
rect 12645 21920 12715 21940
rect 12430 21905 12486 21911
rect 12430 21845 12434 21905
rect 12515 21895 12715 21920
rect 12770 21911 12800 22099
rect 12744 21905 12800 21911
rect 12486 21845 12744 21865
rect 12796 21845 12800 21905
rect 12430 21835 12800 21845
rect 12830 22165 13200 22175
rect 12830 22105 12834 22165
rect 12886 22145 13144 22165
rect 12830 22099 12886 22105
rect 12830 21911 12860 22099
rect 12915 22090 13115 22115
rect 13196 22105 13200 22165
rect 13144 22099 13200 22105
rect 12915 22070 12985 22090
rect 12890 22030 12985 22070
rect 13045 22070 13115 22090
rect 13045 22030 13140 22070
rect 12890 21980 13140 22030
rect 12890 21940 12985 21980
rect 12915 21920 12985 21940
rect 13045 21940 13140 21980
rect 13045 21920 13115 21940
rect 12830 21905 12886 21911
rect 12830 21845 12834 21905
rect 12915 21895 13115 21920
rect 13170 21911 13200 22099
rect 13144 21905 13200 21911
rect 12886 21845 13144 21865
rect 13196 21845 13200 21905
rect 12830 21835 13200 21845
rect -370 21795 0 21805
rect -370 21735 -366 21795
rect -314 21775 -56 21795
rect -370 21729 -314 21735
rect -370 21541 -340 21729
rect -285 21720 -85 21745
rect -4 21735 0 21795
rect -56 21729 0 21735
rect -285 21700 -215 21720
rect -310 21660 -215 21700
rect -155 21700 -85 21720
rect -155 21660 -60 21700
rect -310 21610 -60 21660
rect -310 21570 -215 21610
rect -285 21550 -215 21570
rect -155 21570 -60 21610
rect -155 21550 -85 21570
rect -370 21535 -314 21541
rect -370 21475 -366 21535
rect -285 21525 -85 21550
rect -30 21541 0 21729
rect -56 21535 0 21541
rect -314 21475 -56 21495
rect -4 21475 0 21535
rect -370 21465 0 21475
rect 30 21795 400 21805
rect 30 21735 34 21795
rect 86 21775 344 21795
rect 30 21729 86 21735
rect 30 21541 60 21729
rect 115 21720 315 21745
rect 396 21735 400 21795
rect 344 21729 400 21735
rect 115 21700 185 21720
rect 90 21660 185 21700
rect 245 21700 315 21720
rect 245 21660 340 21700
rect 90 21610 340 21660
rect 90 21570 185 21610
rect 115 21550 185 21570
rect 245 21570 340 21610
rect 245 21550 315 21570
rect 30 21535 86 21541
rect 30 21475 34 21535
rect 115 21525 315 21550
rect 370 21541 400 21729
rect 344 21535 400 21541
rect 86 21475 344 21495
rect 396 21475 400 21535
rect 30 21465 400 21475
rect 430 21795 800 21805
rect 430 21735 434 21795
rect 486 21775 744 21795
rect 430 21729 486 21735
rect 430 21541 460 21729
rect 515 21720 715 21745
rect 796 21735 800 21795
rect 744 21729 800 21735
rect 515 21700 585 21720
rect 490 21660 585 21700
rect 645 21700 715 21720
rect 645 21660 740 21700
rect 490 21610 740 21660
rect 490 21570 585 21610
rect 515 21550 585 21570
rect 645 21570 740 21610
rect 645 21550 715 21570
rect 430 21535 486 21541
rect 430 21475 434 21535
rect 515 21525 715 21550
rect 770 21541 800 21729
rect 744 21535 800 21541
rect 486 21475 744 21495
rect 796 21475 800 21535
rect 430 21465 800 21475
rect 830 21795 1200 21805
rect 830 21735 834 21795
rect 886 21775 1144 21795
rect 830 21729 886 21735
rect 830 21541 860 21729
rect 915 21720 1115 21745
rect 1196 21735 1200 21795
rect 1144 21729 1200 21735
rect 915 21700 985 21720
rect 890 21660 985 21700
rect 1045 21700 1115 21720
rect 1045 21660 1140 21700
rect 890 21610 1140 21660
rect 890 21570 985 21610
rect 915 21550 985 21570
rect 1045 21570 1140 21610
rect 1045 21550 1115 21570
rect 830 21535 886 21541
rect 830 21475 834 21535
rect 915 21525 1115 21550
rect 1170 21541 1200 21729
rect 1144 21535 1200 21541
rect 886 21475 1144 21495
rect 1196 21475 1200 21535
rect 830 21465 1200 21475
rect 1230 21795 1600 21805
rect 1230 21735 1234 21795
rect 1286 21775 1544 21795
rect 1230 21729 1286 21735
rect 1230 21541 1260 21729
rect 1315 21720 1515 21745
rect 1596 21735 1600 21795
rect 1544 21729 1600 21735
rect 1315 21700 1385 21720
rect 1290 21660 1385 21700
rect 1445 21700 1515 21720
rect 1445 21660 1540 21700
rect 1290 21610 1540 21660
rect 1290 21570 1385 21610
rect 1315 21550 1385 21570
rect 1445 21570 1540 21610
rect 1445 21550 1515 21570
rect 1230 21535 1286 21541
rect 1230 21475 1234 21535
rect 1315 21525 1515 21550
rect 1570 21541 1600 21729
rect 1544 21535 1600 21541
rect 1286 21475 1544 21495
rect 1596 21475 1600 21535
rect 1230 21465 1600 21475
rect 1630 21795 2000 21805
rect 1630 21735 1634 21795
rect 1686 21775 1944 21795
rect 1630 21729 1686 21735
rect 1630 21541 1660 21729
rect 1715 21720 1915 21745
rect 1996 21735 2000 21795
rect 1944 21729 2000 21735
rect 1715 21700 1785 21720
rect 1690 21660 1785 21700
rect 1845 21700 1915 21720
rect 1845 21660 1940 21700
rect 1690 21610 1940 21660
rect 1690 21570 1785 21610
rect 1715 21550 1785 21570
rect 1845 21570 1940 21610
rect 1845 21550 1915 21570
rect 1630 21535 1686 21541
rect 1630 21475 1634 21535
rect 1715 21525 1915 21550
rect 1970 21541 2000 21729
rect 1944 21535 2000 21541
rect 1686 21475 1944 21495
rect 1996 21475 2000 21535
rect 1630 21465 2000 21475
rect 2030 21795 2400 21805
rect 2030 21735 2034 21795
rect 2086 21775 2344 21795
rect 2030 21729 2086 21735
rect 2030 21541 2060 21729
rect 2115 21720 2315 21745
rect 2396 21735 2400 21795
rect 2344 21729 2400 21735
rect 2115 21700 2185 21720
rect 2090 21660 2185 21700
rect 2245 21700 2315 21720
rect 2245 21660 2340 21700
rect 2090 21610 2340 21660
rect 2090 21570 2185 21610
rect 2115 21550 2185 21570
rect 2245 21570 2340 21610
rect 2245 21550 2315 21570
rect 2030 21535 2086 21541
rect 2030 21475 2034 21535
rect 2115 21525 2315 21550
rect 2370 21541 2400 21729
rect 2344 21535 2400 21541
rect 2086 21475 2344 21495
rect 2396 21475 2400 21535
rect 2030 21465 2400 21475
rect 2430 21795 2800 21805
rect 2430 21735 2434 21795
rect 2486 21775 2744 21795
rect 2430 21729 2486 21735
rect 2430 21541 2460 21729
rect 2515 21720 2715 21745
rect 2796 21735 2800 21795
rect 2744 21729 2800 21735
rect 2515 21700 2585 21720
rect 2490 21660 2585 21700
rect 2645 21700 2715 21720
rect 2645 21660 2740 21700
rect 2490 21610 2740 21660
rect 2490 21570 2585 21610
rect 2515 21550 2585 21570
rect 2645 21570 2740 21610
rect 2645 21550 2715 21570
rect 2430 21535 2486 21541
rect 2430 21475 2434 21535
rect 2515 21525 2715 21550
rect 2770 21541 2800 21729
rect 2744 21535 2800 21541
rect 2486 21475 2744 21495
rect 2796 21475 2800 21535
rect 2430 21465 2800 21475
rect 2830 21795 3200 21805
rect 2830 21735 2834 21795
rect 2886 21775 3144 21795
rect 2830 21729 2886 21735
rect 2830 21541 2860 21729
rect 2915 21720 3115 21745
rect 3196 21735 3200 21795
rect 3144 21729 3200 21735
rect 2915 21700 2985 21720
rect 2890 21660 2985 21700
rect 3045 21700 3115 21720
rect 3045 21660 3140 21700
rect 2890 21610 3140 21660
rect 2890 21570 2985 21610
rect 2915 21550 2985 21570
rect 3045 21570 3140 21610
rect 3045 21550 3115 21570
rect 2830 21535 2886 21541
rect 2830 21475 2834 21535
rect 2915 21525 3115 21550
rect 3170 21541 3200 21729
rect 3144 21535 3200 21541
rect 2886 21475 3144 21495
rect 3196 21475 3200 21535
rect 2830 21465 3200 21475
rect 3230 21795 3600 21805
rect 3230 21735 3234 21795
rect 3286 21775 3544 21795
rect 3230 21729 3286 21735
rect 3230 21541 3260 21729
rect 3315 21720 3515 21745
rect 3596 21735 3600 21795
rect 3544 21729 3600 21735
rect 3315 21700 3385 21720
rect 3290 21660 3385 21700
rect 3445 21700 3515 21720
rect 3445 21660 3540 21700
rect 3290 21610 3540 21660
rect 3290 21570 3385 21610
rect 3315 21550 3385 21570
rect 3445 21570 3540 21610
rect 3445 21550 3515 21570
rect 3230 21535 3286 21541
rect 3230 21475 3234 21535
rect 3315 21525 3515 21550
rect 3570 21541 3600 21729
rect 3544 21535 3600 21541
rect 3286 21475 3544 21495
rect 3596 21475 3600 21535
rect 3230 21465 3600 21475
rect 3630 21795 4000 21805
rect 3630 21735 3634 21795
rect 3686 21775 3944 21795
rect 3630 21729 3686 21735
rect 3630 21541 3660 21729
rect 3715 21720 3915 21745
rect 3996 21735 4000 21795
rect 3944 21729 4000 21735
rect 3715 21700 3785 21720
rect 3690 21660 3785 21700
rect 3845 21700 3915 21720
rect 3845 21660 3940 21700
rect 3690 21610 3940 21660
rect 3690 21570 3785 21610
rect 3715 21550 3785 21570
rect 3845 21570 3940 21610
rect 3845 21550 3915 21570
rect 3630 21535 3686 21541
rect 3630 21475 3634 21535
rect 3715 21525 3915 21550
rect 3970 21541 4000 21729
rect 3944 21535 4000 21541
rect 3686 21475 3944 21495
rect 3996 21475 4000 21535
rect 3630 21465 4000 21475
rect 4030 21795 4400 21805
rect 4030 21735 4034 21795
rect 4086 21775 4344 21795
rect 4030 21729 4086 21735
rect 4030 21541 4060 21729
rect 4115 21720 4315 21745
rect 4396 21735 4400 21795
rect 4344 21729 4400 21735
rect 4115 21700 4185 21720
rect 4090 21660 4185 21700
rect 4245 21700 4315 21720
rect 4245 21660 4340 21700
rect 4090 21610 4340 21660
rect 4090 21570 4185 21610
rect 4115 21550 4185 21570
rect 4245 21570 4340 21610
rect 4245 21550 4315 21570
rect 4030 21535 4086 21541
rect 4030 21475 4034 21535
rect 4115 21525 4315 21550
rect 4370 21541 4400 21729
rect 4344 21535 4400 21541
rect 4086 21475 4344 21495
rect 4396 21475 4400 21535
rect 4030 21465 4400 21475
rect 4430 21795 4800 21805
rect 4430 21735 4434 21795
rect 4486 21775 4744 21795
rect 4430 21729 4486 21735
rect 4430 21541 4460 21729
rect 4515 21720 4715 21745
rect 4796 21735 4800 21795
rect 4744 21729 4800 21735
rect 4515 21700 4585 21720
rect 4490 21660 4585 21700
rect 4645 21700 4715 21720
rect 4645 21660 4740 21700
rect 4490 21610 4740 21660
rect 4490 21570 4585 21610
rect 4515 21550 4585 21570
rect 4645 21570 4740 21610
rect 4645 21550 4715 21570
rect 4430 21535 4486 21541
rect 4430 21475 4434 21535
rect 4515 21525 4715 21550
rect 4770 21541 4800 21729
rect 4744 21535 4800 21541
rect 4486 21475 4744 21495
rect 4796 21475 4800 21535
rect 4430 21465 4800 21475
rect 4830 21795 5200 21805
rect 4830 21735 4834 21795
rect 4886 21775 5144 21795
rect 4830 21729 4886 21735
rect 4830 21541 4860 21729
rect 4915 21720 5115 21745
rect 5196 21735 5200 21795
rect 5144 21729 5200 21735
rect 4915 21700 4985 21720
rect 4890 21660 4985 21700
rect 5045 21700 5115 21720
rect 5045 21660 5140 21700
rect 4890 21610 5140 21660
rect 4890 21570 4985 21610
rect 4915 21550 4985 21570
rect 5045 21570 5140 21610
rect 5045 21550 5115 21570
rect 4830 21535 4886 21541
rect 4830 21475 4834 21535
rect 4915 21525 5115 21550
rect 5170 21541 5200 21729
rect 5144 21535 5200 21541
rect 4886 21475 5144 21495
rect 5196 21475 5200 21535
rect 4830 21465 5200 21475
rect 5230 21795 5600 21805
rect 5230 21735 5234 21795
rect 5286 21775 5544 21795
rect 5230 21729 5286 21735
rect 5230 21541 5260 21729
rect 5315 21720 5515 21745
rect 5596 21735 5600 21795
rect 5544 21729 5600 21735
rect 5315 21700 5385 21720
rect 5290 21660 5385 21700
rect 5445 21700 5515 21720
rect 5445 21660 5540 21700
rect 5290 21610 5540 21660
rect 5290 21570 5385 21610
rect 5315 21550 5385 21570
rect 5445 21570 5540 21610
rect 5445 21550 5515 21570
rect 5230 21535 5286 21541
rect 5230 21475 5234 21535
rect 5315 21525 5515 21550
rect 5570 21541 5600 21729
rect 5544 21535 5600 21541
rect 5286 21475 5544 21495
rect 5596 21475 5600 21535
rect 5230 21465 5600 21475
rect 5630 21795 6000 21805
rect 5630 21735 5634 21795
rect 5686 21775 5944 21795
rect 5630 21729 5686 21735
rect 5630 21541 5660 21729
rect 5715 21720 5915 21745
rect 5996 21735 6000 21795
rect 5944 21729 6000 21735
rect 5715 21700 5785 21720
rect 5690 21660 5785 21700
rect 5845 21700 5915 21720
rect 5845 21660 5940 21700
rect 5690 21610 5940 21660
rect 5690 21570 5785 21610
rect 5715 21550 5785 21570
rect 5845 21570 5940 21610
rect 5845 21550 5915 21570
rect 5630 21535 5686 21541
rect 5630 21475 5634 21535
rect 5715 21525 5915 21550
rect 5970 21541 6000 21729
rect 5944 21535 6000 21541
rect 5686 21475 5944 21495
rect 5996 21475 6000 21535
rect 5630 21465 6000 21475
rect 6030 21795 6400 21805
rect 6030 21735 6034 21795
rect 6086 21775 6344 21795
rect 6030 21729 6086 21735
rect 6030 21541 6060 21729
rect 6115 21720 6315 21745
rect 6396 21735 6400 21795
rect 6344 21729 6400 21735
rect 6115 21700 6185 21720
rect 6090 21660 6185 21700
rect 6245 21700 6315 21720
rect 6245 21660 6340 21700
rect 6090 21610 6340 21660
rect 6090 21570 6185 21610
rect 6115 21550 6185 21570
rect 6245 21570 6340 21610
rect 6245 21550 6315 21570
rect 6030 21535 6086 21541
rect 6030 21475 6034 21535
rect 6115 21525 6315 21550
rect 6370 21541 6400 21729
rect 6344 21535 6400 21541
rect 6086 21475 6344 21495
rect 6396 21475 6400 21535
rect 6030 21465 6400 21475
rect 6430 21795 6800 21805
rect 6430 21735 6434 21795
rect 6486 21775 6744 21795
rect 6430 21729 6486 21735
rect 6430 21541 6460 21729
rect 6515 21720 6715 21745
rect 6796 21735 6800 21795
rect 6744 21729 6800 21735
rect 6515 21700 6585 21720
rect 6490 21660 6585 21700
rect 6645 21700 6715 21720
rect 6645 21660 6740 21700
rect 6490 21610 6740 21660
rect 6490 21570 6585 21610
rect 6515 21550 6585 21570
rect 6645 21570 6740 21610
rect 6645 21550 6715 21570
rect 6430 21535 6486 21541
rect 6430 21475 6434 21535
rect 6515 21525 6715 21550
rect 6770 21541 6800 21729
rect 6744 21535 6800 21541
rect 6486 21475 6744 21495
rect 6796 21475 6800 21535
rect 6430 21465 6800 21475
rect 6830 21795 7200 21805
rect 6830 21735 6834 21795
rect 6886 21775 7144 21795
rect 6830 21729 6886 21735
rect 6830 21541 6860 21729
rect 6915 21720 7115 21745
rect 7196 21735 7200 21795
rect 7144 21729 7200 21735
rect 6915 21700 6985 21720
rect 6890 21660 6985 21700
rect 7045 21700 7115 21720
rect 7045 21660 7140 21700
rect 6890 21610 7140 21660
rect 6890 21570 6985 21610
rect 6915 21550 6985 21570
rect 7045 21570 7140 21610
rect 7045 21550 7115 21570
rect 6830 21535 6886 21541
rect 6830 21475 6834 21535
rect 6915 21525 7115 21550
rect 7170 21541 7200 21729
rect 7144 21535 7200 21541
rect 6886 21475 7144 21495
rect 7196 21475 7200 21535
rect 6830 21465 7200 21475
rect 7230 21795 7600 21805
rect 7230 21735 7234 21795
rect 7286 21775 7544 21795
rect 7230 21729 7286 21735
rect 7230 21541 7260 21729
rect 7315 21720 7515 21745
rect 7596 21735 7600 21795
rect 7544 21729 7600 21735
rect 7315 21700 7385 21720
rect 7290 21660 7385 21700
rect 7445 21700 7515 21720
rect 7445 21660 7540 21700
rect 7290 21610 7540 21660
rect 7290 21570 7385 21610
rect 7315 21550 7385 21570
rect 7445 21570 7540 21610
rect 7445 21550 7515 21570
rect 7230 21535 7286 21541
rect 7230 21475 7234 21535
rect 7315 21525 7515 21550
rect 7570 21541 7600 21729
rect 7544 21535 7600 21541
rect 7286 21475 7544 21495
rect 7596 21475 7600 21535
rect 7230 21465 7600 21475
rect 7630 21795 8000 21805
rect 7630 21735 7634 21795
rect 7686 21775 7944 21795
rect 7630 21729 7686 21735
rect 7630 21541 7660 21729
rect 7715 21720 7915 21745
rect 7996 21735 8000 21795
rect 7944 21729 8000 21735
rect 7715 21700 7785 21720
rect 7690 21660 7785 21700
rect 7845 21700 7915 21720
rect 7845 21660 7940 21700
rect 7690 21610 7940 21660
rect 7690 21570 7785 21610
rect 7715 21550 7785 21570
rect 7845 21570 7940 21610
rect 7845 21550 7915 21570
rect 7630 21535 7686 21541
rect 7630 21475 7634 21535
rect 7715 21525 7915 21550
rect 7970 21541 8000 21729
rect 7944 21535 8000 21541
rect 7686 21475 7944 21495
rect 7996 21475 8000 21535
rect 7630 21465 8000 21475
rect 8030 21795 8400 21805
rect 8030 21735 8034 21795
rect 8086 21775 8344 21795
rect 8030 21729 8086 21735
rect 8030 21541 8060 21729
rect 8115 21720 8315 21745
rect 8396 21735 8400 21795
rect 8344 21729 8400 21735
rect 8115 21700 8185 21720
rect 8090 21660 8185 21700
rect 8245 21700 8315 21720
rect 8245 21660 8340 21700
rect 8090 21610 8340 21660
rect 8090 21570 8185 21610
rect 8115 21550 8185 21570
rect 8245 21570 8340 21610
rect 8245 21550 8315 21570
rect 8030 21535 8086 21541
rect 8030 21475 8034 21535
rect 8115 21525 8315 21550
rect 8370 21541 8400 21729
rect 8344 21535 8400 21541
rect 8086 21475 8344 21495
rect 8396 21475 8400 21535
rect 8030 21465 8400 21475
rect 8430 21795 8800 21805
rect 8430 21735 8434 21795
rect 8486 21775 8744 21795
rect 8430 21729 8486 21735
rect 8430 21541 8460 21729
rect 8515 21720 8715 21745
rect 8796 21735 8800 21795
rect 8744 21729 8800 21735
rect 8515 21700 8585 21720
rect 8490 21660 8585 21700
rect 8645 21700 8715 21720
rect 8645 21660 8740 21700
rect 8490 21610 8740 21660
rect 8490 21570 8585 21610
rect 8515 21550 8585 21570
rect 8645 21570 8740 21610
rect 8645 21550 8715 21570
rect 8430 21535 8486 21541
rect 8430 21475 8434 21535
rect 8515 21525 8715 21550
rect 8770 21541 8800 21729
rect 8744 21535 8800 21541
rect 8486 21475 8744 21495
rect 8796 21475 8800 21535
rect 8430 21465 8800 21475
rect 8830 21795 9200 21805
rect 8830 21735 8834 21795
rect 8886 21775 9144 21795
rect 8830 21729 8886 21735
rect 8830 21541 8860 21729
rect 8915 21720 9115 21745
rect 9196 21735 9200 21795
rect 9144 21729 9200 21735
rect 8915 21700 8985 21720
rect 8890 21660 8985 21700
rect 9045 21700 9115 21720
rect 9045 21660 9140 21700
rect 8890 21610 9140 21660
rect 8890 21570 8985 21610
rect 8915 21550 8985 21570
rect 9045 21570 9140 21610
rect 9045 21550 9115 21570
rect 8830 21535 8886 21541
rect 8830 21475 8834 21535
rect 8915 21525 9115 21550
rect 9170 21541 9200 21729
rect 9144 21535 9200 21541
rect 8886 21475 9144 21495
rect 9196 21475 9200 21535
rect 8830 21465 9200 21475
rect 9230 21795 9600 21805
rect 9230 21735 9234 21795
rect 9286 21775 9544 21795
rect 9230 21729 9286 21735
rect 9230 21541 9260 21729
rect 9315 21720 9515 21745
rect 9596 21735 9600 21795
rect 9544 21729 9600 21735
rect 9315 21700 9385 21720
rect 9290 21660 9385 21700
rect 9445 21700 9515 21720
rect 9445 21660 9540 21700
rect 9290 21610 9540 21660
rect 9290 21570 9385 21610
rect 9315 21550 9385 21570
rect 9445 21570 9540 21610
rect 9445 21550 9515 21570
rect 9230 21535 9286 21541
rect 9230 21475 9234 21535
rect 9315 21525 9515 21550
rect 9570 21541 9600 21729
rect 9544 21535 9600 21541
rect 9286 21475 9544 21495
rect 9596 21475 9600 21535
rect 9230 21465 9600 21475
rect 9630 21795 10000 21805
rect 9630 21735 9634 21795
rect 9686 21775 9944 21795
rect 9630 21729 9686 21735
rect 9630 21541 9660 21729
rect 9715 21720 9915 21745
rect 9996 21735 10000 21795
rect 9944 21729 10000 21735
rect 9715 21700 9785 21720
rect 9690 21660 9785 21700
rect 9845 21700 9915 21720
rect 9845 21660 9940 21700
rect 9690 21610 9940 21660
rect 9690 21570 9785 21610
rect 9715 21550 9785 21570
rect 9845 21570 9940 21610
rect 9845 21550 9915 21570
rect 9630 21535 9686 21541
rect 9630 21475 9634 21535
rect 9715 21525 9915 21550
rect 9970 21541 10000 21729
rect 9944 21535 10000 21541
rect 9686 21475 9944 21495
rect 9996 21475 10000 21535
rect 9630 21465 10000 21475
rect 10030 21795 10400 21805
rect 10030 21735 10034 21795
rect 10086 21775 10344 21795
rect 10030 21729 10086 21735
rect 10030 21541 10060 21729
rect 10115 21720 10315 21745
rect 10396 21735 10400 21795
rect 10344 21729 10400 21735
rect 10115 21700 10185 21720
rect 10090 21660 10185 21700
rect 10245 21700 10315 21720
rect 10245 21660 10340 21700
rect 10090 21610 10340 21660
rect 10090 21570 10185 21610
rect 10115 21550 10185 21570
rect 10245 21570 10340 21610
rect 10245 21550 10315 21570
rect 10030 21535 10086 21541
rect 10030 21475 10034 21535
rect 10115 21525 10315 21550
rect 10370 21541 10400 21729
rect 10344 21535 10400 21541
rect 10086 21475 10344 21495
rect 10396 21475 10400 21535
rect 10030 21465 10400 21475
rect 10430 21795 10800 21805
rect 10430 21735 10434 21795
rect 10486 21775 10744 21795
rect 10430 21729 10486 21735
rect 10430 21541 10460 21729
rect 10515 21720 10715 21745
rect 10796 21735 10800 21795
rect 10744 21729 10800 21735
rect 10515 21700 10585 21720
rect 10490 21660 10585 21700
rect 10645 21700 10715 21720
rect 10645 21660 10740 21700
rect 10490 21610 10740 21660
rect 10490 21570 10585 21610
rect 10515 21550 10585 21570
rect 10645 21570 10740 21610
rect 10645 21550 10715 21570
rect 10430 21535 10486 21541
rect 10430 21475 10434 21535
rect 10515 21525 10715 21550
rect 10770 21541 10800 21729
rect 10744 21535 10800 21541
rect 10486 21475 10744 21495
rect 10796 21475 10800 21535
rect 10430 21465 10800 21475
rect 10830 21795 11200 21805
rect 10830 21735 10834 21795
rect 10886 21775 11144 21795
rect 10830 21729 10886 21735
rect 10830 21541 10860 21729
rect 10915 21720 11115 21745
rect 11196 21735 11200 21795
rect 11144 21729 11200 21735
rect 10915 21700 10985 21720
rect 10890 21660 10985 21700
rect 11045 21700 11115 21720
rect 11045 21660 11140 21700
rect 10890 21610 11140 21660
rect 10890 21570 10985 21610
rect 10915 21550 10985 21570
rect 11045 21570 11140 21610
rect 11045 21550 11115 21570
rect 10830 21535 10886 21541
rect 10830 21475 10834 21535
rect 10915 21525 11115 21550
rect 11170 21541 11200 21729
rect 11144 21535 11200 21541
rect 10886 21475 11144 21495
rect 11196 21475 11200 21535
rect 10830 21465 11200 21475
rect 11230 21795 11600 21805
rect 11230 21735 11234 21795
rect 11286 21775 11544 21795
rect 11230 21729 11286 21735
rect 11230 21541 11260 21729
rect 11315 21720 11515 21745
rect 11596 21735 11600 21795
rect 11544 21729 11600 21735
rect 11315 21700 11385 21720
rect 11290 21660 11385 21700
rect 11445 21700 11515 21720
rect 11445 21660 11540 21700
rect 11290 21610 11540 21660
rect 11290 21570 11385 21610
rect 11315 21550 11385 21570
rect 11445 21570 11540 21610
rect 11445 21550 11515 21570
rect 11230 21535 11286 21541
rect 11230 21475 11234 21535
rect 11315 21525 11515 21550
rect 11570 21541 11600 21729
rect 11544 21535 11600 21541
rect 11286 21475 11544 21495
rect 11596 21475 11600 21535
rect 11230 21465 11600 21475
rect 11630 21795 12000 21805
rect 11630 21735 11634 21795
rect 11686 21775 11944 21795
rect 11630 21729 11686 21735
rect 11630 21541 11660 21729
rect 11715 21720 11915 21745
rect 11996 21735 12000 21795
rect 11944 21729 12000 21735
rect 11715 21700 11785 21720
rect 11690 21660 11785 21700
rect 11845 21700 11915 21720
rect 11845 21660 11940 21700
rect 11690 21610 11940 21660
rect 11690 21570 11785 21610
rect 11715 21550 11785 21570
rect 11845 21570 11940 21610
rect 11845 21550 11915 21570
rect 11630 21535 11686 21541
rect 11630 21475 11634 21535
rect 11715 21525 11915 21550
rect 11970 21541 12000 21729
rect 11944 21535 12000 21541
rect 11686 21475 11944 21495
rect 11996 21475 12000 21535
rect 11630 21465 12000 21475
rect 12030 21795 12400 21805
rect 12030 21735 12034 21795
rect 12086 21775 12344 21795
rect 12030 21729 12086 21735
rect 12030 21541 12060 21729
rect 12115 21720 12315 21745
rect 12396 21735 12400 21795
rect 12344 21729 12400 21735
rect 12115 21700 12185 21720
rect 12090 21660 12185 21700
rect 12245 21700 12315 21720
rect 12245 21660 12340 21700
rect 12090 21610 12340 21660
rect 12090 21570 12185 21610
rect 12115 21550 12185 21570
rect 12245 21570 12340 21610
rect 12245 21550 12315 21570
rect 12030 21535 12086 21541
rect 12030 21475 12034 21535
rect 12115 21525 12315 21550
rect 12370 21541 12400 21729
rect 12344 21535 12400 21541
rect 12086 21475 12344 21495
rect 12396 21475 12400 21535
rect 12030 21465 12400 21475
rect 12430 21795 12800 21805
rect 12430 21735 12434 21795
rect 12486 21775 12744 21795
rect 12430 21729 12486 21735
rect 12430 21541 12460 21729
rect 12515 21720 12715 21745
rect 12796 21735 12800 21795
rect 12744 21729 12800 21735
rect 12515 21700 12585 21720
rect 12490 21660 12585 21700
rect 12645 21700 12715 21720
rect 12645 21660 12740 21700
rect 12490 21610 12740 21660
rect 12490 21570 12585 21610
rect 12515 21550 12585 21570
rect 12645 21570 12740 21610
rect 12645 21550 12715 21570
rect 12430 21535 12486 21541
rect 12430 21475 12434 21535
rect 12515 21525 12715 21550
rect 12770 21541 12800 21729
rect 12744 21535 12800 21541
rect 12486 21475 12744 21495
rect 12796 21475 12800 21535
rect 12430 21465 12800 21475
rect 12830 21795 13200 21805
rect 12830 21735 12834 21795
rect 12886 21775 13144 21795
rect 12830 21729 12886 21735
rect 12830 21541 12860 21729
rect 12915 21720 13115 21745
rect 13196 21735 13200 21795
rect 13144 21729 13200 21735
rect 12915 21700 12985 21720
rect 12890 21660 12985 21700
rect 13045 21700 13115 21720
rect 13045 21660 13140 21700
rect 12890 21610 13140 21660
rect 12890 21570 12985 21610
rect 12915 21550 12985 21570
rect 13045 21570 13140 21610
rect 13045 21550 13115 21570
rect 12830 21535 12886 21541
rect 12830 21475 12834 21535
rect 12915 21525 13115 21550
rect 13170 21541 13200 21729
rect 13144 21535 13200 21541
rect 12886 21475 13144 21495
rect 13196 21475 13200 21535
rect 12830 21465 13200 21475
rect -370 21425 0 21435
rect -370 21365 -366 21425
rect -314 21405 -56 21425
rect -370 21359 -314 21365
rect -370 21171 -340 21359
rect -285 21350 -85 21375
rect -4 21365 0 21425
rect -56 21359 0 21365
rect -285 21330 -215 21350
rect -310 21290 -215 21330
rect -155 21330 -85 21350
rect -155 21290 -60 21330
rect -310 21240 -60 21290
rect -310 21200 -215 21240
rect -285 21180 -215 21200
rect -155 21200 -60 21240
rect -155 21180 -85 21200
rect -370 21165 -314 21171
rect -370 21105 -366 21165
rect -285 21155 -85 21180
rect -30 21171 0 21359
rect -56 21165 0 21171
rect -314 21105 -56 21125
rect -4 21105 0 21165
rect -370 21095 0 21105
rect 30 21425 400 21435
rect 30 21365 34 21425
rect 86 21405 344 21425
rect 30 21359 86 21365
rect 30 21171 60 21359
rect 115 21350 315 21375
rect 396 21365 400 21425
rect 344 21359 400 21365
rect 115 21330 185 21350
rect 90 21290 185 21330
rect 245 21330 315 21350
rect 245 21290 340 21330
rect 90 21240 340 21290
rect 90 21200 185 21240
rect 115 21180 185 21200
rect 245 21200 340 21240
rect 245 21180 315 21200
rect 30 21165 86 21171
rect 30 21105 34 21165
rect 115 21155 315 21180
rect 370 21171 400 21359
rect 344 21165 400 21171
rect 86 21105 344 21125
rect 396 21105 400 21165
rect 30 21095 400 21105
rect 430 21425 800 21435
rect 430 21365 434 21425
rect 486 21405 744 21425
rect 430 21359 486 21365
rect 430 21171 460 21359
rect 515 21350 715 21375
rect 796 21365 800 21425
rect 744 21359 800 21365
rect 515 21330 585 21350
rect 490 21290 585 21330
rect 645 21330 715 21350
rect 645 21290 740 21330
rect 490 21240 740 21290
rect 490 21200 585 21240
rect 515 21180 585 21200
rect 645 21200 740 21240
rect 645 21180 715 21200
rect 430 21165 486 21171
rect 430 21105 434 21165
rect 515 21155 715 21180
rect 770 21171 800 21359
rect 744 21165 800 21171
rect 486 21105 744 21125
rect 796 21105 800 21165
rect 430 21095 800 21105
rect 830 21425 1200 21435
rect 830 21365 834 21425
rect 886 21405 1144 21425
rect 830 21359 886 21365
rect 830 21171 860 21359
rect 915 21350 1115 21375
rect 1196 21365 1200 21425
rect 1144 21359 1200 21365
rect 915 21330 985 21350
rect 890 21290 985 21330
rect 1045 21330 1115 21350
rect 1045 21290 1140 21330
rect 890 21240 1140 21290
rect 890 21200 985 21240
rect 915 21180 985 21200
rect 1045 21200 1140 21240
rect 1045 21180 1115 21200
rect 830 21165 886 21171
rect 830 21105 834 21165
rect 915 21155 1115 21180
rect 1170 21171 1200 21359
rect 1144 21165 1200 21171
rect 886 21105 1144 21125
rect 1196 21105 1200 21165
rect 830 21095 1200 21105
rect 1230 21425 1600 21435
rect 1230 21365 1234 21425
rect 1286 21405 1544 21425
rect 1230 21359 1286 21365
rect 1230 21171 1260 21359
rect 1315 21350 1515 21375
rect 1596 21365 1600 21425
rect 1544 21359 1600 21365
rect 1315 21330 1385 21350
rect 1290 21290 1385 21330
rect 1445 21330 1515 21350
rect 1445 21290 1540 21330
rect 1290 21240 1540 21290
rect 1290 21200 1385 21240
rect 1315 21180 1385 21200
rect 1445 21200 1540 21240
rect 1445 21180 1515 21200
rect 1230 21165 1286 21171
rect 1230 21105 1234 21165
rect 1315 21155 1515 21180
rect 1570 21171 1600 21359
rect 1544 21165 1600 21171
rect 1286 21105 1544 21125
rect 1596 21105 1600 21165
rect 1230 21095 1600 21105
rect 1630 21425 2000 21435
rect 1630 21365 1634 21425
rect 1686 21405 1944 21425
rect 1630 21359 1686 21365
rect 1630 21171 1660 21359
rect 1715 21350 1915 21375
rect 1996 21365 2000 21425
rect 1944 21359 2000 21365
rect 1715 21330 1785 21350
rect 1690 21290 1785 21330
rect 1845 21330 1915 21350
rect 1845 21290 1940 21330
rect 1690 21240 1940 21290
rect 1690 21200 1785 21240
rect 1715 21180 1785 21200
rect 1845 21200 1940 21240
rect 1845 21180 1915 21200
rect 1630 21165 1686 21171
rect 1630 21105 1634 21165
rect 1715 21155 1915 21180
rect 1970 21171 2000 21359
rect 1944 21165 2000 21171
rect 1686 21105 1944 21125
rect 1996 21105 2000 21165
rect 1630 21095 2000 21105
rect 2030 21425 2400 21435
rect 2030 21365 2034 21425
rect 2086 21405 2344 21425
rect 2030 21359 2086 21365
rect 2030 21171 2060 21359
rect 2115 21350 2315 21375
rect 2396 21365 2400 21425
rect 2344 21359 2400 21365
rect 2115 21330 2185 21350
rect 2090 21290 2185 21330
rect 2245 21330 2315 21350
rect 2245 21290 2340 21330
rect 2090 21240 2340 21290
rect 2090 21200 2185 21240
rect 2115 21180 2185 21200
rect 2245 21200 2340 21240
rect 2245 21180 2315 21200
rect 2030 21165 2086 21171
rect 2030 21105 2034 21165
rect 2115 21155 2315 21180
rect 2370 21171 2400 21359
rect 2344 21165 2400 21171
rect 2086 21105 2344 21125
rect 2396 21105 2400 21165
rect 2030 21095 2400 21105
rect 2430 21425 2800 21435
rect 2430 21365 2434 21425
rect 2486 21405 2744 21425
rect 2430 21359 2486 21365
rect 2430 21171 2460 21359
rect 2515 21350 2715 21375
rect 2796 21365 2800 21425
rect 2744 21359 2800 21365
rect 2515 21330 2585 21350
rect 2490 21290 2585 21330
rect 2645 21330 2715 21350
rect 2645 21290 2740 21330
rect 2490 21240 2740 21290
rect 2490 21200 2585 21240
rect 2515 21180 2585 21200
rect 2645 21200 2740 21240
rect 2645 21180 2715 21200
rect 2430 21165 2486 21171
rect 2430 21105 2434 21165
rect 2515 21155 2715 21180
rect 2770 21171 2800 21359
rect 2744 21165 2800 21171
rect 2486 21105 2744 21125
rect 2796 21105 2800 21165
rect 2430 21095 2800 21105
rect 2830 21425 3200 21435
rect 2830 21365 2834 21425
rect 2886 21405 3144 21425
rect 2830 21359 2886 21365
rect 2830 21171 2860 21359
rect 2915 21350 3115 21375
rect 3196 21365 3200 21425
rect 3144 21359 3200 21365
rect 2915 21330 2985 21350
rect 2890 21290 2985 21330
rect 3045 21330 3115 21350
rect 3045 21290 3140 21330
rect 2890 21240 3140 21290
rect 2890 21200 2985 21240
rect 2915 21180 2985 21200
rect 3045 21200 3140 21240
rect 3045 21180 3115 21200
rect 2830 21165 2886 21171
rect 2830 21105 2834 21165
rect 2915 21155 3115 21180
rect 3170 21171 3200 21359
rect 3144 21165 3200 21171
rect 2886 21105 3144 21125
rect 3196 21105 3200 21165
rect 2830 21095 3200 21105
rect 3230 21425 3600 21435
rect 3230 21365 3234 21425
rect 3286 21405 3544 21425
rect 3230 21359 3286 21365
rect 3230 21171 3260 21359
rect 3315 21350 3515 21375
rect 3596 21365 3600 21425
rect 3544 21359 3600 21365
rect 3315 21330 3385 21350
rect 3290 21290 3385 21330
rect 3445 21330 3515 21350
rect 3445 21290 3540 21330
rect 3290 21240 3540 21290
rect 3290 21200 3385 21240
rect 3315 21180 3385 21200
rect 3445 21200 3540 21240
rect 3445 21180 3515 21200
rect 3230 21165 3286 21171
rect 3230 21105 3234 21165
rect 3315 21155 3515 21180
rect 3570 21171 3600 21359
rect 3544 21165 3600 21171
rect 3286 21105 3544 21125
rect 3596 21105 3600 21165
rect 3230 21095 3600 21105
rect 3630 21425 4000 21435
rect 3630 21365 3634 21425
rect 3686 21405 3944 21425
rect 3630 21359 3686 21365
rect 3630 21171 3660 21359
rect 3715 21350 3915 21375
rect 3996 21365 4000 21425
rect 3944 21359 4000 21365
rect 3715 21330 3785 21350
rect 3690 21290 3785 21330
rect 3845 21330 3915 21350
rect 3845 21290 3940 21330
rect 3690 21240 3940 21290
rect 3690 21200 3785 21240
rect 3715 21180 3785 21200
rect 3845 21200 3940 21240
rect 3845 21180 3915 21200
rect 3630 21165 3686 21171
rect 3630 21105 3634 21165
rect 3715 21155 3915 21180
rect 3970 21171 4000 21359
rect 3944 21165 4000 21171
rect 3686 21105 3944 21125
rect 3996 21105 4000 21165
rect 3630 21095 4000 21105
rect 4030 21425 4400 21435
rect 4030 21365 4034 21425
rect 4086 21405 4344 21425
rect 4030 21359 4086 21365
rect 4030 21171 4060 21359
rect 4115 21350 4315 21375
rect 4396 21365 4400 21425
rect 4344 21359 4400 21365
rect 4115 21330 4185 21350
rect 4090 21290 4185 21330
rect 4245 21330 4315 21350
rect 4245 21290 4340 21330
rect 4090 21240 4340 21290
rect 4090 21200 4185 21240
rect 4115 21180 4185 21200
rect 4245 21200 4340 21240
rect 4245 21180 4315 21200
rect 4030 21165 4086 21171
rect 4030 21105 4034 21165
rect 4115 21155 4315 21180
rect 4370 21171 4400 21359
rect 4344 21165 4400 21171
rect 4086 21105 4344 21125
rect 4396 21105 4400 21165
rect 4030 21095 4400 21105
rect 4430 21425 4800 21435
rect 4430 21365 4434 21425
rect 4486 21405 4744 21425
rect 4430 21359 4486 21365
rect 4430 21171 4460 21359
rect 4515 21350 4715 21375
rect 4796 21365 4800 21425
rect 4744 21359 4800 21365
rect 4515 21330 4585 21350
rect 4490 21290 4585 21330
rect 4645 21330 4715 21350
rect 4645 21290 4740 21330
rect 4490 21240 4740 21290
rect 4490 21200 4585 21240
rect 4515 21180 4585 21200
rect 4645 21200 4740 21240
rect 4645 21180 4715 21200
rect 4430 21165 4486 21171
rect 4430 21105 4434 21165
rect 4515 21155 4715 21180
rect 4770 21171 4800 21359
rect 4744 21165 4800 21171
rect 4486 21105 4744 21125
rect 4796 21105 4800 21165
rect 4430 21095 4800 21105
rect 4830 21425 5200 21435
rect 4830 21365 4834 21425
rect 4886 21405 5144 21425
rect 4830 21359 4886 21365
rect 4830 21171 4860 21359
rect 4915 21350 5115 21375
rect 5196 21365 5200 21425
rect 5144 21359 5200 21365
rect 4915 21330 4985 21350
rect 4890 21290 4985 21330
rect 5045 21330 5115 21350
rect 5045 21290 5140 21330
rect 4890 21240 5140 21290
rect 4890 21200 4985 21240
rect 4915 21180 4985 21200
rect 5045 21200 5140 21240
rect 5045 21180 5115 21200
rect 4830 21165 4886 21171
rect 4830 21105 4834 21165
rect 4915 21155 5115 21180
rect 5170 21171 5200 21359
rect 5144 21165 5200 21171
rect 4886 21105 5144 21125
rect 5196 21105 5200 21165
rect 4830 21095 5200 21105
rect 5230 21425 5600 21435
rect 5230 21365 5234 21425
rect 5286 21405 5544 21425
rect 5230 21359 5286 21365
rect 5230 21171 5260 21359
rect 5315 21350 5515 21375
rect 5596 21365 5600 21425
rect 5544 21359 5600 21365
rect 5315 21330 5385 21350
rect 5290 21290 5385 21330
rect 5445 21330 5515 21350
rect 5445 21290 5540 21330
rect 5290 21240 5540 21290
rect 5290 21200 5385 21240
rect 5315 21180 5385 21200
rect 5445 21200 5540 21240
rect 5445 21180 5515 21200
rect 5230 21165 5286 21171
rect 5230 21105 5234 21165
rect 5315 21155 5515 21180
rect 5570 21171 5600 21359
rect 5544 21165 5600 21171
rect 5286 21105 5544 21125
rect 5596 21105 5600 21165
rect 5230 21095 5600 21105
rect 5630 21425 6000 21435
rect 5630 21365 5634 21425
rect 5686 21405 5944 21425
rect 5630 21359 5686 21365
rect 5630 21171 5660 21359
rect 5715 21350 5915 21375
rect 5996 21365 6000 21425
rect 5944 21359 6000 21365
rect 5715 21330 5785 21350
rect 5690 21290 5785 21330
rect 5845 21330 5915 21350
rect 5845 21290 5940 21330
rect 5690 21240 5940 21290
rect 5690 21200 5785 21240
rect 5715 21180 5785 21200
rect 5845 21200 5940 21240
rect 5845 21180 5915 21200
rect 5630 21165 5686 21171
rect 5630 21105 5634 21165
rect 5715 21155 5915 21180
rect 5970 21171 6000 21359
rect 5944 21165 6000 21171
rect 5686 21105 5944 21125
rect 5996 21105 6000 21165
rect 5630 21095 6000 21105
rect 6030 21425 6400 21435
rect 6030 21365 6034 21425
rect 6086 21405 6344 21425
rect 6030 21359 6086 21365
rect 6030 21171 6060 21359
rect 6115 21350 6315 21375
rect 6396 21365 6400 21425
rect 6344 21359 6400 21365
rect 6115 21330 6185 21350
rect 6090 21290 6185 21330
rect 6245 21330 6315 21350
rect 6245 21290 6340 21330
rect 6090 21240 6340 21290
rect 6090 21200 6185 21240
rect 6115 21180 6185 21200
rect 6245 21200 6340 21240
rect 6245 21180 6315 21200
rect 6030 21165 6086 21171
rect 6030 21105 6034 21165
rect 6115 21155 6315 21180
rect 6370 21171 6400 21359
rect 6344 21165 6400 21171
rect 6086 21105 6344 21125
rect 6396 21105 6400 21165
rect 6030 21095 6400 21105
rect 6430 21425 6800 21435
rect 6430 21365 6434 21425
rect 6486 21405 6744 21425
rect 6430 21359 6486 21365
rect 6430 21171 6460 21359
rect 6515 21350 6715 21375
rect 6796 21365 6800 21425
rect 6744 21359 6800 21365
rect 6515 21330 6585 21350
rect 6490 21290 6585 21330
rect 6645 21330 6715 21350
rect 6645 21290 6740 21330
rect 6490 21240 6740 21290
rect 6490 21200 6585 21240
rect 6515 21180 6585 21200
rect 6645 21200 6740 21240
rect 6645 21180 6715 21200
rect 6430 21165 6486 21171
rect 6430 21105 6434 21165
rect 6515 21155 6715 21180
rect 6770 21171 6800 21359
rect 6744 21165 6800 21171
rect 6486 21105 6744 21125
rect 6796 21105 6800 21165
rect 6430 21095 6800 21105
rect 6830 21425 7200 21435
rect 6830 21365 6834 21425
rect 6886 21405 7144 21425
rect 6830 21359 6886 21365
rect 6830 21171 6860 21359
rect 6915 21350 7115 21375
rect 7196 21365 7200 21425
rect 7144 21359 7200 21365
rect 6915 21330 6985 21350
rect 6890 21290 6985 21330
rect 7045 21330 7115 21350
rect 7045 21290 7140 21330
rect 6890 21240 7140 21290
rect 6890 21200 6985 21240
rect 6915 21180 6985 21200
rect 7045 21200 7140 21240
rect 7045 21180 7115 21200
rect 6830 21165 6886 21171
rect 6830 21105 6834 21165
rect 6915 21155 7115 21180
rect 7170 21171 7200 21359
rect 7144 21165 7200 21171
rect 6886 21105 7144 21125
rect 7196 21105 7200 21165
rect 6830 21095 7200 21105
rect 7230 21425 7600 21435
rect 7230 21365 7234 21425
rect 7286 21405 7544 21425
rect 7230 21359 7286 21365
rect 7230 21171 7260 21359
rect 7315 21350 7515 21375
rect 7596 21365 7600 21425
rect 7544 21359 7600 21365
rect 7315 21330 7385 21350
rect 7290 21290 7385 21330
rect 7445 21330 7515 21350
rect 7445 21290 7540 21330
rect 7290 21240 7540 21290
rect 7290 21200 7385 21240
rect 7315 21180 7385 21200
rect 7445 21200 7540 21240
rect 7445 21180 7515 21200
rect 7230 21165 7286 21171
rect 7230 21105 7234 21165
rect 7315 21155 7515 21180
rect 7570 21171 7600 21359
rect 7544 21165 7600 21171
rect 7286 21105 7544 21125
rect 7596 21105 7600 21165
rect 7230 21095 7600 21105
rect 7630 21425 8000 21435
rect 7630 21365 7634 21425
rect 7686 21405 7944 21425
rect 7630 21359 7686 21365
rect 7630 21171 7660 21359
rect 7715 21350 7915 21375
rect 7996 21365 8000 21425
rect 7944 21359 8000 21365
rect 7715 21330 7785 21350
rect 7690 21290 7785 21330
rect 7845 21330 7915 21350
rect 7845 21290 7940 21330
rect 7690 21240 7940 21290
rect 7690 21200 7785 21240
rect 7715 21180 7785 21200
rect 7845 21200 7940 21240
rect 7845 21180 7915 21200
rect 7630 21165 7686 21171
rect 7630 21105 7634 21165
rect 7715 21155 7915 21180
rect 7970 21171 8000 21359
rect 7944 21165 8000 21171
rect 7686 21105 7944 21125
rect 7996 21105 8000 21165
rect 7630 21095 8000 21105
rect 8030 21425 8400 21435
rect 8030 21365 8034 21425
rect 8086 21405 8344 21425
rect 8030 21359 8086 21365
rect 8030 21171 8060 21359
rect 8115 21350 8315 21375
rect 8396 21365 8400 21425
rect 8344 21359 8400 21365
rect 8115 21330 8185 21350
rect 8090 21290 8185 21330
rect 8245 21330 8315 21350
rect 8245 21290 8340 21330
rect 8090 21240 8340 21290
rect 8090 21200 8185 21240
rect 8115 21180 8185 21200
rect 8245 21200 8340 21240
rect 8245 21180 8315 21200
rect 8030 21165 8086 21171
rect 8030 21105 8034 21165
rect 8115 21155 8315 21180
rect 8370 21171 8400 21359
rect 8344 21165 8400 21171
rect 8086 21105 8344 21125
rect 8396 21105 8400 21165
rect 8030 21095 8400 21105
rect 8430 21425 8800 21435
rect 8430 21365 8434 21425
rect 8486 21405 8744 21425
rect 8430 21359 8486 21365
rect 8430 21171 8460 21359
rect 8515 21350 8715 21375
rect 8796 21365 8800 21425
rect 8744 21359 8800 21365
rect 8515 21330 8585 21350
rect 8490 21290 8585 21330
rect 8645 21330 8715 21350
rect 8645 21290 8740 21330
rect 8490 21240 8740 21290
rect 8490 21200 8585 21240
rect 8515 21180 8585 21200
rect 8645 21200 8740 21240
rect 8645 21180 8715 21200
rect 8430 21165 8486 21171
rect 8430 21105 8434 21165
rect 8515 21155 8715 21180
rect 8770 21171 8800 21359
rect 8744 21165 8800 21171
rect 8486 21105 8744 21125
rect 8796 21105 8800 21165
rect 8430 21095 8800 21105
rect 8830 21425 9200 21435
rect 8830 21365 8834 21425
rect 8886 21405 9144 21425
rect 8830 21359 8886 21365
rect 8830 21171 8860 21359
rect 8915 21350 9115 21375
rect 9196 21365 9200 21425
rect 9144 21359 9200 21365
rect 8915 21330 8985 21350
rect 8890 21290 8985 21330
rect 9045 21330 9115 21350
rect 9045 21290 9140 21330
rect 8890 21240 9140 21290
rect 8890 21200 8985 21240
rect 8915 21180 8985 21200
rect 9045 21200 9140 21240
rect 9045 21180 9115 21200
rect 8830 21165 8886 21171
rect 8830 21105 8834 21165
rect 8915 21155 9115 21180
rect 9170 21171 9200 21359
rect 9144 21165 9200 21171
rect 8886 21105 9144 21125
rect 9196 21105 9200 21165
rect 8830 21095 9200 21105
rect 9230 21425 9600 21435
rect 9230 21365 9234 21425
rect 9286 21405 9544 21425
rect 9230 21359 9286 21365
rect 9230 21171 9260 21359
rect 9315 21350 9515 21375
rect 9596 21365 9600 21425
rect 9544 21359 9600 21365
rect 9315 21330 9385 21350
rect 9290 21290 9385 21330
rect 9445 21330 9515 21350
rect 9445 21290 9540 21330
rect 9290 21240 9540 21290
rect 9290 21200 9385 21240
rect 9315 21180 9385 21200
rect 9445 21200 9540 21240
rect 9445 21180 9515 21200
rect 9230 21165 9286 21171
rect 9230 21105 9234 21165
rect 9315 21155 9515 21180
rect 9570 21171 9600 21359
rect 9544 21165 9600 21171
rect 9286 21105 9544 21125
rect 9596 21105 9600 21165
rect 9230 21095 9600 21105
rect 9630 21425 10000 21435
rect 9630 21365 9634 21425
rect 9686 21405 9944 21425
rect 9630 21359 9686 21365
rect 9630 21171 9660 21359
rect 9715 21350 9915 21375
rect 9996 21365 10000 21425
rect 9944 21359 10000 21365
rect 9715 21330 9785 21350
rect 9690 21290 9785 21330
rect 9845 21330 9915 21350
rect 9845 21290 9940 21330
rect 9690 21240 9940 21290
rect 9690 21200 9785 21240
rect 9715 21180 9785 21200
rect 9845 21200 9940 21240
rect 9845 21180 9915 21200
rect 9630 21165 9686 21171
rect 9630 21105 9634 21165
rect 9715 21155 9915 21180
rect 9970 21171 10000 21359
rect 9944 21165 10000 21171
rect 9686 21105 9944 21125
rect 9996 21105 10000 21165
rect 9630 21095 10000 21105
rect 10030 21425 10400 21435
rect 10030 21365 10034 21425
rect 10086 21405 10344 21425
rect 10030 21359 10086 21365
rect 10030 21171 10060 21359
rect 10115 21350 10315 21375
rect 10396 21365 10400 21425
rect 10344 21359 10400 21365
rect 10115 21330 10185 21350
rect 10090 21290 10185 21330
rect 10245 21330 10315 21350
rect 10245 21290 10340 21330
rect 10090 21240 10340 21290
rect 10090 21200 10185 21240
rect 10115 21180 10185 21200
rect 10245 21200 10340 21240
rect 10245 21180 10315 21200
rect 10030 21165 10086 21171
rect 10030 21105 10034 21165
rect 10115 21155 10315 21180
rect 10370 21171 10400 21359
rect 10344 21165 10400 21171
rect 10086 21105 10344 21125
rect 10396 21105 10400 21165
rect 10030 21095 10400 21105
rect 10430 21425 10800 21435
rect 10430 21365 10434 21425
rect 10486 21405 10744 21425
rect 10430 21359 10486 21365
rect 10430 21171 10460 21359
rect 10515 21350 10715 21375
rect 10796 21365 10800 21425
rect 10744 21359 10800 21365
rect 10515 21330 10585 21350
rect 10490 21290 10585 21330
rect 10645 21330 10715 21350
rect 10645 21290 10740 21330
rect 10490 21240 10740 21290
rect 10490 21200 10585 21240
rect 10515 21180 10585 21200
rect 10645 21200 10740 21240
rect 10645 21180 10715 21200
rect 10430 21165 10486 21171
rect 10430 21105 10434 21165
rect 10515 21155 10715 21180
rect 10770 21171 10800 21359
rect 10744 21165 10800 21171
rect 10486 21105 10744 21125
rect 10796 21105 10800 21165
rect 10430 21095 10800 21105
rect 10830 21425 11200 21435
rect 10830 21365 10834 21425
rect 10886 21405 11144 21425
rect 10830 21359 10886 21365
rect 10830 21171 10860 21359
rect 10915 21350 11115 21375
rect 11196 21365 11200 21425
rect 11144 21359 11200 21365
rect 10915 21330 10985 21350
rect 10890 21290 10985 21330
rect 11045 21330 11115 21350
rect 11045 21290 11140 21330
rect 10890 21240 11140 21290
rect 10890 21200 10985 21240
rect 10915 21180 10985 21200
rect 11045 21200 11140 21240
rect 11045 21180 11115 21200
rect 10830 21165 10886 21171
rect 10830 21105 10834 21165
rect 10915 21155 11115 21180
rect 11170 21171 11200 21359
rect 11144 21165 11200 21171
rect 10886 21105 11144 21125
rect 11196 21105 11200 21165
rect 10830 21095 11200 21105
rect 11230 21425 11600 21435
rect 11230 21365 11234 21425
rect 11286 21405 11544 21425
rect 11230 21359 11286 21365
rect 11230 21171 11260 21359
rect 11315 21350 11515 21375
rect 11596 21365 11600 21425
rect 11544 21359 11600 21365
rect 11315 21330 11385 21350
rect 11290 21290 11385 21330
rect 11445 21330 11515 21350
rect 11445 21290 11540 21330
rect 11290 21240 11540 21290
rect 11290 21200 11385 21240
rect 11315 21180 11385 21200
rect 11445 21200 11540 21240
rect 11445 21180 11515 21200
rect 11230 21165 11286 21171
rect 11230 21105 11234 21165
rect 11315 21155 11515 21180
rect 11570 21171 11600 21359
rect 11544 21165 11600 21171
rect 11286 21105 11544 21125
rect 11596 21105 11600 21165
rect 11230 21095 11600 21105
rect 11630 21425 12000 21435
rect 11630 21365 11634 21425
rect 11686 21405 11944 21425
rect 11630 21359 11686 21365
rect 11630 21171 11660 21359
rect 11715 21350 11915 21375
rect 11996 21365 12000 21425
rect 11944 21359 12000 21365
rect 11715 21330 11785 21350
rect 11690 21290 11785 21330
rect 11845 21330 11915 21350
rect 11845 21290 11940 21330
rect 11690 21240 11940 21290
rect 11690 21200 11785 21240
rect 11715 21180 11785 21200
rect 11845 21200 11940 21240
rect 11845 21180 11915 21200
rect 11630 21165 11686 21171
rect 11630 21105 11634 21165
rect 11715 21155 11915 21180
rect 11970 21171 12000 21359
rect 11944 21165 12000 21171
rect 11686 21105 11944 21125
rect 11996 21105 12000 21165
rect 11630 21095 12000 21105
rect 12030 21425 12400 21435
rect 12030 21365 12034 21425
rect 12086 21405 12344 21425
rect 12030 21359 12086 21365
rect 12030 21171 12060 21359
rect 12115 21350 12315 21375
rect 12396 21365 12400 21425
rect 12344 21359 12400 21365
rect 12115 21330 12185 21350
rect 12090 21290 12185 21330
rect 12245 21330 12315 21350
rect 12245 21290 12340 21330
rect 12090 21240 12340 21290
rect 12090 21200 12185 21240
rect 12115 21180 12185 21200
rect 12245 21200 12340 21240
rect 12245 21180 12315 21200
rect 12030 21165 12086 21171
rect 12030 21105 12034 21165
rect 12115 21155 12315 21180
rect 12370 21171 12400 21359
rect 12344 21165 12400 21171
rect 12086 21105 12344 21125
rect 12396 21105 12400 21165
rect 12030 21095 12400 21105
rect 12430 21425 12800 21435
rect 12430 21365 12434 21425
rect 12486 21405 12744 21425
rect 12430 21359 12486 21365
rect 12430 21171 12460 21359
rect 12515 21350 12715 21375
rect 12796 21365 12800 21425
rect 12744 21359 12800 21365
rect 12515 21330 12585 21350
rect 12490 21290 12585 21330
rect 12645 21330 12715 21350
rect 12645 21290 12740 21330
rect 12490 21240 12740 21290
rect 12490 21200 12585 21240
rect 12515 21180 12585 21200
rect 12645 21200 12740 21240
rect 12645 21180 12715 21200
rect 12430 21165 12486 21171
rect 12430 21105 12434 21165
rect 12515 21155 12715 21180
rect 12770 21171 12800 21359
rect 12744 21165 12800 21171
rect 12486 21105 12744 21125
rect 12796 21105 12800 21165
rect 12430 21095 12800 21105
rect 12830 21425 13200 21435
rect 12830 21365 12834 21425
rect 12886 21405 13144 21425
rect 12830 21359 12886 21365
rect 12830 21171 12860 21359
rect 12915 21350 13115 21375
rect 13196 21365 13200 21425
rect 13144 21359 13200 21365
rect 12915 21330 12985 21350
rect 12890 21290 12985 21330
rect 13045 21330 13115 21350
rect 13045 21290 13140 21330
rect 12890 21240 13140 21290
rect 12890 21200 12985 21240
rect 12915 21180 12985 21200
rect 13045 21200 13140 21240
rect 13045 21180 13115 21200
rect 12830 21165 12886 21171
rect 12830 21105 12834 21165
rect 12915 21155 13115 21180
rect 13170 21171 13200 21359
rect 13144 21165 13200 21171
rect 12886 21105 13144 21125
rect 13196 21105 13200 21165
rect 12830 21095 13200 21105
rect -370 21055 0 21065
rect -370 20995 -366 21055
rect -314 21035 -56 21055
rect -370 20989 -314 20995
rect -370 20801 -340 20989
rect -285 20980 -85 21005
rect -4 20995 0 21055
rect -56 20989 0 20995
rect -285 20960 -215 20980
rect -310 20920 -215 20960
rect -155 20960 -85 20980
rect -155 20920 -60 20960
rect -310 20870 -60 20920
rect -310 20830 -215 20870
rect -285 20810 -215 20830
rect -155 20830 -60 20870
rect -155 20810 -85 20830
rect -370 20795 -314 20801
rect -370 20735 -366 20795
rect -285 20785 -85 20810
rect -30 20801 0 20989
rect -56 20795 0 20801
rect -314 20735 -56 20755
rect -4 20735 0 20795
rect -370 20725 0 20735
rect 30 21055 400 21065
rect 30 20995 34 21055
rect 86 21035 344 21055
rect 30 20989 86 20995
rect 30 20801 60 20989
rect 115 20980 315 21005
rect 396 20995 400 21055
rect 344 20989 400 20995
rect 115 20960 185 20980
rect 90 20920 185 20960
rect 245 20960 315 20980
rect 245 20920 340 20960
rect 90 20870 340 20920
rect 90 20830 185 20870
rect 115 20810 185 20830
rect 245 20830 340 20870
rect 245 20810 315 20830
rect 30 20795 86 20801
rect 30 20735 34 20795
rect 115 20785 315 20810
rect 370 20801 400 20989
rect 344 20795 400 20801
rect 86 20735 344 20755
rect 396 20735 400 20795
rect 30 20725 400 20735
rect 430 21055 800 21065
rect 430 20995 434 21055
rect 486 21035 744 21055
rect 430 20989 486 20995
rect 430 20801 460 20989
rect 515 20980 715 21005
rect 796 20995 800 21055
rect 744 20989 800 20995
rect 515 20960 585 20980
rect 490 20920 585 20960
rect 645 20960 715 20980
rect 645 20920 740 20960
rect 490 20870 740 20920
rect 490 20830 585 20870
rect 515 20810 585 20830
rect 645 20830 740 20870
rect 645 20810 715 20830
rect 430 20795 486 20801
rect 430 20735 434 20795
rect 515 20785 715 20810
rect 770 20801 800 20989
rect 744 20795 800 20801
rect 486 20735 744 20755
rect 796 20735 800 20795
rect 430 20725 800 20735
rect 830 21055 1200 21065
rect 830 20995 834 21055
rect 886 21035 1144 21055
rect 830 20989 886 20995
rect 830 20801 860 20989
rect 915 20980 1115 21005
rect 1196 20995 1200 21055
rect 1144 20989 1200 20995
rect 915 20960 985 20980
rect 890 20920 985 20960
rect 1045 20960 1115 20980
rect 1045 20920 1140 20960
rect 890 20870 1140 20920
rect 890 20830 985 20870
rect 915 20810 985 20830
rect 1045 20830 1140 20870
rect 1045 20810 1115 20830
rect 830 20795 886 20801
rect 830 20735 834 20795
rect 915 20785 1115 20810
rect 1170 20801 1200 20989
rect 1144 20795 1200 20801
rect 886 20735 1144 20755
rect 1196 20735 1200 20795
rect 830 20725 1200 20735
rect 1230 21055 1600 21065
rect 1230 20995 1234 21055
rect 1286 21035 1544 21055
rect 1230 20989 1286 20995
rect 1230 20801 1260 20989
rect 1315 20980 1515 21005
rect 1596 20995 1600 21055
rect 1544 20989 1600 20995
rect 1315 20960 1385 20980
rect 1290 20920 1385 20960
rect 1445 20960 1515 20980
rect 1445 20920 1540 20960
rect 1290 20870 1540 20920
rect 1290 20830 1385 20870
rect 1315 20810 1385 20830
rect 1445 20830 1540 20870
rect 1445 20810 1515 20830
rect 1230 20795 1286 20801
rect 1230 20735 1234 20795
rect 1315 20785 1515 20810
rect 1570 20801 1600 20989
rect 1544 20795 1600 20801
rect 1286 20735 1544 20755
rect 1596 20735 1600 20795
rect 1230 20725 1600 20735
rect 1630 21055 2000 21065
rect 1630 20995 1634 21055
rect 1686 21035 1944 21055
rect 1630 20989 1686 20995
rect 1630 20801 1660 20989
rect 1715 20980 1915 21005
rect 1996 20995 2000 21055
rect 1944 20989 2000 20995
rect 1715 20960 1785 20980
rect 1690 20920 1785 20960
rect 1845 20960 1915 20980
rect 1845 20920 1940 20960
rect 1690 20870 1940 20920
rect 1690 20830 1785 20870
rect 1715 20810 1785 20830
rect 1845 20830 1940 20870
rect 1845 20810 1915 20830
rect 1630 20795 1686 20801
rect 1630 20735 1634 20795
rect 1715 20785 1915 20810
rect 1970 20801 2000 20989
rect 1944 20795 2000 20801
rect 1686 20735 1944 20755
rect 1996 20735 2000 20795
rect 1630 20725 2000 20735
rect 2030 21055 2400 21065
rect 2030 20995 2034 21055
rect 2086 21035 2344 21055
rect 2030 20989 2086 20995
rect 2030 20801 2060 20989
rect 2115 20980 2315 21005
rect 2396 20995 2400 21055
rect 2344 20989 2400 20995
rect 2115 20960 2185 20980
rect 2090 20920 2185 20960
rect 2245 20960 2315 20980
rect 2245 20920 2340 20960
rect 2090 20870 2340 20920
rect 2090 20830 2185 20870
rect 2115 20810 2185 20830
rect 2245 20830 2340 20870
rect 2245 20810 2315 20830
rect 2030 20795 2086 20801
rect 2030 20735 2034 20795
rect 2115 20785 2315 20810
rect 2370 20801 2400 20989
rect 2344 20795 2400 20801
rect 2086 20735 2344 20755
rect 2396 20735 2400 20795
rect 2030 20725 2400 20735
rect 2430 21055 2800 21065
rect 2430 20995 2434 21055
rect 2486 21035 2744 21055
rect 2430 20989 2486 20995
rect 2430 20801 2460 20989
rect 2515 20980 2715 21005
rect 2796 20995 2800 21055
rect 2744 20989 2800 20995
rect 2515 20960 2585 20980
rect 2490 20920 2585 20960
rect 2645 20960 2715 20980
rect 2645 20920 2740 20960
rect 2490 20870 2740 20920
rect 2490 20830 2585 20870
rect 2515 20810 2585 20830
rect 2645 20830 2740 20870
rect 2645 20810 2715 20830
rect 2430 20795 2486 20801
rect 2430 20735 2434 20795
rect 2515 20785 2715 20810
rect 2770 20801 2800 20989
rect 2744 20795 2800 20801
rect 2486 20735 2744 20755
rect 2796 20735 2800 20795
rect 2430 20725 2800 20735
rect 2830 21055 3200 21065
rect 2830 20995 2834 21055
rect 2886 21035 3144 21055
rect 2830 20989 2886 20995
rect 2830 20801 2860 20989
rect 2915 20980 3115 21005
rect 3196 20995 3200 21055
rect 3144 20989 3200 20995
rect 2915 20960 2985 20980
rect 2890 20920 2985 20960
rect 3045 20960 3115 20980
rect 3045 20920 3140 20960
rect 2890 20870 3140 20920
rect 2890 20830 2985 20870
rect 2915 20810 2985 20830
rect 3045 20830 3140 20870
rect 3045 20810 3115 20830
rect 2830 20795 2886 20801
rect 2830 20735 2834 20795
rect 2915 20785 3115 20810
rect 3170 20801 3200 20989
rect 3144 20795 3200 20801
rect 2886 20735 3144 20755
rect 3196 20735 3200 20795
rect 2830 20725 3200 20735
rect 3230 21055 3600 21065
rect 3230 20995 3234 21055
rect 3286 21035 3544 21055
rect 3230 20989 3286 20995
rect 3230 20801 3260 20989
rect 3315 20980 3515 21005
rect 3596 20995 3600 21055
rect 3544 20989 3600 20995
rect 3315 20960 3385 20980
rect 3290 20920 3385 20960
rect 3445 20960 3515 20980
rect 3445 20920 3540 20960
rect 3290 20870 3540 20920
rect 3290 20830 3385 20870
rect 3315 20810 3385 20830
rect 3445 20830 3540 20870
rect 3445 20810 3515 20830
rect 3230 20795 3286 20801
rect 3230 20735 3234 20795
rect 3315 20785 3515 20810
rect 3570 20801 3600 20989
rect 3544 20795 3600 20801
rect 3286 20735 3544 20755
rect 3596 20735 3600 20795
rect 3230 20725 3600 20735
rect 3630 21055 4000 21065
rect 3630 20995 3634 21055
rect 3686 21035 3944 21055
rect 3630 20989 3686 20995
rect 3630 20801 3660 20989
rect 3715 20980 3915 21005
rect 3996 20995 4000 21055
rect 3944 20989 4000 20995
rect 3715 20960 3785 20980
rect 3690 20920 3785 20960
rect 3845 20960 3915 20980
rect 3845 20920 3940 20960
rect 3690 20870 3940 20920
rect 3690 20830 3785 20870
rect 3715 20810 3785 20830
rect 3845 20830 3940 20870
rect 3845 20810 3915 20830
rect 3630 20795 3686 20801
rect 3630 20735 3634 20795
rect 3715 20785 3915 20810
rect 3970 20801 4000 20989
rect 3944 20795 4000 20801
rect 3686 20735 3944 20755
rect 3996 20735 4000 20795
rect 3630 20725 4000 20735
rect 4030 21055 4400 21065
rect 4030 20995 4034 21055
rect 4086 21035 4344 21055
rect 4030 20989 4086 20995
rect 4030 20801 4060 20989
rect 4115 20980 4315 21005
rect 4396 20995 4400 21055
rect 4344 20989 4400 20995
rect 4115 20960 4185 20980
rect 4090 20920 4185 20960
rect 4245 20960 4315 20980
rect 4245 20920 4340 20960
rect 4090 20870 4340 20920
rect 4090 20830 4185 20870
rect 4115 20810 4185 20830
rect 4245 20830 4340 20870
rect 4245 20810 4315 20830
rect 4030 20795 4086 20801
rect 4030 20735 4034 20795
rect 4115 20785 4315 20810
rect 4370 20801 4400 20989
rect 4344 20795 4400 20801
rect 4086 20735 4344 20755
rect 4396 20735 4400 20795
rect 4030 20725 4400 20735
rect 4430 21055 4800 21065
rect 4430 20995 4434 21055
rect 4486 21035 4744 21055
rect 4430 20989 4486 20995
rect 4430 20801 4460 20989
rect 4515 20980 4715 21005
rect 4796 20995 4800 21055
rect 4744 20989 4800 20995
rect 4515 20960 4585 20980
rect 4490 20920 4585 20960
rect 4645 20960 4715 20980
rect 4645 20920 4740 20960
rect 4490 20870 4740 20920
rect 4490 20830 4585 20870
rect 4515 20810 4585 20830
rect 4645 20830 4740 20870
rect 4645 20810 4715 20830
rect 4430 20795 4486 20801
rect 4430 20735 4434 20795
rect 4515 20785 4715 20810
rect 4770 20801 4800 20989
rect 4744 20795 4800 20801
rect 4486 20735 4744 20755
rect 4796 20735 4800 20795
rect 4430 20725 4800 20735
rect 4830 21055 5200 21065
rect 4830 20995 4834 21055
rect 4886 21035 5144 21055
rect 4830 20989 4886 20995
rect 4830 20801 4860 20989
rect 4915 20980 5115 21005
rect 5196 20995 5200 21055
rect 5144 20989 5200 20995
rect 4915 20960 4985 20980
rect 4890 20920 4985 20960
rect 5045 20960 5115 20980
rect 5045 20920 5140 20960
rect 4890 20870 5140 20920
rect 4890 20830 4985 20870
rect 4915 20810 4985 20830
rect 5045 20830 5140 20870
rect 5045 20810 5115 20830
rect 4830 20795 4886 20801
rect 4830 20735 4834 20795
rect 4915 20785 5115 20810
rect 5170 20801 5200 20989
rect 5144 20795 5200 20801
rect 4886 20735 5144 20755
rect 5196 20735 5200 20795
rect 4830 20725 5200 20735
rect 5230 21055 5600 21065
rect 5230 20995 5234 21055
rect 5286 21035 5544 21055
rect 5230 20989 5286 20995
rect 5230 20801 5260 20989
rect 5315 20980 5515 21005
rect 5596 20995 5600 21055
rect 5544 20989 5600 20995
rect 5315 20960 5385 20980
rect 5290 20920 5385 20960
rect 5445 20960 5515 20980
rect 5445 20920 5540 20960
rect 5290 20870 5540 20920
rect 5290 20830 5385 20870
rect 5315 20810 5385 20830
rect 5445 20830 5540 20870
rect 5445 20810 5515 20830
rect 5230 20795 5286 20801
rect 5230 20735 5234 20795
rect 5315 20785 5515 20810
rect 5570 20801 5600 20989
rect 5544 20795 5600 20801
rect 5286 20735 5544 20755
rect 5596 20735 5600 20795
rect 5230 20725 5600 20735
rect 5630 21055 6000 21065
rect 5630 20995 5634 21055
rect 5686 21035 5944 21055
rect 5630 20989 5686 20995
rect 5630 20801 5660 20989
rect 5715 20980 5915 21005
rect 5996 20995 6000 21055
rect 5944 20989 6000 20995
rect 5715 20960 5785 20980
rect 5690 20920 5785 20960
rect 5845 20960 5915 20980
rect 5845 20920 5940 20960
rect 5690 20870 5940 20920
rect 5690 20830 5785 20870
rect 5715 20810 5785 20830
rect 5845 20830 5940 20870
rect 5845 20810 5915 20830
rect 5630 20795 5686 20801
rect 5630 20735 5634 20795
rect 5715 20785 5915 20810
rect 5970 20801 6000 20989
rect 5944 20795 6000 20801
rect 5686 20735 5944 20755
rect 5996 20735 6000 20795
rect 5630 20725 6000 20735
rect 6030 21055 6400 21065
rect 6030 20995 6034 21055
rect 6086 21035 6344 21055
rect 6030 20989 6086 20995
rect 6030 20801 6060 20989
rect 6115 20980 6315 21005
rect 6396 20995 6400 21055
rect 6344 20989 6400 20995
rect 6115 20960 6185 20980
rect 6090 20920 6185 20960
rect 6245 20960 6315 20980
rect 6245 20920 6340 20960
rect 6090 20870 6340 20920
rect 6090 20830 6185 20870
rect 6115 20810 6185 20830
rect 6245 20830 6340 20870
rect 6245 20810 6315 20830
rect 6030 20795 6086 20801
rect 6030 20735 6034 20795
rect 6115 20785 6315 20810
rect 6370 20801 6400 20989
rect 6344 20795 6400 20801
rect 6086 20735 6344 20755
rect 6396 20735 6400 20795
rect 6030 20725 6400 20735
rect 6430 21055 6800 21065
rect 6430 20995 6434 21055
rect 6486 21035 6744 21055
rect 6430 20989 6486 20995
rect 6430 20801 6460 20989
rect 6515 20980 6715 21005
rect 6796 20995 6800 21055
rect 6744 20989 6800 20995
rect 6515 20960 6585 20980
rect 6490 20920 6585 20960
rect 6645 20960 6715 20980
rect 6645 20920 6740 20960
rect 6490 20870 6740 20920
rect 6490 20830 6585 20870
rect 6515 20810 6585 20830
rect 6645 20830 6740 20870
rect 6645 20810 6715 20830
rect 6430 20795 6486 20801
rect 6430 20735 6434 20795
rect 6515 20785 6715 20810
rect 6770 20801 6800 20989
rect 6744 20795 6800 20801
rect 6486 20735 6744 20755
rect 6796 20735 6800 20795
rect 6430 20725 6800 20735
rect 6830 21055 7200 21065
rect 6830 20995 6834 21055
rect 6886 21035 7144 21055
rect 6830 20989 6886 20995
rect 6830 20801 6860 20989
rect 6915 20980 7115 21005
rect 7196 20995 7200 21055
rect 7144 20989 7200 20995
rect 6915 20960 6985 20980
rect 6890 20920 6985 20960
rect 7045 20960 7115 20980
rect 7045 20920 7140 20960
rect 6890 20870 7140 20920
rect 6890 20830 6985 20870
rect 6915 20810 6985 20830
rect 7045 20830 7140 20870
rect 7045 20810 7115 20830
rect 6830 20795 6886 20801
rect 6830 20735 6834 20795
rect 6915 20785 7115 20810
rect 7170 20801 7200 20989
rect 7144 20795 7200 20801
rect 6886 20735 7144 20755
rect 7196 20735 7200 20795
rect 6830 20725 7200 20735
rect 7230 21055 7600 21065
rect 7230 20995 7234 21055
rect 7286 21035 7544 21055
rect 7230 20989 7286 20995
rect 7230 20801 7260 20989
rect 7315 20980 7515 21005
rect 7596 20995 7600 21055
rect 7544 20989 7600 20995
rect 7315 20960 7385 20980
rect 7290 20920 7385 20960
rect 7445 20960 7515 20980
rect 7445 20920 7540 20960
rect 7290 20870 7540 20920
rect 7290 20830 7385 20870
rect 7315 20810 7385 20830
rect 7445 20830 7540 20870
rect 7445 20810 7515 20830
rect 7230 20795 7286 20801
rect 7230 20735 7234 20795
rect 7315 20785 7515 20810
rect 7570 20801 7600 20989
rect 7544 20795 7600 20801
rect 7286 20735 7544 20755
rect 7596 20735 7600 20795
rect 7230 20725 7600 20735
rect 7630 21055 8000 21065
rect 7630 20995 7634 21055
rect 7686 21035 7944 21055
rect 7630 20989 7686 20995
rect 7630 20801 7660 20989
rect 7715 20980 7915 21005
rect 7996 20995 8000 21055
rect 7944 20989 8000 20995
rect 7715 20960 7785 20980
rect 7690 20920 7785 20960
rect 7845 20960 7915 20980
rect 7845 20920 7940 20960
rect 7690 20870 7940 20920
rect 7690 20830 7785 20870
rect 7715 20810 7785 20830
rect 7845 20830 7940 20870
rect 7845 20810 7915 20830
rect 7630 20795 7686 20801
rect 7630 20735 7634 20795
rect 7715 20785 7915 20810
rect 7970 20801 8000 20989
rect 7944 20795 8000 20801
rect 7686 20735 7944 20755
rect 7996 20735 8000 20795
rect 7630 20725 8000 20735
rect 8030 21055 8400 21065
rect 8030 20995 8034 21055
rect 8086 21035 8344 21055
rect 8030 20989 8086 20995
rect 8030 20801 8060 20989
rect 8115 20980 8315 21005
rect 8396 20995 8400 21055
rect 8344 20989 8400 20995
rect 8115 20960 8185 20980
rect 8090 20920 8185 20960
rect 8245 20960 8315 20980
rect 8245 20920 8340 20960
rect 8090 20870 8340 20920
rect 8090 20830 8185 20870
rect 8115 20810 8185 20830
rect 8245 20830 8340 20870
rect 8245 20810 8315 20830
rect 8030 20795 8086 20801
rect 8030 20735 8034 20795
rect 8115 20785 8315 20810
rect 8370 20801 8400 20989
rect 8344 20795 8400 20801
rect 8086 20735 8344 20755
rect 8396 20735 8400 20795
rect 8030 20725 8400 20735
rect 8430 21055 8800 21065
rect 8430 20995 8434 21055
rect 8486 21035 8744 21055
rect 8430 20989 8486 20995
rect 8430 20801 8460 20989
rect 8515 20980 8715 21005
rect 8796 20995 8800 21055
rect 8744 20989 8800 20995
rect 8515 20960 8585 20980
rect 8490 20920 8585 20960
rect 8645 20960 8715 20980
rect 8645 20920 8740 20960
rect 8490 20870 8740 20920
rect 8490 20830 8585 20870
rect 8515 20810 8585 20830
rect 8645 20830 8740 20870
rect 8645 20810 8715 20830
rect 8430 20795 8486 20801
rect 8430 20735 8434 20795
rect 8515 20785 8715 20810
rect 8770 20801 8800 20989
rect 8744 20795 8800 20801
rect 8486 20735 8744 20755
rect 8796 20735 8800 20795
rect 8430 20725 8800 20735
rect 8830 21055 9200 21065
rect 8830 20995 8834 21055
rect 8886 21035 9144 21055
rect 8830 20989 8886 20995
rect 8830 20801 8860 20989
rect 8915 20980 9115 21005
rect 9196 20995 9200 21055
rect 9144 20989 9200 20995
rect 8915 20960 8985 20980
rect 8890 20920 8985 20960
rect 9045 20960 9115 20980
rect 9045 20920 9140 20960
rect 8890 20870 9140 20920
rect 8890 20830 8985 20870
rect 8915 20810 8985 20830
rect 9045 20830 9140 20870
rect 9045 20810 9115 20830
rect 8830 20795 8886 20801
rect 8830 20735 8834 20795
rect 8915 20785 9115 20810
rect 9170 20801 9200 20989
rect 9144 20795 9200 20801
rect 8886 20735 9144 20755
rect 9196 20735 9200 20795
rect 8830 20725 9200 20735
rect 9230 21055 9600 21065
rect 9230 20995 9234 21055
rect 9286 21035 9544 21055
rect 9230 20989 9286 20995
rect 9230 20801 9260 20989
rect 9315 20980 9515 21005
rect 9596 20995 9600 21055
rect 9544 20989 9600 20995
rect 9315 20960 9385 20980
rect 9290 20920 9385 20960
rect 9445 20960 9515 20980
rect 9445 20920 9540 20960
rect 9290 20870 9540 20920
rect 9290 20830 9385 20870
rect 9315 20810 9385 20830
rect 9445 20830 9540 20870
rect 9445 20810 9515 20830
rect 9230 20795 9286 20801
rect 9230 20735 9234 20795
rect 9315 20785 9515 20810
rect 9570 20801 9600 20989
rect 9544 20795 9600 20801
rect 9286 20735 9544 20755
rect 9596 20735 9600 20795
rect 9230 20725 9600 20735
rect 9630 21055 10000 21065
rect 9630 20995 9634 21055
rect 9686 21035 9944 21055
rect 9630 20989 9686 20995
rect 9630 20801 9660 20989
rect 9715 20980 9915 21005
rect 9996 20995 10000 21055
rect 9944 20989 10000 20995
rect 9715 20960 9785 20980
rect 9690 20920 9785 20960
rect 9845 20960 9915 20980
rect 9845 20920 9940 20960
rect 9690 20870 9940 20920
rect 9690 20830 9785 20870
rect 9715 20810 9785 20830
rect 9845 20830 9940 20870
rect 9845 20810 9915 20830
rect 9630 20795 9686 20801
rect 9630 20735 9634 20795
rect 9715 20785 9915 20810
rect 9970 20801 10000 20989
rect 9944 20795 10000 20801
rect 9686 20735 9944 20755
rect 9996 20735 10000 20795
rect 9630 20725 10000 20735
rect 10030 21055 10400 21065
rect 10030 20995 10034 21055
rect 10086 21035 10344 21055
rect 10030 20989 10086 20995
rect 10030 20801 10060 20989
rect 10115 20980 10315 21005
rect 10396 20995 10400 21055
rect 10344 20989 10400 20995
rect 10115 20960 10185 20980
rect 10090 20920 10185 20960
rect 10245 20960 10315 20980
rect 10245 20920 10340 20960
rect 10090 20870 10340 20920
rect 10090 20830 10185 20870
rect 10115 20810 10185 20830
rect 10245 20830 10340 20870
rect 10245 20810 10315 20830
rect 10030 20795 10086 20801
rect 10030 20735 10034 20795
rect 10115 20785 10315 20810
rect 10370 20801 10400 20989
rect 10344 20795 10400 20801
rect 10086 20735 10344 20755
rect 10396 20735 10400 20795
rect 10030 20725 10400 20735
rect 10430 21055 10800 21065
rect 10430 20995 10434 21055
rect 10486 21035 10744 21055
rect 10430 20989 10486 20995
rect 10430 20801 10460 20989
rect 10515 20980 10715 21005
rect 10796 20995 10800 21055
rect 10744 20989 10800 20995
rect 10515 20960 10585 20980
rect 10490 20920 10585 20960
rect 10645 20960 10715 20980
rect 10645 20920 10740 20960
rect 10490 20870 10740 20920
rect 10490 20830 10585 20870
rect 10515 20810 10585 20830
rect 10645 20830 10740 20870
rect 10645 20810 10715 20830
rect 10430 20795 10486 20801
rect 10430 20735 10434 20795
rect 10515 20785 10715 20810
rect 10770 20801 10800 20989
rect 10744 20795 10800 20801
rect 10486 20735 10744 20755
rect 10796 20735 10800 20795
rect 10430 20725 10800 20735
rect 10830 21055 11200 21065
rect 10830 20995 10834 21055
rect 10886 21035 11144 21055
rect 10830 20989 10886 20995
rect 10830 20801 10860 20989
rect 10915 20980 11115 21005
rect 11196 20995 11200 21055
rect 11144 20989 11200 20995
rect 10915 20960 10985 20980
rect 10890 20920 10985 20960
rect 11045 20960 11115 20980
rect 11045 20920 11140 20960
rect 10890 20870 11140 20920
rect 10890 20830 10985 20870
rect 10915 20810 10985 20830
rect 11045 20830 11140 20870
rect 11045 20810 11115 20830
rect 10830 20795 10886 20801
rect 10830 20735 10834 20795
rect 10915 20785 11115 20810
rect 11170 20801 11200 20989
rect 11144 20795 11200 20801
rect 10886 20735 11144 20755
rect 11196 20735 11200 20795
rect 10830 20725 11200 20735
rect 11230 21055 11600 21065
rect 11230 20995 11234 21055
rect 11286 21035 11544 21055
rect 11230 20989 11286 20995
rect 11230 20801 11260 20989
rect 11315 20980 11515 21005
rect 11596 20995 11600 21055
rect 11544 20989 11600 20995
rect 11315 20960 11385 20980
rect 11290 20920 11385 20960
rect 11445 20960 11515 20980
rect 11445 20920 11540 20960
rect 11290 20870 11540 20920
rect 11290 20830 11385 20870
rect 11315 20810 11385 20830
rect 11445 20830 11540 20870
rect 11445 20810 11515 20830
rect 11230 20795 11286 20801
rect 11230 20735 11234 20795
rect 11315 20785 11515 20810
rect 11570 20801 11600 20989
rect 11544 20795 11600 20801
rect 11286 20735 11544 20755
rect 11596 20735 11600 20795
rect 11230 20725 11600 20735
rect 11630 21055 12000 21065
rect 11630 20995 11634 21055
rect 11686 21035 11944 21055
rect 11630 20989 11686 20995
rect 11630 20801 11660 20989
rect 11715 20980 11915 21005
rect 11996 20995 12000 21055
rect 11944 20989 12000 20995
rect 11715 20960 11785 20980
rect 11690 20920 11785 20960
rect 11845 20960 11915 20980
rect 11845 20920 11940 20960
rect 11690 20870 11940 20920
rect 11690 20830 11785 20870
rect 11715 20810 11785 20830
rect 11845 20830 11940 20870
rect 11845 20810 11915 20830
rect 11630 20795 11686 20801
rect 11630 20735 11634 20795
rect 11715 20785 11915 20810
rect 11970 20801 12000 20989
rect 11944 20795 12000 20801
rect 11686 20735 11944 20755
rect 11996 20735 12000 20795
rect 11630 20725 12000 20735
rect 12030 21055 12400 21065
rect 12030 20995 12034 21055
rect 12086 21035 12344 21055
rect 12030 20989 12086 20995
rect 12030 20801 12060 20989
rect 12115 20980 12315 21005
rect 12396 20995 12400 21055
rect 12344 20989 12400 20995
rect 12115 20960 12185 20980
rect 12090 20920 12185 20960
rect 12245 20960 12315 20980
rect 12245 20920 12340 20960
rect 12090 20870 12340 20920
rect 12090 20830 12185 20870
rect 12115 20810 12185 20830
rect 12245 20830 12340 20870
rect 12245 20810 12315 20830
rect 12030 20795 12086 20801
rect 12030 20735 12034 20795
rect 12115 20785 12315 20810
rect 12370 20801 12400 20989
rect 12344 20795 12400 20801
rect 12086 20735 12344 20755
rect 12396 20735 12400 20795
rect 12030 20725 12400 20735
rect 12430 21055 12800 21065
rect 12430 20995 12434 21055
rect 12486 21035 12744 21055
rect 12430 20989 12486 20995
rect 12430 20801 12460 20989
rect 12515 20980 12715 21005
rect 12796 20995 12800 21055
rect 12744 20989 12800 20995
rect 12515 20960 12585 20980
rect 12490 20920 12585 20960
rect 12645 20960 12715 20980
rect 12645 20920 12740 20960
rect 12490 20870 12740 20920
rect 12490 20830 12585 20870
rect 12515 20810 12585 20830
rect 12645 20830 12740 20870
rect 12645 20810 12715 20830
rect 12430 20795 12486 20801
rect 12430 20735 12434 20795
rect 12515 20785 12715 20810
rect 12770 20801 12800 20989
rect 12744 20795 12800 20801
rect 12486 20735 12744 20755
rect 12796 20735 12800 20795
rect 12430 20725 12800 20735
rect 12830 21055 13200 21065
rect 12830 20995 12834 21055
rect 12886 21035 13144 21055
rect 12830 20989 12886 20995
rect 12830 20801 12860 20989
rect 12915 20980 13115 21005
rect 13196 20995 13200 21055
rect 13144 20989 13200 20995
rect 12915 20960 12985 20980
rect 12890 20920 12985 20960
rect 13045 20960 13115 20980
rect 13045 20920 13140 20960
rect 12890 20870 13140 20920
rect 12890 20830 12985 20870
rect 12915 20810 12985 20830
rect 13045 20830 13140 20870
rect 13045 20810 13115 20830
rect 12830 20795 12886 20801
rect 12830 20735 12834 20795
rect 12915 20785 13115 20810
rect 13170 20801 13200 20989
rect 13144 20795 13200 20801
rect 12886 20735 13144 20755
rect 13196 20735 13200 20795
rect 12830 20725 13200 20735
rect -370 20685 0 20695
rect -370 20625 -366 20685
rect -314 20665 -56 20685
rect -370 20619 -314 20625
rect -370 20431 -340 20619
rect -285 20610 -85 20635
rect -4 20625 0 20685
rect -56 20619 0 20625
rect -285 20590 -215 20610
rect -310 20550 -215 20590
rect -155 20590 -85 20610
rect -155 20550 -60 20590
rect -310 20500 -60 20550
rect -310 20460 -215 20500
rect -285 20440 -215 20460
rect -155 20460 -60 20500
rect -155 20440 -85 20460
rect -370 20425 -314 20431
rect -370 20365 -366 20425
rect -285 20415 -85 20440
rect -30 20431 0 20619
rect -56 20425 0 20431
rect -314 20365 -56 20385
rect -4 20365 0 20425
rect -370 20355 0 20365
rect 30 20685 400 20695
rect 30 20625 34 20685
rect 86 20665 344 20685
rect 30 20619 86 20625
rect 30 20431 60 20619
rect 115 20610 315 20635
rect 396 20625 400 20685
rect 344 20619 400 20625
rect 115 20590 185 20610
rect 90 20550 185 20590
rect 245 20590 315 20610
rect 245 20550 340 20590
rect 90 20500 340 20550
rect 90 20460 185 20500
rect 115 20440 185 20460
rect 245 20460 340 20500
rect 245 20440 315 20460
rect 30 20425 86 20431
rect 30 20365 34 20425
rect 115 20415 315 20440
rect 370 20431 400 20619
rect 344 20425 400 20431
rect 86 20365 344 20385
rect 396 20365 400 20425
rect 30 20355 400 20365
rect 430 20685 800 20695
rect 430 20625 434 20685
rect 486 20665 744 20685
rect 430 20619 486 20625
rect 430 20431 460 20619
rect 515 20610 715 20635
rect 796 20625 800 20685
rect 744 20619 800 20625
rect 515 20590 585 20610
rect 490 20550 585 20590
rect 645 20590 715 20610
rect 645 20550 740 20590
rect 490 20500 740 20550
rect 490 20460 585 20500
rect 515 20440 585 20460
rect 645 20460 740 20500
rect 645 20440 715 20460
rect 430 20425 486 20431
rect 430 20365 434 20425
rect 515 20415 715 20440
rect 770 20431 800 20619
rect 744 20425 800 20431
rect 486 20365 744 20385
rect 796 20365 800 20425
rect 430 20355 800 20365
rect 830 20685 1200 20695
rect 830 20625 834 20685
rect 886 20665 1144 20685
rect 830 20619 886 20625
rect 830 20431 860 20619
rect 915 20610 1115 20635
rect 1196 20625 1200 20685
rect 1144 20619 1200 20625
rect 915 20590 985 20610
rect 890 20550 985 20590
rect 1045 20590 1115 20610
rect 1045 20550 1140 20590
rect 890 20500 1140 20550
rect 890 20460 985 20500
rect 915 20440 985 20460
rect 1045 20460 1140 20500
rect 1045 20440 1115 20460
rect 830 20425 886 20431
rect 830 20365 834 20425
rect 915 20415 1115 20440
rect 1170 20431 1200 20619
rect 1144 20425 1200 20431
rect 886 20365 1144 20385
rect 1196 20365 1200 20425
rect 830 20355 1200 20365
rect 1230 20685 1600 20695
rect 1230 20625 1234 20685
rect 1286 20665 1544 20685
rect 1230 20619 1286 20625
rect 1230 20431 1260 20619
rect 1315 20610 1515 20635
rect 1596 20625 1600 20685
rect 1544 20619 1600 20625
rect 1315 20590 1385 20610
rect 1290 20550 1385 20590
rect 1445 20590 1515 20610
rect 1445 20550 1540 20590
rect 1290 20500 1540 20550
rect 1290 20460 1385 20500
rect 1315 20440 1385 20460
rect 1445 20460 1540 20500
rect 1445 20440 1515 20460
rect 1230 20425 1286 20431
rect 1230 20365 1234 20425
rect 1315 20415 1515 20440
rect 1570 20431 1600 20619
rect 1544 20425 1600 20431
rect 1286 20365 1544 20385
rect 1596 20365 1600 20425
rect 1230 20355 1600 20365
rect 1630 20685 2000 20695
rect 1630 20625 1634 20685
rect 1686 20665 1944 20685
rect 1630 20619 1686 20625
rect 1630 20431 1660 20619
rect 1715 20610 1915 20635
rect 1996 20625 2000 20685
rect 1944 20619 2000 20625
rect 1715 20590 1785 20610
rect 1690 20550 1785 20590
rect 1845 20590 1915 20610
rect 1845 20550 1940 20590
rect 1690 20500 1940 20550
rect 1690 20460 1785 20500
rect 1715 20440 1785 20460
rect 1845 20460 1940 20500
rect 1845 20440 1915 20460
rect 1630 20425 1686 20431
rect 1630 20365 1634 20425
rect 1715 20415 1915 20440
rect 1970 20431 2000 20619
rect 1944 20425 2000 20431
rect 1686 20365 1944 20385
rect 1996 20365 2000 20425
rect 1630 20355 2000 20365
rect 2030 20685 2400 20695
rect 2030 20625 2034 20685
rect 2086 20665 2344 20685
rect 2030 20619 2086 20625
rect 2030 20431 2060 20619
rect 2115 20610 2315 20635
rect 2396 20625 2400 20685
rect 2344 20619 2400 20625
rect 2115 20590 2185 20610
rect 2090 20550 2185 20590
rect 2245 20590 2315 20610
rect 2245 20550 2340 20590
rect 2090 20500 2340 20550
rect 2090 20460 2185 20500
rect 2115 20440 2185 20460
rect 2245 20460 2340 20500
rect 2245 20440 2315 20460
rect 2030 20425 2086 20431
rect 2030 20365 2034 20425
rect 2115 20415 2315 20440
rect 2370 20431 2400 20619
rect 2344 20425 2400 20431
rect 2086 20365 2344 20385
rect 2396 20365 2400 20425
rect 2030 20355 2400 20365
rect 2430 20685 2800 20695
rect 2430 20625 2434 20685
rect 2486 20665 2744 20685
rect 2430 20619 2486 20625
rect 2430 20431 2460 20619
rect 2515 20610 2715 20635
rect 2796 20625 2800 20685
rect 2744 20619 2800 20625
rect 2515 20590 2585 20610
rect 2490 20550 2585 20590
rect 2645 20590 2715 20610
rect 2645 20550 2740 20590
rect 2490 20500 2740 20550
rect 2490 20460 2585 20500
rect 2515 20440 2585 20460
rect 2645 20460 2740 20500
rect 2645 20440 2715 20460
rect 2430 20425 2486 20431
rect 2430 20365 2434 20425
rect 2515 20415 2715 20440
rect 2770 20431 2800 20619
rect 2744 20425 2800 20431
rect 2486 20365 2744 20385
rect 2796 20365 2800 20425
rect 2430 20355 2800 20365
rect 2830 20685 3200 20695
rect 2830 20625 2834 20685
rect 2886 20665 3144 20685
rect 2830 20619 2886 20625
rect 2830 20431 2860 20619
rect 2915 20610 3115 20635
rect 3196 20625 3200 20685
rect 3144 20619 3200 20625
rect 2915 20590 2985 20610
rect 2890 20550 2985 20590
rect 3045 20590 3115 20610
rect 3045 20550 3140 20590
rect 2890 20500 3140 20550
rect 2890 20460 2985 20500
rect 2915 20440 2985 20460
rect 3045 20460 3140 20500
rect 3045 20440 3115 20460
rect 2830 20425 2886 20431
rect 2830 20365 2834 20425
rect 2915 20415 3115 20440
rect 3170 20431 3200 20619
rect 3144 20425 3200 20431
rect 2886 20365 3144 20385
rect 3196 20365 3200 20425
rect 2830 20355 3200 20365
rect 3230 20685 3600 20695
rect 3230 20625 3234 20685
rect 3286 20665 3544 20685
rect 3230 20619 3286 20625
rect 3230 20431 3260 20619
rect 3315 20610 3515 20635
rect 3596 20625 3600 20685
rect 3544 20619 3600 20625
rect 3315 20590 3385 20610
rect 3290 20550 3385 20590
rect 3445 20590 3515 20610
rect 3445 20550 3540 20590
rect 3290 20500 3540 20550
rect 3290 20460 3385 20500
rect 3315 20440 3385 20460
rect 3445 20460 3540 20500
rect 3445 20440 3515 20460
rect 3230 20425 3286 20431
rect 3230 20365 3234 20425
rect 3315 20415 3515 20440
rect 3570 20431 3600 20619
rect 3544 20425 3600 20431
rect 3286 20365 3544 20385
rect 3596 20365 3600 20425
rect 3230 20355 3600 20365
rect 3630 20685 4000 20695
rect 3630 20625 3634 20685
rect 3686 20665 3944 20685
rect 3630 20619 3686 20625
rect 3630 20431 3660 20619
rect 3715 20610 3915 20635
rect 3996 20625 4000 20685
rect 3944 20619 4000 20625
rect 3715 20590 3785 20610
rect 3690 20550 3785 20590
rect 3845 20590 3915 20610
rect 3845 20550 3940 20590
rect 3690 20500 3940 20550
rect 3690 20460 3785 20500
rect 3715 20440 3785 20460
rect 3845 20460 3940 20500
rect 3845 20440 3915 20460
rect 3630 20425 3686 20431
rect 3630 20365 3634 20425
rect 3715 20415 3915 20440
rect 3970 20431 4000 20619
rect 3944 20425 4000 20431
rect 3686 20365 3944 20385
rect 3996 20365 4000 20425
rect 3630 20355 4000 20365
rect 4030 20685 4400 20695
rect 4030 20625 4034 20685
rect 4086 20665 4344 20685
rect 4030 20619 4086 20625
rect 4030 20431 4060 20619
rect 4115 20610 4315 20635
rect 4396 20625 4400 20685
rect 4344 20619 4400 20625
rect 4115 20590 4185 20610
rect 4090 20550 4185 20590
rect 4245 20590 4315 20610
rect 4245 20550 4340 20590
rect 4090 20500 4340 20550
rect 4090 20460 4185 20500
rect 4115 20440 4185 20460
rect 4245 20460 4340 20500
rect 4245 20440 4315 20460
rect 4030 20425 4086 20431
rect 4030 20365 4034 20425
rect 4115 20415 4315 20440
rect 4370 20431 4400 20619
rect 4344 20425 4400 20431
rect 4086 20365 4344 20385
rect 4396 20365 4400 20425
rect 4030 20355 4400 20365
rect 4430 20685 4800 20695
rect 4430 20625 4434 20685
rect 4486 20665 4744 20685
rect 4430 20619 4486 20625
rect 4430 20431 4460 20619
rect 4515 20610 4715 20635
rect 4796 20625 4800 20685
rect 4744 20619 4800 20625
rect 4515 20590 4585 20610
rect 4490 20550 4585 20590
rect 4645 20590 4715 20610
rect 4645 20550 4740 20590
rect 4490 20500 4740 20550
rect 4490 20460 4585 20500
rect 4515 20440 4585 20460
rect 4645 20460 4740 20500
rect 4645 20440 4715 20460
rect 4430 20425 4486 20431
rect 4430 20365 4434 20425
rect 4515 20415 4715 20440
rect 4770 20431 4800 20619
rect 4744 20425 4800 20431
rect 4486 20365 4744 20385
rect 4796 20365 4800 20425
rect 4430 20355 4800 20365
rect 4830 20685 5200 20695
rect 4830 20625 4834 20685
rect 4886 20665 5144 20685
rect 4830 20619 4886 20625
rect 4830 20431 4860 20619
rect 4915 20610 5115 20635
rect 5196 20625 5200 20685
rect 5144 20619 5200 20625
rect 4915 20590 4985 20610
rect 4890 20550 4985 20590
rect 5045 20590 5115 20610
rect 5045 20550 5140 20590
rect 4890 20500 5140 20550
rect 4890 20460 4985 20500
rect 4915 20440 4985 20460
rect 5045 20460 5140 20500
rect 5045 20440 5115 20460
rect 4830 20425 4886 20431
rect 4830 20365 4834 20425
rect 4915 20415 5115 20440
rect 5170 20431 5200 20619
rect 5144 20425 5200 20431
rect 4886 20365 5144 20385
rect 5196 20365 5200 20425
rect 4830 20355 5200 20365
rect 5230 20685 5600 20695
rect 5230 20625 5234 20685
rect 5286 20665 5544 20685
rect 5230 20619 5286 20625
rect 5230 20431 5260 20619
rect 5315 20610 5515 20635
rect 5596 20625 5600 20685
rect 5544 20619 5600 20625
rect 5315 20590 5385 20610
rect 5290 20550 5385 20590
rect 5445 20590 5515 20610
rect 5445 20550 5540 20590
rect 5290 20500 5540 20550
rect 5290 20460 5385 20500
rect 5315 20440 5385 20460
rect 5445 20460 5540 20500
rect 5445 20440 5515 20460
rect 5230 20425 5286 20431
rect 5230 20365 5234 20425
rect 5315 20415 5515 20440
rect 5570 20431 5600 20619
rect 5544 20425 5600 20431
rect 5286 20365 5544 20385
rect 5596 20365 5600 20425
rect 5230 20355 5600 20365
rect 5630 20685 6000 20695
rect 5630 20625 5634 20685
rect 5686 20665 5944 20685
rect 5630 20619 5686 20625
rect 5630 20431 5660 20619
rect 5715 20610 5915 20635
rect 5996 20625 6000 20685
rect 5944 20619 6000 20625
rect 5715 20590 5785 20610
rect 5690 20550 5785 20590
rect 5845 20590 5915 20610
rect 5845 20550 5940 20590
rect 5690 20500 5940 20550
rect 5690 20460 5785 20500
rect 5715 20440 5785 20460
rect 5845 20460 5940 20500
rect 5845 20440 5915 20460
rect 5630 20425 5686 20431
rect 5630 20365 5634 20425
rect 5715 20415 5915 20440
rect 5970 20431 6000 20619
rect 5944 20425 6000 20431
rect 5686 20365 5944 20385
rect 5996 20365 6000 20425
rect 5630 20355 6000 20365
rect 6030 20685 6400 20695
rect 6030 20625 6034 20685
rect 6086 20665 6344 20685
rect 6030 20619 6086 20625
rect 6030 20431 6060 20619
rect 6115 20610 6315 20635
rect 6396 20625 6400 20685
rect 6344 20619 6400 20625
rect 6115 20590 6185 20610
rect 6090 20550 6185 20590
rect 6245 20590 6315 20610
rect 6245 20550 6340 20590
rect 6090 20500 6340 20550
rect 6090 20460 6185 20500
rect 6115 20440 6185 20460
rect 6245 20460 6340 20500
rect 6245 20440 6315 20460
rect 6030 20425 6086 20431
rect 6030 20365 6034 20425
rect 6115 20415 6315 20440
rect 6370 20431 6400 20619
rect 6344 20425 6400 20431
rect 6086 20365 6344 20385
rect 6396 20365 6400 20425
rect 6030 20355 6400 20365
rect 6430 20685 6800 20695
rect 6430 20625 6434 20685
rect 6486 20665 6744 20685
rect 6430 20619 6486 20625
rect 6430 20431 6460 20619
rect 6515 20610 6715 20635
rect 6796 20625 6800 20685
rect 6744 20619 6800 20625
rect 6515 20590 6585 20610
rect 6490 20550 6585 20590
rect 6645 20590 6715 20610
rect 6645 20550 6740 20590
rect 6490 20500 6740 20550
rect 6490 20460 6585 20500
rect 6515 20440 6585 20460
rect 6645 20460 6740 20500
rect 6645 20440 6715 20460
rect 6430 20425 6486 20431
rect 6430 20365 6434 20425
rect 6515 20415 6715 20440
rect 6770 20431 6800 20619
rect 6744 20425 6800 20431
rect 6486 20365 6744 20385
rect 6796 20365 6800 20425
rect 6430 20355 6800 20365
rect 6830 20685 7200 20695
rect 6830 20625 6834 20685
rect 6886 20665 7144 20685
rect 6830 20619 6886 20625
rect 6830 20431 6860 20619
rect 6915 20610 7115 20635
rect 7196 20625 7200 20685
rect 7144 20619 7200 20625
rect 6915 20590 6985 20610
rect 6890 20550 6985 20590
rect 7045 20590 7115 20610
rect 7045 20550 7140 20590
rect 6890 20500 7140 20550
rect 6890 20460 6985 20500
rect 6915 20440 6985 20460
rect 7045 20460 7140 20500
rect 7045 20440 7115 20460
rect 6830 20425 6886 20431
rect 6830 20365 6834 20425
rect 6915 20415 7115 20440
rect 7170 20431 7200 20619
rect 7144 20425 7200 20431
rect 6886 20365 7144 20385
rect 7196 20365 7200 20425
rect 6830 20355 7200 20365
rect 7230 20685 7600 20695
rect 7230 20625 7234 20685
rect 7286 20665 7544 20685
rect 7230 20619 7286 20625
rect 7230 20431 7260 20619
rect 7315 20610 7515 20635
rect 7596 20625 7600 20685
rect 7544 20619 7600 20625
rect 7315 20590 7385 20610
rect 7290 20550 7385 20590
rect 7445 20590 7515 20610
rect 7445 20550 7540 20590
rect 7290 20500 7540 20550
rect 7290 20460 7385 20500
rect 7315 20440 7385 20460
rect 7445 20460 7540 20500
rect 7445 20440 7515 20460
rect 7230 20425 7286 20431
rect 7230 20365 7234 20425
rect 7315 20415 7515 20440
rect 7570 20431 7600 20619
rect 7544 20425 7600 20431
rect 7286 20365 7544 20385
rect 7596 20365 7600 20425
rect 7230 20355 7600 20365
rect 7630 20685 8000 20695
rect 7630 20625 7634 20685
rect 7686 20665 7944 20685
rect 7630 20619 7686 20625
rect 7630 20431 7660 20619
rect 7715 20610 7915 20635
rect 7996 20625 8000 20685
rect 7944 20619 8000 20625
rect 7715 20590 7785 20610
rect 7690 20550 7785 20590
rect 7845 20590 7915 20610
rect 7845 20550 7940 20590
rect 7690 20500 7940 20550
rect 7690 20460 7785 20500
rect 7715 20440 7785 20460
rect 7845 20460 7940 20500
rect 7845 20440 7915 20460
rect 7630 20425 7686 20431
rect 7630 20365 7634 20425
rect 7715 20415 7915 20440
rect 7970 20431 8000 20619
rect 7944 20425 8000 20431
rect 7686 20365 7944 20385
rect 7996 20365 8000 20425
rect 7630 20355 8000 20365
rect 8030 20685 8400 20695
rect 8030 20625 8034 20685
rect 8086 20665 8344 20685
rect 8030 20619 8086 20625
rect 8030 20431 8060 20619
rect 8115 20610 8315 20635
rect 8396 20625 8400 20685
rect 8344 20619 8400 20625
rect 8115 20590 8185 20610
rect 8090 20550 8185 20590
rect 8245 20590 8315 20610
rect 8245 20550 8340 20590
rect 8090 20500 8340 20550
rect 8090 20460 8185 20500
rect 8115 20440 8185 20460
rect 8245 20460 8340 20500
rect 8245 20440 8315 20460
rect 8030 20425 8086 20431
rect 8030 20365 8034 20425
rect 8115 20415 8315 20440
rect 8370 20431 8400 20619
rect 8344 20425 8400 20431
rect 8086 20365 8344 20385
rect 8396 20365 8400 20425
rect 8030 20355 8400 20365
rect 8430 20685 8800 20695
rect 8430 20625 8434 20685
rect 8486 20665 8744 20685
rect 8430 20619 8486 20625
rect 8430 20431 8460 20619
rect 8515 20610 8715 20635
rect 8796 20625 8800 20685
rect 8744 20619 8800 20625
rect 8515 20590 8585 20610
rect 8490 20550 8585 20590
rect 8645 20590 8715 20610
rect 8645 20550 8740 20590
rect 8490 20500 8740 20550
rect 8490 20460 8585 20500
rect 8515 20440 8585 20460
rect 8645 20460 8740 20500
rect 8645 20440 8715 20460
rect 8430 20425 8486 20431
rect 8430 20365 8434 20425
rect 8515 20415 8715 20440
rect 8770 20431 8800 20619
rect 8744 20425 8800 20431
rect 8486 20365 8744 20385
rect 8796 20365 8800 20425
rect 8430 20355 8800 20365
rect 8830 20685 9200 20695
rect 8830 20625 8834 20685
rect 8886 20665 9144 20685
rect 8830 20619 8886 20625
rect 8830 20431 8860 20619
rect 8915 20610 9115 20635
rect 9196 20625 9200 20685
rect 9144 20619 9200 20625
rect 8915 20590 8985 20610
rect 8890 20550 8985 20590
rect 9045 20590 9115 20610
rect 9045 20550 9140 20590
rect 8890 20500 9140 20550
rect 8890 20460 8985 20500
rect 8915 20440 8985 20460
rect 9045 20460 9140 20500
rect 9045 20440 9115 20460
rect 8830 20425 8886 20431
rect 8830 20365 8834 20425
rect 8915 20415 9115 20440
rect 9170 20431 9200 20619
rect 9144 20425 9200 20431
rect 8886 20365 9144 20385
rect 9196 20365 9200 20425
rect 8830 20355 9200 20365
rect 9230 20685 9600 20695
rect 9230 20625 9234 20685
rect 9286 20665 9544 20685
rect 9230 20619 9286 20625
rect 9230 20431 9260 20619
rect 9315 20610 9515 20635
rect 9596 20625 9600 20685
rect 9544 20619 9600 20625
rect 9315 20590 9385 20610
rect 9290 20550 9385 20590
rect 9445 20590 9515 20610
rect 9445 20550 9540 20590
rect 9290 20500 9540 20550
rect 9290 20460 9385 20500
rect 9315 20440 9385 20460
rect 9445 20460 9540 20500
rect 9445 20440 9515 20460
rect 9230 20425 9286 20431
rect 9230 20365 9234 20425
rect 9315 20415 9515 20440
rect 9570 20431 9600 20619
rect 9544 20425 9600 20431
rect 9286 20365 9544 20385
rect 9596 20365 9600 20425
rect 9230 20355 9600 20365
rect 9630 20685 10000 20695
rect 9630 20625 9634 20685
rect 9686 20665 9944 20685
rect 9630 20619 9686 20625
rect 9630 20431 9660 20619
rect 9715 20610 9915 20635
rect 9996 20625 10000 20685
rect 9944 20619 10000 20625
rect 9715 20590 9785 20610
rect 9690 20550 9785 20590
rect 9845 20590 9915 20610
rect 9845 20550 9940 20590
rect 9690 20500 9940 20550
rect 9690 20460 9785 20500
rect 9715 20440 9785 20460
rect 9845 20460 9940 20500
rect 9845 20440 9915 20460
rect 9630 20425 9686 20431
rect 9630 20365 9634 20425
rect 9715 20415 9915 20440
rect 9970 20431 10000 20619
rect 9944 20425 10000 20431
rect 9686 20365 9944 20385
rect 9996 20365 10000 20425
rect 9630 20355 10000 20365
rect 10030 20685 10400 20695
rect 10030 20625 10034 20685
rect 10086 20665 10344 20685
rect 10030 20619 10086 20625
rect 10030 20431 10060 20619
rect 10115 20610 10315 20635
rect 10396 20625 10400 20685
rect 10344 20619 10400 20625
rect 10115 20590 10185 20610
rect 10090 20550 10185 20590
rect 10245 20590 10315 20610
rect 10245 20550 10340 20590
rect 10090 20500 10340 20550
rect 10090 20460 10185 20500
rect 10115 20440 10185 20460
rect 10245 20460 10340 20500
rect 10245 20440 10315 20460
rect 10030 20425 10086 20431
rect 10030 20365 10034 20425
rect 10115 20415 10315 20440
rect 10370 20431 10400 20619
rect 10344 20425 10400 20431
rect 10086 20365 10344 20385
rect 10396 20365 10400 20425
rect 10030 20355 10400 20365
rect 10430 20685 10800 20695
rect 10430 20625 10434 20685
rect 10486 20665 10744 20685
rect 10430 20619 10486 20625
rect 10430 20431 10460 20619
rect 10515 20610 10715 20635
rect 10796 20625 10800 20685
rect 10744 20619 10800 20625
rect 10515 20590 10585 20610
rect 10490 20550 10585 20590
rect 10645 20590 10715 20610
rect 10645 20550 10740 20590
rect 10490 20500 10740 20550
rect 10490 20460 10585 20500
rect 10515 20440 10585 20460
rect 10645 20460 10740 20500
rect 10645 20440 10715 20460
rect 10430 20425 10486 20431
rect 10430 20365 10434 20425
rect 10515 20415 10715 20440
rect 10770 20431 10800 20619
rect 10744 20425 10800 20431
rect 10486 20365 10744 20385
rect 10796 20365 10800 20425
rect 10430 20355 10800 20365
rect 10830 20685 11200 20695
rect 10830 20625 10834 20685
rect 10886 20665 11144 20685
rect 10830 20619 10886 20625
rect 10830 20431 10860 20619
rect 10915 20610 11115 20635
rect 11196 20625 11200 20685
rect 11144 20619 11200 20625
rect 10915 20590 10985 20610
rect 10890 20550 10985 20590
rect 11045 20590 11115 20610
rect 11045 20550 11140 20590
rect 10890 20500 11140 20550
rect 10890 20460 10985 20500
rect 10915 20440 10985 20460
rect 11045 20460 11140 20500
rect 11045 20440 11115 20460
rect 10830 20425 10886 20431
rect 10830 20365 10834 20425
rect 10915 20415 11115 20440
rect 11170 20431 11200 20619
rect 11144 20425 11200 20431
rect 10886 20365 11144 20385
rect 11196 20365 11200 20425
rect 10830 20355 11200 20365
rect 11230 20685 11600 20695
rect 11230 20625 11234 20685
rect 11286 20665 11544 20685
rect 11230 20619 11286 20625
rect 11230 20431 11260 20619
rect 11315 20610 11515 20635
rect 11596 20625 11600 20685
rect 11544 20619 11600 20625
rect 11315 20590 11385 20610
rect 11290 20550 11385 20590
rect 11445 20590 11515 20610
rect 11445 20550 11540 20590
rect 11290 20500 11540 20550
rect 11290 20460 11385 20500
rect 11315 20440 11385 20460
rect 11445 20460 11540 20500
rect 11445 20440 11515 20460
rect 11230 20425 11286 20431
rect 11230 20365 11234 20425
rect 11315 20415 11515 20440
rect 11570 20431 11600 20619
rect 11544 20425 11600 20431
rect 11286 20365 11544 20385
rect 11596 20365 11600 20425
rect 11230 20355 11600 20365
rect 11630 20685 12000 20695
rect 11630 20625 11634 20685
rect 11686 20665 11944 20685
rect 11630 20619 11686 20625
rect 11630 20431 11660 20619
rect 11715 20610 11915 20635
rect 11996 20625 12000 20685
rect 11944 20619 12000 20625
rect 11715 20590 11785 20610
rect 11690 20550 11785 20590
rect 11845 20590 11915 20610
rect 11845 20550 11940 20590
rect 11690 20500 11940 20550
rect 11690 20460 11785 20500
rect 11715 20440 11785 20460
rect 11845 20460 11940 20500
rect 11845 20440 11915 20460
rect 11630 20425 11686 20431
rect 11630 20365 11634 20425
rect 11715 20415 11915 20440
rect 11970 20431 12000 20619
rect 11944 20425 12000 20431
rect 11686 20365 11944 20385
rect 11996 20365 12000 20425
rect 11630 20355 12000 20365
rect 12030 20685 12400 20695
rect 12030 20625 12034 20685
rect 12086 20665 12344 20685
rect 12030 20619 12086 20625
rect 12030 20431 12060 20619
rect 12115 20610 12315 20635
rect 12396 20625 12400 20685
rect 12344 20619 12400 20625
rect 12115 20590 12185 20610
rect 12090 20550 12185 20590
rect 12245 20590 12315 20610
rect 12245 20550 12340 20590
rect 12090 20500 12340 20550
rect 12090 20460 12185 20500
rect 12115 20440 12185 20460
rect 12245 20460 12340 20500
rect 12245 20440 12315 20460
rect 12030 20425 12086 20431
rect 12030 20365 12034 20425
rect 12115 20415 12315 20440
rect 12370 20431 12400 20619
rect 12344 20425 12400 20431
rect 12086 20365 12344 20385
rect 12396 20365 12400 20425
rect 12030 20355 12400 20365
rect 12430 20685 12800 20695
rect 12430 20625 12434 20685
rect 12486 20665 12744 20685
rect 12430 20619 12486 20625
rect 12430 20431 12460 20619
rect 12515 20610 12715 20635
rect 12796 20625 12800 20685
rect 12744 20619 12800 20625
rect 12515 20590 12585 20610
rect 12490 20550 12585 20590
rect 12645 20590 12715 20610
rect 12645 20550 12740 20590
rect 12490 20500 12740 20550
rect 12490 20460 12585 20500
rect 12515 20440 12585 20460
rect 12645 20460 12740 20500
rect 12645 20440 12715 20460
rect 12430 20425 12486 20431
rect 12430 20365 12434 20425
rect 12515 20415 12715 20440
rect 12770 20431 12800 20619
rect 12744 20425 12800 20431
rect 12486 20365 12744 20385
rect 12796 20365 12800 20425
rect 12430 20355 12800 20365
rect 12830 20685 13200 20695
rect 12830 20625 12834 20685
rect 12886 20665 13144 20685
rect 12830 20619 12886 20625
rect 12830 20431 12860 20619
rect 12915 20610 13115 20635
rect 13196 20625 13200 20685
rect 13144 20619 13200 20625
rect 12915 20590 12985 20610
rect 12890 20550 12985 20590
rect 13045 20590 13115 20610
rect 13045 20550 13140 20590
rect 12890 20500 13140 20550
rect 12890 20460 12985 20500
rect 12915 20440 12985 20460
rect 13045 20460 13140 20500
rect 13045 20440 13115 20460
rect 12830 20425 12886 20431
rect 12830 20365 12834 20425
rect 12915 20415 13115 20440
rect 13170 20431 13200 20619
rect 13144 20425 13200 20431
rect 12886 20365 13144 20385
rect 13196 20365 13200 20425
rect 12830 20355 13200 20365
rect -370 20315 0 20325
rect -370 20255 -366 20315
rect -314 20295 -56 20315
rect -370 20249 -314 20255
rect -370 20061 -340 20249
rect -285 20240 -85 20265
rect -4 20255 0 20315
rect -56 20249 0 20255
rect -285 20220 -215 20240
rect -310 20180 -215 20220
rect -155 20220 -85 20240
rect -155 20180 -60 20220
rect -310 20130 -60 20180
rect -310 20090 -215 20130
rect -285 20070 -215 20090
rect -155 20090 -60 20130
rect -155 20070 -85 20090
rect -370 20055 -314 20061
rect -370 19995 -366 20055
rect -285 20045 -85 20070
rect -30 20061 0 20249
rect -56 20055 0 20061
rect -314 19995 -56 20015
rect -4 19995 0 20055
rect -370 19985 0 19995
rect 30 20315 400 20325
rect 30 20255 34 20315
rect 86 20295 344 20315
rect 30 20249 86 20255
rect 30 20061 60 20249
rect 115 20240 315 20265
rect 396 20255 400 20315
rect 344 20249 400 20255
rect 115 20220 185 20240
rect 90 20180 185 20220
rect 245 20220 315 20240
rect 245 20180 340 20220
rect 90 20130 340 20180
rect 90 20090 185 20130
rect 115 20070 185 20090
rect 245 20090 340 20130
rect 245 20070 315 20090
rect 30 20055 86 20061
rect 30 19995 34 20055
rect 115 20045 315 20070
rect 370 20061 400 20249
rect 344 20055 400 20061
rect 86 19995 344 20015
rect 396 19995 400 20055
rect 30 19985 400 19995
rect 430 20315 800 20325
rect 430 20255 434 20315
rect 486 20295 744 20315
rect 430 20249 486 20255
rect 430 20061 460 20249
rect 515 20240 715 20265
rect 796 20255 800 20315
rect 744 20249 800 20255
rect 515 20220 585 20240
rect 490 20180 585 20220
rect 645 20220 715 20240
rect 645 20180 740 20220
rect 490 20130 740 20180
rect 490 20090 585 20130
rect 515 20070 585 20090
rect 645 20090 740 20130
rect 645 20070 715 20090
rect 430 20055 486 20061
rect 430 19995 434 20055
rect 515 20045 715 20070
rect 770 20061 800 20249
rect 744 20055 800 20061
rect 486 19995 744 20015
rect 796 19995 800 20055
rect 430 19985 800 19995
rect 830 20315 1200 20325
rect 830 20255 834 20315
rect 886 20295 1144 20315
rect 830 20249 886 20255
rect 830 20061 860 20249
rect 915 20240 1115 20265
rect 1196 20255 1200 20315
rect 1144 20249 1200 20255
rect 915 20220 985 20240
rect 890 20180 985 20220
rect 1045 20220 1115 20240
rect 1045 20180 1140 20220
rect 890 20130 1140 20180
rect 890 20090 985 20130
rect 915 20070 985 20090
rect 1045 20090 1140 20130
rect 1045 20070 1115 20090
rect 830 20055 886 20061
rect 830 19995 834 20055
rect 915 20045 1115 20070
rect 1170 20061 1200 20249
rect 1144 20055 1200 20061
rect 886 19995 1144 20015
rect 1196 19995 1200 20055
rect 830 19985 1200 19995
rect 1230 20315 1600 20325
rect 1230 20255 1234 20315
rect 1286 20295 1544 20315
rect 1230 20249 1286 20255
rect 1230 20061 1260 20249
rect 1315 20240 1515 20265
rect 1596 20255 1600 20315
rect 1544 20249 1600 20255
rect 1315 20220 1385 20240
rect 1290 20180 1385 20220
rect 1445 20220 1515 20240
rect 1445 20180 1540 20220
rect 1290 20130 1540 20180
rect 1290 20090 1385 20130
rect 1315 20070 1385 20090
rect 1445 20090 1540 20130
rect 1445 20070 1515 20090
rect 1230 20055 1286 20061
rect 1230 19995 1234 20055
rect 1315 20045 1515 20070
rect 1570 20061 1600 20249
rect 1544 20055 1600 20061
rect 1286 19995 1544 20015
rect 1596 19995 1600 20055
rect 1230 19985 1600 19995
rect 1630 20315 2000 20325
rect 1630 20255 1634 20315
rect 1686 20295 1944 20315
rect 1630 20249 1686 20255
rect 1630 20061 1660 20249
rect 1715 20240 1915 20265
rect 1996 20255 2000 20315
rect 1944 20249 2000 20255
rect 1715 20220 1785 20240
rect 1690 20180 1785 20220
rect 1845 20220 1915 20240
rect 1845 20180 1940 20220
rect 1690 20130 1940 20180
rect 1690 20090 1785 20130
rect 1715 20070 1785 20090
rect 1845 20090 1940 20130
rect 1845 20070 1915 20090
rect 1630 20055 1686 20061
rect 1630 19995 1634 20055
rect 1715 20045 1915 20070
rect 1970 20061 2000 20249
rect 1944 20055 2000 20061
rect 1686 19995 1944 20015
rect 1996 19995 2000 20055
rect 1630 19985 2000 19995
rect 2030 20315 2400 20325
rect 2030 20255 2034 20315
rect 2086 20295 2344 20315
rect 2030 20249 2086 20255
rect 2030 20061 2060 20249
rect 2115 20240 2315 20265
rect 2396 20255 2400 20315
rect 2344 20249 2400 20255
rect 2115 20220 2185 20240
rect 2090 20180 2185 20220
rect 2245 20220 2315 20240
rect 2245 20180 2340 20220
rect 2090 20130 2340 20180
rect 2090 20090 2185 20130
rect 2115 20070 2185 20090
rect 2245 20090 2340 20130
rect 2245 20070 2315 20090
rect 2030 20055 2086 20061
rect 2030 19995 2034 20055
rect 2115 20045 2315 20070
rect 2370 20061 2400 20249
rect 2344 20055 2400 20061
rect 2086 19995 2344 20015
rect 2396 19995 2400 20055
rect 2030 19985 2400 19995
rect 2430 20315 2800 20325
rect 2430 20255 2434 20315
rect 2486 20295 2744 20315
rect 2430 20249 2486 20255
rect 2430 20061 2460 20249
rect 2515 20240 2715 20265
rect 2796 20255 2800 20315
rect 2744 20249 2800 20255
rect 2515 20220 2585 20240
rect 2490 20180 2585 20220
rect 2645 20220 2715 20240
rect 2645 20180 2740 20220
rect 2490 20130 2740 20180
rect 2490 20090 2585 20130
rect 2515 20070 2585 20090
rect 2645 20090 2740 20130
rect 2645 20070 2715 20090
rect 2430 20055 2486 20061
rect 2430 19995 2434 20055
rect 2515 20045 2715 20070
rect 2770 20061 2800 20249
rect 2744 20055 2800 20061
rect 2486 19995 2744 20015
rect 2796 19995 2800 20055
rect 2430 19985 2800 19995
rect 2830 20315 3200 20325
rect 2830 20255 2834 20315
rect 2886 20295 3144 20315
rect 2830 20249 2886 20255
rect 2830 20061 2860 20249
rect 2915 20240 3115 20265
rect 3196 20255 3200 20315
rect 3144 20249 3200 20255
rect 2915 20220 2985 20240
rect 2890 20180 2985 20220
rect 3045 20220 3115 20240
rect 3045 20180 3140 20220
rect 2890 20130 3140 20180
rect 2890 20090 2985 20130
rect 2915 20070 2985 20090
rect 3045 20090 3140 20130
rect 3045 20070 3115 20090
rect 2830 20055 2886 20061
rect 2830 19995 2834 20055
rect 2915 20045 3115 20070
rect 3170 20061 3200 20249
rect 3144 20055 3200 20061
rect 2886 19995 3144 20015
rect 3196 19995 3200 20055
rect 2830 19985 3200 19995
rect 3230 20315 3600 20325
rect 3230 20255 3234 20315
rect 3286 20295 3544 20315
rect 3230 20249 3286 20255
rect 3230 20061 3260 20249
rect 3315 20240 3515 20265
rect 3596 20255 3600 20315
rect 3544 20249 3600 20255
rect 3315 20220 3385 20240
rect 3290 20180 3385 20220
rect 3445 20220 3515 20240
rect 3445 20180 3540 20220
rect 3290 20130 3540 20180
rect 3290 20090 3385 20130
rect 3315 20070 3385 20090
rect 3445 20090 3540 20130
rect 3445 20070 3515 20090
rect 3230 20055 3286 20061
rect 3230 19995 3234 20055
rect 3315 20045 3515 20070
rect 3570 20061 3600 20249
rect 3544 20055 3600 20061
rect 3286 19995 3544 20015
rect 3596 19995 3600 20055
rect 3230 19985 3600 19995
rect 3630 20315 4000 20325
rect 3630 20255 3634 20315
rect 3686 20295 3944 20315
rect 3630 20249 3686 20255
rect 3630 20061 3660 20249
rect 3715 20240 3915 20265
rect 3996 20255 4000 20315
rect 3944 20249 4000 20255
rect 3715 20220 3785 20240
rect 3690 20180 3785 20220
rect 3845 20220 3915 20240
rect 3845 20180 3940 20220
rect 3690 20130 3940 20180
rect 3690 20090 3785 20130
rect 3715 20070 3785 20090
rect 3845 20090 3940 20130
rect 3845 20070 3915 20090
rect 3630 20055 3686 20061
rect 3630 19995 3634 20055
rect 3715 20045 3915 20070
rect 3970 20061 4000 20249
rect 3944 20055 4000 20061
rect 3686 19995 3944 20015
rect 3996 19995 4000 20055
rect 3630 19985 4000 19995
rect 4030 20315 4400 20325
rect 4030 20255 4034 20315
rect 4086 20295 4344 20315
rect 4030 20249 4086 20255
rect 4030 20061 4060 20249
rect 4115 20240 4315 20265
rect 4396 20255 4400 20315
rect 4344 20249 4400 20255
rect 4115 20220 4185 20240
rect 4090 20180 4185 20220
rect 4245 20220 4315 20240
rect 4245 20180 4340 20220
rect 4090 20130 4340 20180
rect 4090 20090 4185 20130
rect 4115 20070 4185 20090
rect 4245 20090 4340 20130
rect 4245 20070 4315 20090
rect 4030 20055 4086 20061
rect 4030 19995 4034 20055
rect 4115 20045 4315 20070
rect 4370 20061 4400 20249
rect 4344 20055 4400 20061
rect 4086 19995 4344 20015
rect 4396 19995 4400 20055
rect 4030 19985 4400 19995
rect 4430 20315 4800 20325
rect 4430 20255 4434 20315
rect 4486 20295 4744 20315
rect 4430 20249 4486 20255
rect 4430 20061 4460 20249
rect 4515 20240 4715 20265
rect 4796 20255 4800 20315
rect 4744 20249 4800 20255
rect 4515 20220 4585 20240
rect 4490 20180 4585 20220
rect 4645 20220 4715 20240
rect 4645 20180 4740 20220
rect 4490 20130 4740 20180
rect 4490 20090 4585 20130
rect 4515 20070 4585 20090
rect 4645 20090 4740 20130
rect 4645 20070 4715 20090
rect 4430 20055 4486 20061
rect 4430 19995 4434 20055
rect 4515 20045 4715 20070
rect 4770 20061 4800 20249
rect 4744 20055 4800 20061
rect 4486 19995 4744 20015
rect 4796 19995 4800 20055
rect 4430 19985 4800 19995
rect 4830 20315 5200 20325
rect 4830 20255 4834 20315
rect 4886 20295 5144 20315
rect 4830 20249 4886 20255
rect 4830 20061 4860 20249
rect 4915 20240 5115 20265
rect 5196 20255 5200 20315
rect 5144 20249 5200 20255
rect 4915 20220 4985 20240
rect 4890 20180 4985 20220
rect 5045 20220 5115 20240
rect 5045 20180 5140 20220
rect 4890 20130 5140 20180
rect 4890 20090 4985 20130
rect 4915 20070 4985 20090
rect 5045 20090 5140 20130
rect 5045 20070 5115 20090
rect 4830 20055 4886 20061
rect 4830 19995 4834 20055
rect 4915 20045 5115 20070
rect 5170 20061 5200 20249
rect 5144 20055 5200 20061
rect 4886 19995 5144 20015
rect 5196 19995 5200 20055
rect 4830 19985 5200 19995
rect 5230 20315 5600 20325
rect 5230 20255 5234 20315
rect 5286 20295 5544 20315
rect 5230 20249 5286 20255
rect 5230 20061 5260 20249
rect 5315 20240 5515 20265
rect 5596 20255 5600 20315
rect 5544 20249 5600 20255
rect 5315 20220 5385 20240
rect 5290 20180 5385 20220
rect 5445 20220 5515 20240
rect 5445 20180 5540 20220
rect 5290 20130 5540 20180
rect 5290 20090 5385 20130
rect 5315 20070 5385 20090
rect 5445 20090 5540 20130
rect 5445 20070 5515 20090
rect 5230 20055 5286 20061
rect 5230 19995 5234 20055
rect 5315 20045 5515 20070
rect 5570 20061 5600 20249
rect 5544 20055 5600 20061
rect 5286 19995 5544 20015
rect 5596 19995 5600 20055
rect 5230 19985 5600 19995
rect 5630 20315 6000 20325
rect 5630 20255 5634 20315
rect 5686 20295 5944 20315
rect 5630 20249 5686 20255
rect 5630 20061 5660 20249
rect 5715 20240 5915 20265
rect 5996 20255 6000 20315
rect 5944 20249 6000 20255
rect 5715 20220 5785 20240
rect 5690 20180 5785 20220
rect 5845 20220 5915 20240
rect 5845 20180 5940 20220
rect 5690 20130 5940 20180
rect 5690 20090 5785 20130
rect 5715 20070 5785 20090
rect 5845 20090 5940 20130
rect 5845 20070 5915 20090
rect 5630 20055 5686 20061
rect 5630 19995 5634 20055
rect 5715 20045 5915 20070
rect 5970 20061 6000 20249
rect 5944 20055 6000 20061
rect 5686 19995 5944 20015
rect 5996 19995 6000 20055
rect 5630 19985 6000 19995
rect 6030 20315 6400 20325
rect 6030 20255 6034 20315
rect 6086 20295 6344 20315
rect 6030 20249 6086 20255
rect 6030 20061 6060 20249
rect 6115 20240 6315 20265
rect 6396 20255 6400 20315
rect 6344 20249 6400 20255
rect 6115 20220 6185 20240
rect 6090 20180 6185 20220
rect 6245 20220 6315 20240
rect 6245 20180 6340 20220
rect 6090 20130 6340 20180
rect 6090 20090 6185 20130
rect 6115 20070 6185 20090
rect 6245 20090 6340 20130
rect 6245 20070 6315 20090
rect 6030 20055 6086 20061
rect 6030 19995 6034 20055
rect 6115 20045 6315 20070
rect 6370 20061 6400 20249
rect 6344 20055 6400 20061
rect 6086 19995 6344 20015
rect 6396 19995 6400 20055
rect 6030 19985 6400 19995
rect 6430 20315 6800 20325
rect 6430 20255 6434 20315
rect 6486 20295 6744 20315
rect 6430 20249 6486 20255
rect 6430 20061 6460 20249
rect 6515 20240 6715 20265
rect 6796 20255 6800 20315
rect 6744 20249 6800 20255
rect 6515 20220 6585 20240
rect 6490 20180 6585 20220
rect 6645 20220 6715 20240
rect 6645 20180 6740 20220
rect 6490 20130 6740 20180
rect 6490 20090 6585 20130
rect 6515 20070 6585 20090
rect 6645 20090 6740 20130
rect 6645 20070 6715 20090
rect 6430 20055 6486 20061
rect 6430 19995 6434 20055
rect 6515 20045 6715 20070
rect 6770 20061 6800 20249
rect 6744 20055 6800 20061
rect 6486 19995 6744 20015
rect 6796 19995 6800 20055
rect 6430 19985 6800 19995
rect 6830 20315 7200 20325
rect 6830 20255 6834 20315
rect 6886 20295 7144 20315
rect 6830 20249 6886 20255
rect 6830 20061 6860 20249
rect 6915 20240 7115 20265
rect 7196 20255 7200 20315
rect 7144 20249 7200 20255
rect 6915 20220 6985 20240
rect 6890 20180 6985 20220
rect 7045 20220 7115 20240
rect 7045 20180 7140 20220
rect 6890 20130 7140 20180
rect 6890 20090 6985 20130
rect 6915 20070 6985 20090
rect 7045 20090 7140 20130
rect 7045 20070 7115 20090
rect 6830 20055 6886 20061
rect 6830 19995 6834 20055
rect 6915 20045 7115 20070
rect 7170 20061 7200 20249
rect 7144 20055 7200 20061
rect 6886 19995 7144 20015
rect 7196 19995 7200 20055
rect 6830 19985 7200 19995
rect 7230 20315 7600 20325
rect 7230 20255 7234 20315
rect 7286 20295 7544 20315
rect 7230 20249 7286 20255
rect 7230 20061 7260 20249
rect 7315 20240 7515 20265
rect 7596 20255 7600 20315
rect 7544 20249 7600 20255
rect 7315 20220 7385 20240
rect 7290 20180 7385 20220
rect 7445 20220 7515 20240
rect 7445 20180 7540 20220
rect 7290 20130 7540 20180
rect 7290 20090 7385 20130
rect 7315 20070 7385 20090
rect 7445 20090 7540 20130
rect 7445 20070 7515 20090
rect 7230 20055 7286 20061
rect 7230 19995 7234 20055
rect 7315 20045 7515 20070
rect 7570 20061 7600 20249
rect 7544 20055 7600 20061
rect 7286 19995 7544 20015
rect 7596 19995 7600 20055
rect 7230 19985 7600 19995
rect 7630 20315 8000 20325
rect 7630 20255 7634 20315
rect 7686 20295 7944 20315
rect 7630 20249 7686 20255
rect 7630 20061 7660 20249
rect 7715 20240 7915 20265
rect 7996 20255 8000 20315
rect 7944 20249 8000 20255
rect 7715 20220 7785 20240
rect 7690 20180 7785 20220
rect 7845 20220 7915 20240
rect 7845 20180 7940 20220
rect 7690 20130 7940 20180
rect 7690 20090 7785 20130
rect 7715 20070 7785 20090
rect 7845 20090 7940 20130
rect 7845 20070 7915 20090
rect 7630 20055 7686 20061
rect 7630 19995 7634 20055
rect 7715 20045 7915 20070
rect 7970 20061 8000 20249
rect 7944 20055 8000 20061
rect 7686 19995 7944 20015
rect 7996 19995 8000 20055
rect 7630 19985 8000 19995
rect 8030 20315 8400 20325
rect 8030 20255 8034 20315
rect 8086 20295 8344 20315
rect 8030 20249 8086 20255
rect 8030 20061 8060 20249
rect 8115 20240 8315 20265
rect 8396 20255 8400 20315
rect 8344 20249 8400 20255
rect 8115 20220 8185 20240
rect 8090 20180 8185 20220
rect 8245 20220 8315 20240
rect 8245 20180 8340 20220
rect 8090 20130 8340 20180
rect 8090 20090 8185 20130
rect 8115 20070 8185 20090
rect 8245 20090 8340 20130
rect 8245 20070 8315 20090
rect 8030 20055 8086 20061
rect 8030 19995 8034 20055
rect 8115 20045 8315 20070
rect 8370 20061 8400 20249
rect 8344 20055 8400 20061
rect 8086 19995 8344 20015
rect 8396 19995 8400 20055
rect 8030 19985 8400 19995
rect 8430 20315 8800 20325
rect 8430 20255 8434 20315
rect 8486 20295 8744 20315
rect 8430 20249 8486 20255
rect 8430 20061 8460 20249
rect 8515 20240 8715 20265
rect 8796 20255 8800 20315
rect 8744 20249 8800 20255
rect 8515 20220 8585 20240
rect 8490 20180 8585 20220
rect 8645 20220 8715 20240
rect 8645 20180 8740 20220
rect 8490 20130 8740 20180
rect 8490 20090 8585 20130
rect 8515 20070 8585 20090
rect 8645 20090 8740 20130
rect 8645 20070 8715 20090
rect 8430 20055 8486 20061
rect 8430 19995 8434 20055
rect 8515 20045 8715 20070
rect 8770 20061 8800 20249
rect 8744 20055 8800 20061
rect 8486 19995 8744 20015
rect 8796 19995 8800 20055
rect 8430 19985 8800 19995
rect 8830 20315 9200 20325
rect 8830 20255 8834 20315
rect 8886 20295 9144 20315
rect 8830 20249 8886 20255
rect 8830 20061 8860 20249
rect 8915 20240 9115 20265
rect 9196 20255 9200 20315
rect 9144 20249 9200 20255
rect 8915 20220 8985 20240
rect 8890 20180 8985 20220
rect 9045 20220 9115 20240
rect 9045 20180 9140 20220
rect 8890 20130 9140 20180
rect 8890 20090 8985 20130
rect 8915 20070 8985 20090
rect 9045 20090 9140 20130
rect 9045 20070 9115 20090
rect 8830 20055 8886 20061
rect 8830 19995 8834 20055
rect 8915 20045 9115 20070
rect 9170 20061 9200 20249
rect 9144 20055 9200 20061
rect 8886 19995 9144 20015
rect 9196 19995 9200 20055
rect 8830 19985 9200 19995
rect 9230 20315 9600 20325
rect 9230 20255 9234 20315
rect 9286 20295 9544 20315
rect 9230 20249 9286 20255
rect 9230 20061 9260 20249
rect 9315 20240 9515 20265
rect 9596 20255 9600 20315
rect 9544 20249 9600 20255
rect 9315 20220 9385 20240
rect 9290 20180 9385 20220
rect 9445 20220 9515 20240
rect 9445 20180 9540 20220
rect 9290 20130 9540 20180
rect 9290 20090 9385 20130
rect 9315 20070 9385 20090
rect 9445 20090 9540 20130
rect 9445 20070 9515 20090
rect 9230 20055 9286 20061
rect 9230 19995 9234 20055
rect 9315 20045 9515 20070
rect 9570 20061 9600 20249
rect 9544 20055 9600 20061
rect 9286 19995 9544 20015
rect 9596 19995 9600 20055
rect 9230 19985 9600 19995
rect 9630 20315 10000 20325
rect 9630 20255 9634 20315
rect 9686 20295 9944 20315
rect 9630 20249 9686 20255
rect 9630 20061 9660 20249
rect 9715 20240 9915 20265
rect 9996 20255 10000 20315
rect 9944 20249 10000 20255
rect 9715 20220 9785 20240
rect 9690 20180 9785 20220
rect 9845 20220 9915 20240
rect 9845 20180 9940 20220
rect 9690 20130 9940 20180
rect 9690 20090 9785 20130
rect 9715 20070 9785 20090
rect 9845 20090 9940 20130
rect 9845 20070 9915 20090
rect 9630 20055 9686 20061
rect 9630 19995 9634 20055
rect 9715 20045 9915 20070
rect 9970 20061 10000 20249
rect 9944 20055 10000 20061
rect 9686 19995 9944 20015
rect 9996 19995 10000 20055
rect 9630 19985 10000 19995
rect 10030 20315 10400 20325
rect 10030 20255 10034 20315
rect 10086 20295 10344 20315
rect 10030 20249 10086 20255
rect 10030 20061 10060 20249
rect 10115 20240 10315 20265
rect 10396 20255 10400 20315
rect 10344 20249 10400 20255
rect 10115 20220 10185 20240
rect 10090 20180 10185 20220
rect 10245 20220 10315 20240
rect 10245 20180 10340 20220
rect 10090 20130 10340 20180
rect 10090 20090 10185 20130
rect 10115 20070 10185 20090
rect 10245 20090 10340 20130
rect 10245 20070 10315 20090
rect 10030 20055 10086 20061
rect 10030 19995 10034 20055
rect 10115 20045 10315 20070
rect 10370 20061 10400 20249
rect 10344 20055 10400 20061
rect 10086 19995 10344 20015
rect 10396 19995 10400 20055
rect 10030 19985 10400 19995
rect 10430 20315 10800 20325
rect 10430 20255 10434 20315
rect 10486 20295 10744 20315
rect 10430 20249 10486 20255
rect 10430 20061 10460 20249
rect 10515 20240 10715 20265
rect 10796 20255 10800 20315
rect 10744 20249 10800 20255
rect 10515 20220 10585 20240
rect 10490 20180 10585 20220
rect 10645 20220 10715 20240
rect 10645 20180 10740 20220
rect 10490 20130 10740 20180
rect 10490 20090 10585 20130
rect 10515 20070 10585 20090
rect 10645 20090 10740 20130
rect 10645 20070 10715 20090
rect 10430 20055 10486 20061
rect 10430 19995 10434 20055
rect 10515 20045 10715 20070
rect 10770 20061 10800 20249
rect 10744 20055 10800 20061
rect 10486 19995 10744 20015
rect 10796 19995 10800 20055
rect 10430 19985 10800 19995
rect 10830 20315 11200 20325
rect 10830 20255 10834 20315
rect 10886 20295 11144 20315
rect 10830 20249 10886 20255
rect 10830 20061 10860 20249
rect 10915 20240 11115 20265
rect 11196 20255 11200 20315
rect 11144 20249 11200 20255
rect 10915 20220 10985 20240
rect 10890 20180 10985 20220
rect 11045 20220 11115 20240
rect 11045 20180 11140 20220
rect 10890 20130 11140 20180
rect 10890 20090 10985 20130
rect 10915 20070 10985 20090
rect 11045 20090 11140 20130
rect 11045 20070 11115 20090
rect 10830 20055 10886 20061
rect 10830 19995 10834 20055
rect 10915 20045 11115 20070
rect 11170 20061 11200 20249
rect 11144 20055 11200 20061
rect 10886 19995 11144 20015
rect 11196 19995 11200 20055
rect 10830 19985 11200 19995
rect 11230 20315 11600 20325
rect 11230 20255 11234 20315
rect 11286 20295 11544 20315
rect 11230 20249 11286 20255
rect 11230 20061 11260 20249
rect 11315 20240 11515 20265
rect 11596 20255 11600 20315
rect 11544 20249 11600 20255
rect 11315 20220 11385 20240
rect 11290 20180 11385 20220
rect 11445 20220 11515 20240
rect 11445 20180 11540 20220
rect 11290 20130 11540 20180
rect 11290 20090 11385 20130
rect 11315 20070 11385 20090
rect 11445 20090 11540 20130
rect 11445 20070 11515 20090
rect 11230 20055 11286 20061
rect 11230 19995 11234 20055
rect 11315 20045 11515 20070
rect 11570 20061 11600 20249
rect 11544 20055 11600 20061
rect 11286 19995 11544 20015
rect 11596 19995 11600 20055
rect 11230 19985 11600 19995
rect 11630 20315 12000 20325
rect 11630 20255 11634 20315
rect 11686 20295 11944 20315
rect 11630 20249 11686 20255
rect 11630 20061 11660 20249
rect 11715 20240 11915 20265
rect 11996 20255 12000 20315
rect 11944 20249 12000 20255
rect 11715 20220 11785 20240
rect 11690 20180 11785 20220
rect 11845 20220 11915 20240
rect 11845 20180 11940 20220
rect 11690 20130 11940 20180
rect 11690 20090 11785 20130
rect 11715 20070 11785 20090
rect 11845 20090 11940 20130
rect 11845 20070 11915 20090
rect 11630 20055 11686 20061
rect 11630 19995 11634 20055
rect 11715 20045 11915 20070
rect 11970 20061 12000 20249
rect 11944 20055 12000 20061
rect 11686 19995 11944 20015
rect 11996 19995 12000 20055
rect 11630 19985 12000 19995
rect 12030 20315 12400 20325
rect 12030 20255 12034 20315
rect 12086 20295 12344 20315
rect 12030 20249 12086 20255
rect 12030 20061 12060 20249
rect 12115 20240 12315 20265
rect 12396 20255 12400 20315
rect 12344 20249 12400 20255
rect 12115 20220 12185 20240
rect 12090 20180 12185 20220
rect 12245 20220 12315 20240
rect 12245 20180 12340 20220
rect 12090 20130 12340 20180
rect 12090 20090 12185 20130
rect 12115 20070 12185 20090
rect 12245 20090 12340 20130
rect 12245 20070 12315 20090
rect 12030 20055 12086 20061
rect 12030 19995 12034 20055
rect 12115 20045 12315 20070
rect 12370 20061 12400 20249
rect 12344 20055 12400 20061
rect 12086 19995 12344 20015
rect 12396 19995 12400 20055
rect 12030 19985 12400 19995
rect 12430 20315 12800 20325
rect 12430 20255 12434 20315
rect 12486 20295 12744 20315
rect 12430 20249 12486 20255
rect 12430 20061 12460 20249
rect 12515 20240 12715 20265
rect 12796 20255 12800 20315
rect 12744 20249 12800 20255
rect 12515 20220 12585 20240
rect 12490 20180 12585 20220
rect 12645 20220 12715 20240
rect 12645 20180 12740 20220
rect 12490 20130 12740 20180
rect 12490 20090 12585 20130
rect 12515 20070 12585 20090
rect 12645 20090 12740 20130
rect 12645 20070 12715 20090
rect 12430 20055 12486 20061
rect 12430 19995 12434 20055
rect 12515 20045 12715 20070
rect 12770 20061 12800 20249
rect 12744 20055 12800 20061
rect 12486 19995 12744 20015
rect 12796 19995 12800 20055
rect 12430 19985 12800 19995
rect 12830 20315 13200 20325
rect 12830 20255 12834 20315
rect 12886 20295 13144 20315
rect 12830 20249 12886 20255
rect 12830 20061 12860 20249
rect 12915 20240 13115 20265
rect 13196 20255 13200 20315
rect 13144 20249 13200 20255
rect 12915 20220 12985 20240
rect 12890 20180 12985 20220
rect 13045 20220 13115 20240
rect 13045 20180 13140 20220
rect 12890 20130 13140 20180
rect 12890 20090 12985 20130
rect 12915 20070 12985 20090
rect 13045 20090 13140 20130
rect 13045 20070 13115 20090
rect 12830 20055 12886 20061
rect 12830 19995 12834 20055
rect 12915 20045 13115 20070
rect 13170 20061 13200 20249
rect 13144 20055 13200 20061
rect 12886 19995 13144 20015
rect 13196 19995 13200 20055
rect 12830 19985 13200 19995
rect -370 19945 0 19955
rect -370 19885 -366 19945
rect -314 19925 -56 19945
rect -370 19879 -314 19885
rect -370 19691 -340 19879
rect -285 19870 -85 19895
rect -4 19885 0 19945
rect -56 19879 0 19885
rect -285 19850 -215 19870
rect -310 19810 -215 19850
rect -155 19850 -85 19870
rect -155 19810 -60 19850
rect -310 19760 -60 19810
rect -310 19720 -215 19760
rect -285 19700 -215 19720
rect -155 19720 -60 19760
rect -155 19700 -85 19720
rect -370 19685 -314 19691
rect -370 19625 -366 19685
rect -285 19675 -85 19700
rect -30 19691 0 19879
rect -56 19685 0 19691
rect -314 19625 -56 19645
rect -4 19625 0 19685
rect -370 19615 0 19625
rect 30 19945 400 19955
rect 30 19885 34 19945
rect 86 19925 344 19945
rect 30 19879 86 19885
rect 30 19691 60 19879
rect 115 19870 315 19895
rect 396 19885 400 19945
rect 344 19879 400 19885
rect 115 19850 185 19870
rect 90 19810 185 19850
rect 245 19850 315 19870
rect 245 19810 340 19850
rect 90 19760 340 19810
rect 90 19720 185 19760
rect 115 19700 185 19720
rect 245 19720 340 19760
rect 245 19700 315 19720
rect 30 19685 86 19691
rect 30 19625 34 19685
rect 115 19675 315 19700
rect 370 19691 400 19879
rect 344 19685 400 19691
rect 86 19625 344 19645
rect 396 19625 400 19685
rect 30 19615 400 19625
rect 430 19945 800 19955
rect 430 19885 434 19945
rect 486 19925 744 19945
rect 430 19879 486 19885
rect 430 19691 460 19879
rect 515 19870 715 19895
rect 796 19885 800 19945
rect 744 19879 800 19885
rect 515 19850 585 19870
rect 490 19810 585 19850
rect 645 19850 715 19870
rect 645 19810 740 19850
rect 490 19760 740 19810
rect 490 19720 585 19760
rect 515 19700 585 19720
rect 645 19720 740 19760
rect 645 19700 715 19720
rect 430 19685 486 19691
rect 430 19625 434 19685
rect 515 19675 715 19700
rect 770 19691 800 19879
rect 744 19685 800 19691
rect 486 19625 744 19645
rect 796 19625 800 19685
rect 430 19615 800 19625
rect 830 19945 1200 19955
rect 830 19885 834 19945
rect 886 19925 1144 19945
rect 830 19879 886 19885
rect 830 19691 860 19879
rect 915 19870 1115 19895
rect 1196 19885 1200 19945
rect 1144 19879 1200 19885
rect 915 19850 985 19870
rect 890 19810 985 19850
rect 1045 19850 1115 19870
rect 1045 19810 1140 19850
rect 890 19760 1140 19810
rect 890 19720 985 19760
rect 915 19700 985 19720
rect 1045 19720 1140 19760
rect 1045 19700 1115 19720
rect 830 19685 886 19691
rect 830 19625 834 19685
rect 915 19675 1115 19700
rect 1170 19691 1200 19879
rect 1144 19685 1200 19691
rect 886 19625 1144 19645
rect 1196 19625 1200 19685
rect 830 19615 1200 19625
rect 1230 19945 1600 19955
rect 1230 19885 1234 19945
rect 1286 19925 1544 19945
rect 1230 19879 1286 19885
rect 1230 19691 1260 19879
rect 1315 19870 1515 19895
rect 1596 19885 1600 19945
rect 1544 19879 1600 19885
rect 1315 19850 1385 19870
rect 1290 19810 1385 19850
rect 1445 19850 1515 19870
rect 1445 19810 1540 19850
rect 1290 19760 1540 19810
rect 1290 19720 1385 19760
rect 1315 19700 1385 19720
rect 1445 19720 1540 19760
rect 1445 19700 1515 19720
rect 1230 19685 1286 19691
rect 1230 19625 1234 19685
rect 1315 19675 1515 19700
rect 1570 19691 1600 19879
rect 1544 19685 1600 19691
rect 1286 19625 1544 19645
rect 1596 19625 1600 19685
rect 1230 19615 1600 19625
rect 1630 19945 2000 19955
rect 1630 19885 1634 19945
rect 1686 19925 1944 19945
rect 1630 19879 1686 19885
rect 1630 19691 1660 19879
rect 1715 19870 1915 19895
rect 1996 19885 2000 19945
rect 1944 19879 2000 19885
rect 1715 19850 1785 19870
rect 1690 19810 1785 19850
rect 1845 19850 1915 19870
rect 1845 19810 1940 19850
rect 1690 19760 1940 19810
rect 1690 19720 1785 19760
rect 1715 19700 1785 19720
rect 1845 19720 1940 19760
rect 1845 19700 1915 19720
rect 1630 19685 1686 19691
rect 1630 19625 1634 19685
rect 1715 19675 1915 19700
rect 1970 19691 2000 19879
rect 1944 19685 2000 19691
rect 1686 19625 1944 19645
rect 1996 19625 2000 19685
rect 1630 19615 2000 19625
rect 2030 19945 2400 19955
rect 2030 19885 2034 19945
rect 2086 19925 2344 19945
rect 2030 19879 2086 19885
rect 2030 19691 2060 19879
rect 2115 19870 2315 19895
rect 2396 19885 2400 19945
rect 2344 19879 2400 19885
rect 2115 19850 2185 19870
rect 2090 19810 2185 19850
rect 2245 19850 2315 19870
rect 2245 19810 2340 19850
rect 2090 19760 2340 19810
rect 2090 19720 2185 19760
rect 2115 19700 2185 19720
rect 2245 19720 2340 19760
rect 2245 19700 2315 19720
rect 2030 19685 2086 19691
rect 2030 19625 2034 19685
rect 2115 19675 2315 19700
rect 2370 19691 2400 19879
rect 2344 19685 2400 19691
rect 2086 19625 2344 19645
rect 2396 19625 2400 19685
rect 2030 19615 2400 19625
rect 2430 19945 2800 19955
rect 2430 19885 2434 19945
rect 2486 19925 2744 19945
rect 2430 19879 2486 19885
rect 2430 19691 2460 19879
rect 2515 19870 2715 19895
rect 2796 19885 2800 19945
rect 2744 19879 2800 19885
rect 2515 19850 2585 19870
rect 2490 19810 2585 19850
rect 2645 19850 2715 19870
rect 2645 19810 2740 19850
rect 2490 19760 2740 19810
rect 2490 19720 2585 19760
rect 2515 19700 2585 19720
rect 2645 19720 2740 19760
rect 2645 19700 2715 19720
rect 2430 19685 2486 19691
rect 2430 19625 2434 19685
rect 2515 19675 2715 19700
rect 2770 19691 2800 19879
rect 2744 19685 2800 19691
rect 2486 19625 2744 19645
rect 2796 19625 2800 19685
rect 2430 19615 2800 19625
rect 2830 19945 3200 19955
rect 2830 19885 2834 19945
rect 2886 19925 3144 19945
rect 2830 19879 2886 19885
rect 2830 19691 2860 19879
rect 2915 19870 3115 19895
rect 3196 19885 3200 19945
rect 3144 19879 3200 19885
rect 2915 19850 2985 19870
rect 2890 19810 2985 19850
rect 3045 19850 3115 19870
rect 3045 19810 3140 19850
rect 2890 19760 3140 19810
rect 2890 19720 2985 19760
rect 2915 19700 2985 19720
rect 3045 19720 3140 19760
rect 3045 19700 3115 19720
rect 2830 19685 2886 19691
rect 2830 19625 2834 19685
rect 2915 19675 3115 19700
rect 3170 19691 3200 19879
rect 3144 19685 3200 19691
rect 2886 19625 3144 19645
rect 3196 19625 3200 19685
rect 2830 19615 3200 19625
rect 3230 19945 3600 19955
rect 3230 19885 3234 19945
rect 3286 19925 3544 19945
rect 3230 19879 3286 19885
rect 3230 19691 3260 19879
rect 3315 19870 3515 19895
rect 3596 19885 3600 19945
rect 3544 19879 3600 19885
rect 3315 19850 3385 19870
rect 3290 19810 3385 19850
rect 3445 19850 3515 19870
rect 3445 19810 3540 19850
rect 3290 19760 3540 19810
rect 3290 19720 3385 19760
rect 3315 19700 3385 19720
rect 3445 19720 3540 19760
rect 3445 19700 3515 19720
rect 3230 19685 3286 19691
rect 3230 19625 3234 19685
rect 3315 19675 3515 19700
rect 3570 19691 3600 19879
rect 3544 19685 3600 19691
rect 3286 19625 3544 19645
rect 3596 19625 3600 19685
rect 3230 19615 3600 19625
rect 3630 19945 4000 19955
rect 3630 19885 3634 19945
rect 3686 19925 3944 19945
rect 3630 19879 3686 19885
rect 3630 19691 3660 19879
rect 3715 19870 3915 19895
rect 3996 19885 4000 19945
rect 3944 19879 4000 19885
rect 3715 19850 3785 19870
rect 3690 19810 3785 19850
rect 3845 19850 3915 19870
rect 3845 19810 3940 19850
rect 3690 19760 3940 19810
rect 3690 19720 3785 19760
rect 3715 19700 3785 19720
rect 3845 19720 3940 19760
rect 3845 19700 3915 19720
rect 3630 19685 3686 19691
rect 3630 19625 3634 19685
rect 3715 19675 3915 19700
rect 3970 19691 4000 19879
rect 3944 19685 4000 19691
rect 3686 19625 3944 19645
rect 3996 19625 4000 19685
rect 3630 19615 4000 19625
rect 4030 19945 4400 19955
rect 4030 19885 4034 19945
rect 4086 19925 4344 19945
rect 4030 19879 4086 19885
rect 4030 19691 4060 19879
rect 4115 19870 4315 19895
rect 4396 19885 4400 19945
rect 4344 19879 4400 19885
rect 4115 19850 4185 19870
rect 4090 19810 4185 19850
rect 4245 19850 4315 19870
rect 4245 19810 4340 19850
rect 4090 19760 4340 19810
rect 4090 19720 4185 19760
rect 4115 19700 4185 19720
rect 4245 19720 4340 19760
rect 4245 19700 4315 19720
rect 4030 19685 4086 19691
rect 4030 19625 4034 19685
rect 4115 19675 4315 19700
rect 4370 19691 4400 19879
rect 4344 19685 4400 19691
rect 4086 19625 4344 19645
rect 4396 19625 4400 19685
rect 4030 19615 4400 19625
rect 4430 19945 4800 19955
rect 4430 19885 4434 19945
rect 4486 19925 4744 19945
rect 4430 19879 4486 19885
rect 4430 19691 4460 19879
rect 4515 19870 4715 19895
rect 4796 19885 4800 19945
rect 4744 19879 4800 19885
rect 4515 19850 4585 19870
rect 4490 19810 4585 19850
rect 4645 19850 4715 19870
rect 4645 19810 4740 19850
rect 4490 19760 4740 19810
rect 4490 19720 4585 19760
rect 4515 19700 4585 19720
rect 4645 19720 4740 19760
rect 4645 19700 4715 19720
rect 4430 19685 4486 19691
rect 4430 19625 4434 19685
rect 4515 19675 4715 19700
rect 4770 19691 4800 19879
rect 4744 19685 4800 19691
rect 4486 19625 4744 19645
rect 4796 19625 4800 19685
rect 4430 19615 4800 19625
rect 4830 19945 5200 19955
rect 4830 19885 4834 19945
rect 4886 19925 5144 19945
rect 4830 19879 4886 19885
rect 4830 19691 4860 19879
rect 4915 19870 5115 19895
rect 5196 19885 5200 19945
rect 5144 19879 5200 19885
rect 4915 19850 4985 19870
rect 4890 19810 4985 19850
rect 5045 19850 5115 19870
rect 5045 19810 5140 19850
rect 4890 19760 5140 19810
rect 4890 19720 4985 19760
rect 4915 19700 4985 19720
rect 5045 19720 5140 19760
rect 5045 19700 5115 19720
rect 4830 19685 4886 19691
rect 4830 19625 4834 19685
rect 4915 19675 5115 19700
rect 5170 19691 5200 19879
rect 5144 19685 5200 19691
rect 4886 19625 5144 19645
rect 5196 19625 5200 19685
rect 4830 19615 5200 19625
rect 5230 19945 5600 19955
rect 5230 19885 5234 19945
rect 5286 19925 5544 19945
rect 5230 19879 5286 19885
rect 5230 19691 5260 19879
rect 5315 19870 5515 19895
rect 5596 19885 5600 19945
rect 5544 19879 5600 19885
rect 5315 19850 5385 19870
rect 5290 19810 5385 19850
rect 5445 19850 5515 19870
rect 5445 19810 5540 19850
rect 5290 19760 5540 19810
rect 5290 19720 5385 19760
rect 5315 19700 5385 19720
rect 5445 19720 5540 19760
rect 5445 19700 5515 19720
rect 5230 19685 5286 19691
rect 5230 19625 5234 19685
rect 5315 19675 5515 19700
rect 5570 19691 5600 19879
rect 5544 19685 5600 19691
rect 5286 19625 5544 19645
rect 5596 19625 5600 19685
rect 5230 19615 5600 19625
rect 5630 19945 6000 19955
rect 5630 19885 5634 19945
rect 5686 19925 5944 19945
rect 5630 19879 5686 19885
rect 5630 19691 5660 19879
rect 5715 19870 5915 19895
rect 5996 19885 6000 19945
rect 5944 19879 6000 19885
rect 5715 19850 5785 19870
rect 5690 19810 5785 19850
rect 5845 19850 5915 19870
rect 5845 19810 5940 19850
rect 5690 19760 5940 19810
rect 5690 19720 5785 19760
rect 5715 19700 5785 19720
rect 5845 19720 5940 19760
rect 5845 19700 5915 19720
rect 5630 19685 5686 19691
rect 5630 19625 5634 19685
rect 5715 19675 5915 19700
rect 5970 19691 6000 19879
rect 5944 19685 6000 19691
rect 5686 19625 5944 19645
rect 5996 19625 6000 19685
rect 5630 19615 6000 19625
rect 6030 19945 6400 19955
rect 6030 19885 6034 19945
rect 6086 19925 6344 19945
rect 6030 19879 6086 19885
rect 6030 19691 6060 19879
rect 6115 19870 6315 19895
rect 6396 19885 6400 19945
rect 6344 19879 6400 19885
rect 6115 19850 6185 19870
rect 6090 19810 6185 19850
rect 6245 19850 6315 19870
rect 6245 19810 6340 19850
rect 6090 19760 6340 19810
rect 6090 19720 6185 19760
rect 6115 19700 6185 19720
rect 6245 19720 6340 19760
rect 6245 19700 6315 19720
rect 6030 19685 6086 19691
rect 6030 19625 6034 19685
rect 6115 19675 6315 19700
rect 6370 19691 6400 19879
rect 6344 19685 6400 19691
rect 6086 19625 6344 19645
rect 6396 19625 6400 19685
rect 6030 19615 6400 19625
rect 6430 19945 6800 19955
rect 6430 19885 6434 19945
rect 6486 19925 6744 19945
rect 6430 19879 6486 19885
rect 6430 19691 6460 19879
rect 6515 19870 6715 19895
rect 6796 19885 6800 19945
rect 6744 19879 6800 19885
rect 6515 19850 6585 19870
rect 6490 19810 6585 19850
rect 6645 19850 6715 19870
rect 6645 19810 6740 19850
rect 6490 19760 6740 19810
rect 6490 19720 6585 19760
rect 6515 19700 6585 19720
rect 6645 19720 6740 19760
rect 6645 19700 6715 19720
rect 6430 19685 6486 19691
rect 6430 19625 6434 19685
rect 6515 19675 6715 19700
rect 6770 19691 6800 19879
rect 6744 19685 6800 19691
rect 6486 19625 6744 19645
rect 6796 19625 6800 19685
rect 6430 19615 6800 19625
rect 6830 19945 7200 19955
rect 6830 19885 6834 19945
rect 6886 19925 7144 19945
rect 6830 19879 6886 19885
rect 6830 19691 6860 19879
rect 6915 19870 7115 19895
rect 7196 19885 7200 19945
rect 7144 19879 7200 19885
rect 6915 19850 6985 19870
rect 6890 19810 6985 19850
rect 7045 19850 7115 19870
rect 7045 19810 7140 19850
rect 6890 19760 7140 19810
rect 6890 19720 6985 19760
rect 6915 19700 6985 19720
rect 7045 19720 7140 19760
rect 7045 19700 7115 19720
rect 6830 19685 6886 19691
rect 6830 19625 6834 19685
rect 6915 19675 7115 19700
rect 7170 19691 7200 19879
rect 7144 19685 7200 19691
rect 6886 19625 7144 19645
rect 7196 19625 7200 19685
rect 6830 19615 7200 19625
rect 7230 19945 7600 19955
rect 7230 19885 7234 19945
rect 7286 19925 7544 19945
rect 7230 19879 7286 19885
rect 7230 19691 7260 19879
rect 7315 19870 7515 19895
rect 7596 19885 7600 19945
rect 7544 19879 7600 19885
rect 7315 19850 7385 19870
rect 7290 19810 7385 19850
rect 7445 19850 7515 19870
rect 7445 19810 7540 19850
rect 7290 19760 7540 19810
rect 7290 19720 7385 19760
rect 7315 19700 7385 19720
rect 7445 19720 7540 19760
rect 7445 19700 7515 19720
rect 7230 19685 7286 19691
rect 7230 19625 7234 19685
rect 7315 19675 7515 19700
rect 7570 19691 7600 19879
rect 7544 19685 7600 19691
rect 7286 19625 7544 19645
rect 7596 19625 7600 19685
rect 7230 19615 7600 19625
rect 7630 19945 8000 19955
rect 7630 19885 7634 19945
rect 7686 19925 7944 19945
rect 7630 19879 7686 19885
rect 7630 19691 7660 19879
rect 7715 19870 7915 19895
rect 7996 19885 8000 19945
rect 7944 19879 8000 19885
rect 7715 19850 7785 19870
rect 7690 19810 7785 19850
rect 7845 19850 7915 19870
rect 7845 19810 7940 19850
rect 7690 19760 7940 19810
rect 7690 19720 7785 19760
rect 7715 19700 7785 19720
rect 7845 19720 7940 19760
rect 7845 19700 7915 19720
rect 7630 19685 7686 19691
rect 7630 19625 7634 19685
rect 7715 19675 7915 19700
rect 7970 19691 8000 19879
rect 7944 19685 8000 19691
rect 7686 19625 7944 19645
rect 7996 19625 8000 19685
rect 7630 19615 8000 19625
rect 8030 19945 8400 19955
rect 8030 19885 8034 19945
rect 8086 19925 8344 19945
rect 8030 19879 8086 19885
rect 8030 19691 8060 19879
rect 8115 19870 8315 19895
rect 8396 19885 8400 19945
rect 8344 19879 8400 19885
rect 8115 19850 8185 19870
rect 8090 19810 8185 19850
rect 8245 19850 8315 19870
rect 8245 19810 8340 19850
rect 8090 19760 8340 19810
rect 8090 19720 8185 19760
rect 8115 19700 8185 19720
rect 8245 19720 8340 19760
rect 8245 19700 8315 19720
rect 8030 19685 8086 19691
rect 8030 19625 8034 19685
rect 8115 19675 8315 19700
rect 8370 19691 8400 19879
rect 8344 19685 8400 19691
rect 8086 19625 8344 19645
rect 8396 19625 8400 19685
rect 8030 19615 8400 19625
rect 8430 19945 8800 19955
rect 8430 19885 8434 19945
rect 8486 19925 8744 19945
rect 8430 19879 8486 19885
rect 8430 19691 8460 19879
rect 8515 19870 8715 19895
rect 8796 19885 8800 19945
rect 8744 19879 8800 19885
rect 8515 19850 8585 19870
rect 8490 19810 8585 19850
rect 8645 19850 8715 19870
rect 8645 19810 8740 19850
rect 8490 19760 8740 19810
rect 8490 19720 8585 19760
rect 8515 19700 8585 19720
rect 8645 19720 8740 19760
rect 8645 19700 8715 19720
rect 8430 19685 8486 19691
rect 8430 19625 8434 19685
rect 8515 19675 8715 19700
rect 8770 19691 8800 19879
rect 8744 19685 8800 19691
rect 8486 19625 8744 19645
rect 8796 19625 8800 19685
rect 8430 19615 8800 19625
rect 8830 19945 9200 19955
rect 8830 19885 8834 19945
rect 8886 19925 9144 19945
rect 8830 19879 8886 19885
rect 8830 19691 8860 19879
rect 8915 19870 9115 19895
rect 9196 19885 9200 19945
rect 9144 19879 9200 19885
rect 8915 19850 8985 19870
rect 8890 19810 8985 19850
rect 9045 19850 9115 19870
rect 9045 19810 9140 19850
rect 8890 19760 9140 19810
rect 8890 19720 8985 19760
rect 8915 19700 8985 19720
rect 9045 19720 9140 19760
rect 9045 19700 9115 19720
rect 8830 19685 8886 19691
rect 8830 19625 8834 19685
rect 8915 19675 9115 19700
rect 9170 19691 9200 19879
rect 9144 19685 9200 19691
rect 8886 19625 9144 19645
rect 9196 19625 9200 19685
rect 8830 19615 9200 19625
rect 9230 19945 9600 19955
rect 9230 19885 9234 19945
rect 9286 19925 9544 19945
rect 9230 19879 9286 19885
rect 9230 19691 9260 19879
rect 9315 19870 9515 19895
rect 9596 19885 9600 19945
rect 9544 19879 9600 19885
rect 9315 19850 9385 19870
rect 9290 19810 9385 19850
rect 9445 19850 9515 19870
rect 9445 19810 9540 19850
rect 9290 19760 9540 19810
rect 9290 19720 9385 19760
rect 9315 19700 9385 19720
rect 9445 19720 9540 19760
rect 9445 19700 9515 19720
rect 9230 19685 9286 19691
rect 9230 19625 9234 19685
rect 9315 19675 9515 19700
rect 9570 19691 9600 19879
rect 9544 19685 9600 19691
rect 9286 19625 9544 19645
rect 9596 19625 9600 19685
rect 9230 19615 9600 19625
rect 9630 19945 10000 19955
rect 9630 19885 9634 19945
rect 9686 19925 9944 19945
rect 9630 19879 9686 19885
rect 9630 19691 9660 19879
rect 9715 19870 9915 19895
rect 9996 19885 10000 19945
rect 9944 19879 10000 19885
rect 9715 19850 9785 19870
rect 9690 19810 9785 19850
rect 9845 19850 9915 19870
rect 9845 19810 9940 19850
rect 9690 19760 9940 19810
rect 9690 19720 9785 19760
rect 9715 19700 9785 19720
rect 9845 19720 9940 19760
rect 9845 19700 9915 19720
rect 9630 19685 9686 19691
rect 9630 19625 9634 19685
rect 9715 19675 9915 19700
rect 9970 19691 10000 19879
rect 9944 19685 10000 19691
rect 9686 19625 9944 19645
rect 9996 19625 10000 19685
rect 9630 19615 10000 19625
rect 10030 19945 10400 19955
rect 10030 19885 10034 19945
rect 10086 19925 10344 19945
rect 10030 19879 10086 19885
rect 10030 19691 10060 19879
rect 10115 19870 10315 19895
rect 10396 19885 10400 19945
rect 10344 19879 10400 19885
rect 10115 19850 10185 19870
rect 10090 19810 10185 19850
rect 10245 19850 10315 19870
rect 10245 19810 10340 19850
rect 10090 19760 10340 19810
rect 10090 19720 10185 19760
rect 10115 19700 10185 19720
rect 10245 19720 10340 19760
rect 10245 19700 10315 19720
rect 10030 19685 10086 19691
rect 10030 19625 10034 19685
rect 10115 19675 10315 19700
rect 10370 19691 10400 19879
rect 10344 19685 10400 19691
rect 10086 19625 10344 19645
rect 10396 19625 10400 19685
rect 10030 19615 10400 19625
rect 10430 19945 10800 19955
rect 10430 19885 10434 19945
rect 10486 19925 10744 19945
rect 10430 19879 10486 19885
rect 10430 19691 10460 19879
rect 10515 19870 10715 19895
rect 10796 19885 10800 19945
rect 10744 19879 10800 19885
rect 10515 19850 10585 19870
rect 10490 19810 10585 19850
rect 10645 19850 10715 19870
rect 10645 19810 10740 19850
rect 10490 19760 10740 19810
rect 10490 19720 10585 19760
rect 10515 19700 10585 19720
rect 10645 19720 10740 19760
rect 10645 19700 10715 19720
rect 10430 19685 10486 19691
rect 10430 19625 10434 19685
rect 10515 19675 10715 19700
rect 10770 19691 10800 19879
rect 10744 19685 10800 19691
rect 10486 19625 10744 19645
rect 10796 19625 10800 19685
rect 10430 19615 10800 19625
rect 10830 19945 11200 19955
rect 10830 19885 10834 19945
rect 10886 19925 11144 19945
rect 10830 19879 10886 19885
rect 10830 19691 10860 19879
rect 10915 19870 11115 19895
rect 11196 19885 11200 19945
rect 11144 19879 11200 19885
rect 10915 19850 10985 19870
rect 10890 19810 10985 19850
rect 11045 19850 11115 19870
rect 11045 19810 11140 19850
rect 10890 19760 11140 19810
rect 10890 19720 10985 19760
rect 10915 19700 10985 19720
rect 11045 19720 11140 19760
rect 11045 19700 11115 19720
rect 10830 19685 10886 19691
rect 10830 19625 10834 19685
rect 10915 19675 11115 19700
rect 11170 19691 11200 19879
rect 11144 19685 11200 19691
rect 10886 19625 11144 19645
rect 11196 19625 11200 19685
rect 10830 19615 11200 19625
rect 11230 19945 11600 19955
rect 11230 19885 11234 19945
rect 11286 19925 11544 19945
rect 11230 19879 11286 19885
rect 11230 19691 11260 19879
rect 11315 19870 11515 19895
rect 11596 19885 11600 19945
rect 11544 19879 11600 19885
rect 11315 19850 11385 19870
rect 11290 19810 11385 19850
rect 11445 19850 11515 19870
rect 11445 19810 11540 19850
rect 11290 19760 11540 19810
rect 11290 19720 11385 19760
rect 11315 19700 11385 19720
rect 11445 19720 11540 19760
rect 11445 19700 11515 19720
rect 11230 19685 11286 19691
rect 11230 19625 11234 19685
rect 11315 19675 11515 19700
rect 11570 19691 11600 19879
rect 11544 19685 11600 19691
rect 11286 19625 11544 19645
rect 11596 19625 11600 19685
rect 11230 19615 11600 19625
rect 11630 19945 12000 19955
rect 11630 19885 11634 19945
rect 11686 19925 11944 19945
rect 11630 19879 11686 19885
rect 11630 19691 11660 19879
rect 11715 19870 11915 19895
rect 11996 19885 12000 19945
rect 11944 19879 12000 19885
rect 11715 19850 11785 19870
rect 11690 19810 11785 19850
rect 11845 19850 11915 19870
rect 11845 19810 11940 19850
rect 11690 19760 11940 19810
rect 11690 19720 11785 19760
rect 11715 19700 11785 19720
rect 11845 19720 11940 19760
rect 11845 19700 11915 19720
rect 11630 19685 11686 19691
rect 11630 19625 11634 19685
rect 11715 19675 11915 19700
rect 11970 19691 12000 19879
rect 11944 19685 12000 19691
rect 11686 19625 11944 19645
rect 11996 19625 12000 19685
rect 11630 19615 12000 19625
rect 12030 19945 12400 19955
rect 12030 19885 12034 19945
rect 12086 19925 12344 19945
rect 12030 19879 12086 19885
rect 12030 19691 12060 19879
rect 12115 19870 12315 19895
rect 12396 19885 12400 19945
rect 12344 19879 12400 19885
rect 12115 19850 12185 19870
rect 12090 19810 12185 19850
rect 12245 19850 12315 19870
rect 12245 19810 12340 19850
rect 12090 19760 12340 19810
rect 12090 19720 12185 19760
rect 12115 19700 12185 19720
rect 12245 19720 12340 19760
rect 12245 19700 12315 19720
rect 12030 19685 12086 19691
rect 12030 19625 12034 19685
rect 12115 19675 12315 19700
rect 12370 19691 12400 19879
rect 12344 19685 12400 19691
rect 12086 19625 12344 19645
rect 12396 19625 12400 19685
rect 12030 19615 12400 19625
rect 12430 19945 12800 19955
rect 12430 19885 12434 19945
rect 12486 19925 12744 19945
rect 12430 19879 12486 19885
rect 12430 19691 12460 19879
rect 12515 19870 12715 19895
rect 12796 19885 12800 19945
rect 12744 19879 12800 19885
rect 12515 19850 12585 19870
rect 12490 19810 12585 19850
rect 12645 19850 12715 19870
rect 12645 19810 12740 19850
rect 12490 19760 12740 19810
rect 12490 19720 12585 19760
rect 12515 19700 12585 19720
rect 12645 19720 12740 19760
rect 12645 19700 12715 19720
rect 12430 19685 12486 19691
rect 12430 19625 12434 19685
rect 12515 19675 12715 19700
rect 12770 19691 12800 19879
rect 12744 19685 12800 19691
rect 12486 19625 12744 19645
rect 12796 19625 12800 19685
rect 12430 19615 12800 19625
rect 12830 19945 13200 19955
rect 12830 19885 12834 19945
rect 12886 19925 13144 19945
rect 12830 19879 12886 19885
rect 12830 19691 12860 19879
rect 12915 19870 13115 19895
rect 13196 19885 13200 19945
rect 13144 19879 13200 19885
rect 12915 19850 12985 19870
rect 12890 19810 12985 19850
rect 13045 19850 13115 19870
rect 13045 19810 13140 19850
rect 12890 19760 13140 19810
rect 12890 19720 12985 19760
rect 12915 19700 12985 19720
rect 13045 19720 13140 19760
rect 13045 19700 13115 19720
rect 12830 19685 12886 19691
rect 12830 19625 12834 19685
rect 12915 19675 13115 19700
rect 13170 19691 13200 19879
rect 13144 19685 13200 19691
rect 12886 19625 13144 19645
rect 13196 19625 13200 19685
rect 12830 19615 13200 19625
rect -370 19575 0 19585
rect -370 19515 -366 19575
rect -314 19555 -56 19575
rect -370 19509 -314 19515
rect -370 19321 -340 19509
rect -285 19500 -85 19525
rect -4 19515 0 19575
rect -56 19509 0 19515
rect -285 19480 -215 19500
rect -310 19440 -215 19480
rect -155 19480 -85 19500
rect -155 19440 -60 19480
rect -310 19390 -60 19440
rect -310 19350 -215 19390
rect -285 19330 -215 19350
rect -155 19350 -60 19390
rect -155 19330 -85 19350
rect -370 19315 -314 19321
rect -370 19255 -366 19315
rect -285 19305 -85 19330
rect -30 19321 0 19509
rect -56 19315 0 19321
rect -314 19255 -56 19275
rect -4 19255 0 19315
rect -370 19245 0 19255
rect 30 19575 400 19585
rect 30 19515 34 19575
rect 86 19555 344 19575
rect 30 19509 86 19515
rect 30 19321 60 19509
rect 115 19500 315 19525
rect 396 19515 400 19575
rect 344 19509 400 19515
rect 115 19480 185 19500
rect 90 19440 185 19480
rect 245 19480 315 19500
rect 245 19440 340 19480
rect 90 19390 340 19440
rect 90 19350 185 19390
rect 115 19330 185 19350
rect 245 19350 340 19390
rect 245 19330 315 19350
rect 30 19315 86 19321
rect 30 19255 34 19315
rect 115 19305 315 19330
rect 370 19321 400 19509
rect 344 19315 400 19321
rect 86 19255 344 19275
rect 396 19255 400 19315
rect 30 19245 400 19255
rect 430 19575 800 19585
rect 430 19515 434 19575
rect 486 19555 744 19575
rect 430 19509 486 19515
rect 430 19321 460 19509
rect 515 19500 715 19525
rect 796 19515 800 19575
rect 744 19509 800 19515
rect 515 19480 585 19500
rect 490 19440 585 19480
rect 645 19480 715 19500
rect 645 19440 740 19480
rect 490 19390 740 19440
rect 490 19350 585 19390
rect 515 19330 585 19350
rect 645 19350 740 19390
rect 645 19330 715 19350
rect 430 19315 486 19321
rect 430 19255 434 19315
rect 515 19305 715 19330
rect 770 19321 800 19509
rect 744 19315 800 19321
rect 486 19255 744 19275
rect 796 19255 800 19315
rect 430 19245 800 19255
rect 830 19575 1200 19585
rect 830 19515 834 19575
rect 886 19555 1144 19575
rect 830 19509 886 19515
rect 830 19321 860 19509
rect 915 19500 1115 19525
rect 1196 19515 1200 19575
rect 1144 19509 1200 19515
rect 915 19480 985 19500
rect 890 19440 985 19480
rect 1045 19480 1115 19500
rect 1045 19440 1140 19480
rect 890 19390 1140 19440
rect 890 19350 985 19390
rect 915 19330 985 19350
rect 1045 19350 1140 19390
rect 1045 19330 1115 19350
rect 830 19315 886 19321
rect 830 19255 834 19315
rect 915 19305 1115 19330
rect 1170 19321 1200 19509
rect 1144 19315 1200 19321
rect 886 19255 1144 19275
rect 1196 19255 1200 19315
rect 830 19245 1200 19255
rect 1230 19575 1600 19585
rect 1230 19515 1234 19575
rect 1286 19555 1544 19575
rect 1230 19509 1286 19515
rect 1230 19321 1260 19509
rect 1315 19500 1515 19525
rect 1596 19515 1600 19575
rect 1544 19509 1600 19515
rect 1315 19480 1385 19500
rect 1290 19440 1385 19480
rect 1445 19480 1515 19500
rect 1445 19440 1540 19480
rect 1290 19390 1540 19440
rect 1290 19350 1385 19390
rect 1315 19330 1385 19350
rect 1445 19350 1540 19390
rect 1445 19330 1515 19350
rect 1230 19315 1286 19321
rect 1230 19255 1234 19315
rect 1315 19305 1515 19330
rect 1570 19321 1600 19509
rect 1544 19315 1600 19321
rect 1286 19255 1544 19275
rect 1596 19255 1600 19315
rect 1230 19245 1600 19255
rect 1630 19575 2000 19585
rect 1630 19515 1634 19575
rect 1686 19555 1944 19575
rect 1630 19509 1686 19515
rect 1630 19321 1660 19509
rect 1715 19500 1915 19525
rect 1996 19515 2000 19575
rect 1944 19509 2000 19515
rect 1715 19480 1785 19500
rect 1690 19440 1785 19480
rect 1845 19480 1915 19500
rect 1845 19440 1940 19480
rect 1690 19390 1940 19440
rect 1690 19350 1785 19390
rect 1715 19330 1785 19350
rect 1845 19350 1940 19390
rect 1845 19330 1915 19350
rect 1630 19315 1686 19321
rect 1630 19255 1634 19315
rect 1715 19305 1915 19330
rect 1970 19321 2000 19509
rect 1944 19315 2000 19321
rect 1686 19255 1944 19275
rect 1996 19255 2000 19315
rect 1630 19245 2000 19255
rect 2030 19575 2400 19585
rect 2030 19515 2034 19575
rect 2086 19555 2344 19575
rect 2030 19509 2086 19515
rect 2030 19321 2060 19509
rect 2115 19500 2315 19525
rect 2396 19515 2400 19575
rect 2344 19509 2400 19515
rect 2115 19480 2185 19500
rect 2090 19440 2185 19480
rect 2245 19480 2315 19500
rect 2245 19440 2340 19480
rect 2090 19390 2340 19440
rect 2090 19350 2185 19390
rect 2115 19330 2185 19350
rect 2245 19350 2340 19390
rect 2245 19330 2315 19350
rect 2030 19315 2086 19321
rect 2030 19255 2034 19315
rect 2115 19305 2315 19330
rect 2370 19321 2400 19509
rect 2344 19315 2400 19321
rect 2086 19255 2344 19275
rect 2396 19255 2400 19315
rect 2030 19245 2400 19255
rect 2430 19575 2800 19585
rect 2430 19515 2434 19575
rect 2486 19555 2744 19575
rect 2430 19509 2486 19515
rect 2430 19321 2460 19509
rect 2515 19500 2715 19525
rect 2796 19515 2800 19575
rect 2744 19509 2800 19515
rect 2515 19480 2585 19500
rect 2490 19440 2585 19480
rect 2645 19480 2715 19500
rect 2645 19440 2740 19480
rect 2490 19390 2740 19440
rect 2490 19350 2585 19390
rect 2515 19330 2585 19350
rect 2645 19350 2740 19390
rect 2645 19330 2715 19350
rect 2430 19315 2486 19321
rect 2430 19255 2434 19315
rect 2515 19305 2715 19330
rect 2770 19321 2800 19509
rect 2744 19315 2800 19321
rect 2486 19255 2744 19275
rect 2796 19255 2800 19315
rect 2430 19245 2800 19255
rect 2830 19575 3200 19585
rect 2830 19515 2834 19575
rect 2886 19555 3144 19575
rect 2830 19509 2886 19515
rect 2830 19321 2860 19509
rect 2915 19500 3115 19525
rect 3196 19515 3200 19575
rect 3144 19509 3200 19515
rect 2915 19480 2985 19500
rect 2890 19440 2985 19480
rect 3045 19480 3115 19500
rect 3045 19440 3140 19480
rect 2890 19390 3140 19440
rect 2890 19350 2985 19390
rect 2915 19330 2985 19350
rect 3045 19350 3140 19390
rect 3045 19330 3115 19350
rect 2830 19315 2886 19321
rect 2830 19255 2834 19315
rect 2915 19305 3115 19330
rect 3170 19321 3200 19509
rect 3144 19315 3200 19321
rect 2886 19255 3144 19275
rect 3196 19255 3200 19315
rect 2830 19245 3200 19255
rect 3230 19575 3600 19585
rect 3230 19515 3234 19575
rect 3286 19555 3544 19575
rect 3230 19509 3286 19515
rect 3230 19321 3260 19509
rect 3315 19500 3515 19525
rect 3596 19515 3600 19575
rect 3544 19509 3600 19515
rect 3315 19480 3385 19500
rect 3290 19440 3385 19480
rect 3445 19480 3515 19500
rect 3445 19440 3540 19480
rect 3290 19390 3540 19440
rect 3290 19350 3385 19390
rect 3315 19330 3385 19350
rect 3445 19350 3540 19390
rect 3445 19330 3515 19350
rect 3230 19315 3286 19321
rect 3230 19255 3234 19315
rect 3315 19305 3515 19330
rect 3570 19321 3600 19509
rect 3544 19315 3600 19321
rect 3286 19255 3544 19275
rect 3596 19255 3600 19315
rect 3230 19245 3600 19255
rect 3630 19575 4000 19585
rect 3630 19515 3634 19575
rect 3686 19555 3944 19575
rect 3630 19509 3686 19515
rect 3630 19321 3660 19509
rect 3715 19500 3915 19525
rect 3996 19515 4000 19575
rect 3944 19509 4000 19515
rect 3715 19480 3785 19500
rect 3690 19440 3785 19480
rect 3845 19480 3915 19500
rect 3845 19440 3940 19480
rect 3690 19390 3940 19440
rect 3690 19350 3785 19390
rect 3715 19330 3785 19350
rect 3845 19350 3940 19390
rect 3845 19330 3915 19350
rect 3630 19315 3686 19321
rect 3630 19255 3634 19315
rect 3715 19305 3915 19330
rect 3970 19321 4000 19509
rect 3944 19315 4000 19321
rect 3686 19255 3944 19275
rect 3996 19255 4000 19315
rect 3630 19245 4000 19255
rect 4030 19575 4400 19585
rect 4030 19515 4034 19575
rect 4086 19555 4344 19575
rect 4030 19509 4086 19515
rect 4030 19321 4060 19509
rect 4115 19500 4315 19525
rect 4396 19515 4400 19575
rect 4344 19509 4400 19515
rect 4115 19480 4185 19500
rect 4090 19440 4185 19480
rect 4245 19480 4315 19500
rect 4245 19440 4340 19480
rect 4090 19390 4340 19440
rect 4090 19350 4185 19390
rect 4115 19330 4185 19350
rect 4245 19350 4340 19390
rect 4245 19330 4315 19350
rect 4030 19315 4086 19321
rect 4030 19255 4034 19315
rect 4115 19305 4315 19330
rect 4370 19321 4400 19509
rect 4344 19315 4400 19321
rect 4086 19255 4344 19275
rect 4396 19255 4400 19315
rect 4030 19245 4400 19255
rect 4430 19575 4800 19585
rect 4430 19515 4434 19575
rect 4486 19555 4744 19575
rect 4430 19509 4486 19515
rect 4430 19321 4460 19509
rect 4515 19500 4715 19525
rect 4796 19515 4800 19575
rect 4744 19509 4800 19515
rect 4515 19480 4585 19500
rect 4490 19440 4585 19480
rect 4645 19480 4715 19500
rect 4645 19440 4740 19480
rect 4490 19390 4740 19440
rect 4490 19350 4585 19390
rect 4515 19330 4585 19350
rect 4645 19350 4740 19390
rect 4645 19330 4715 19350
rect 4430 19315 4486 19321
rect 4430 19255 4434 19315
rect 4515 19305 4715 19330
rect 4770 19321 4800 19509
rect 4744 19315 4800 19321
rect 4486 19255 4744 19275
rect 4796 19255 4800 19315
rect 4430 19245 4800 19255
rect 4830 19575 5200 19585
rect 4830 19515 4834 19575
rect 4886 19555 5144 19575
rect 4830 19509 4886 19515
rect 4830 19321 4860 19509
rect 4915 19500 5115 19525
rect 5196 19515 5200 19575
rect 5144 19509 5200 19515
rect 4915 19480 4985 19500
rect 4890 19440 4985 19480
rect 5045 19480 5115 19500
rect 5045 19440 5140 19480
rect 4890 19390 5140 19440
rect 4890 19350 4985 19390
rect 4915 19330 4985 19350
rect 5045 19350 5140 19390
rect 5045 19330 5115 19350
rect 4830 19315 4886 19321
rect 4830 19255 4834 19315
rect 4915 19305 5115 19330
rect 5170 19321 5200 19509
rect 5144 19315 5200 19321
rect 4886 19255 5144 19275
rect 5196 19255 5200 19315
rect 4830 19245 5200 19255
rect 5230 19575 5600 19585
rect 5230 19515 5234 19575
rect 5286 19555 5544 19575
rect 5230 19509 5286 19515
rect 5230 19321 5260 19509
rect 5315 19500 5515 19525
rect 5596 19515 5600 19575
rect 5544 19509 5600 19515
rect 5315 19480 5385 19500
rect 5290 19440 5385 19480
rect 5445 19480 5515 19500
rect 5445 19440 5540 19480
rect 5290 19390 5540 19440
rect 5290 19350 5385 19390
rect 5315 19330 5385 19350
rect 5445 19350 5540 19390
rect 5445 19330 5515 19350
rect 5230 19315 5286 19321
rect 5230 19255 5234 19315
rect 5315 19305 5515 19330
rect 5570 19321 5600 19509
rect 5544 19315 5600 19321
rect 5286 19255 5544 19275
rect 5596 19255 5600 19315
rect 5230 19245 5600 19255
rect 5630 19575 6000 19585
rect 5630 19515 5634 19575
rect 5686 19555 5944 19575
rect 5630 19509 5686 19515
rect 5630 19321 5660 19509
rect 5715 19500 5915 19525
rect 5996 19515 6000 19575
rect 5944 19509 6000 19515
rect 5715 19480 5785 19500
rect 5690 19440 5785 19480
rect 5845 19480 5915 19500
rect 5845 19440 5940 19480
rect 5690 19390 5940 19440
rect 5690 19350 5785 19390
rect 5715 19330 5785 19350
rect 5845 19350 5940 19390
rect 5845 19330 5915 19350
rect 5630 19315 5686 19321
rect 5630 19255 5634 19315
rect 5715 19305 5915 19330
rect 5970 19321 6000 19509
rect 5944 19315 6000 19321
rect 5686 19255 5944 19275
rect 5996 19255 6000 19315
rect 5630 19245 6000 19255
rect 6030 19575 6400 19585
rect 6030 19515 6034 19575
rect 6086 19555 6344 19575
rect 6030 19509 6086 19515
rect 6030 19321 6060 19509
rect 6115 19500 6315 19525
rect 6396 19515 6400 19575
rect 6344 19509 6400 19515
rect 6115 19480 6185 19500
rect 6090 19440 6185 19480
rect 6245 19480 6315 19500
rect 6245 19440 6340 19480
rect 6090 19390 6340 19440
rect 6090 19350 6185 19390
rect 6115 19330 6185 19350
rect 6245 19350 6340 19390
rect 6245 19330 6315 19350
rect 6030 19315 6086 19321
rect 6030 19255 6034 19315
rect 6115 19305 6315 19330
rect 6370 19321 6400 19509
rect 6344 19315 6400 19321
rect 6086 19255 6344 19275
rect 6396 19255 6400 19315
rect 6030 19245 6400 19255
rect 6430 19575 6800 19585
rect 6430 19515 6434 19575
rect 6486 19555 6744 19575
rect 6430 19509 6486 19515
rect 6430 19321 6460 19509
rect 6515 19500 6715 19525
rect 6796 19515 6800 19575
rect 6744 19509 6800 19515
rect 6515 19480 6585 19500
rect 6490 19440 6585 19480
rect 6645 19480 6715 19500
rect 6645 19440 6740 19480
rect 6490 19390 6740 19440
rect 6490 19350 6585 19390
rect 6515 19330 6585 19350
rect 6645 19350 6740 19390
rect 6645 19330 6715 19350
rect 6430 19315 6486 19321
rect 6430 19255 6434 19315
rect 6515 19305 6715 19330
rect 6770 19321 6800 19509
rect 6744 19315 6800 19321
rect 6486 19255 6744 19275
rect 6796 19255 6800 19315
rect 6430 19245 6800 19255
rect 6830 19575 7200 19585
rect 6830 19515 6834 19575
rect 6886 19555 7144 19575
rect 6830 19509 6886 19515
rect 6830 19321 6860 19509
rect 6915 19500 7115 19525
rect 7196 19515 7200 19575
rect 7144 19509 7200 19515
rect 6915 19480 6985 19500
rect 6890 19440 6985 19480
rect 7045 19480 7115 19500
rect 7045 19440 7140 19480
rect 6890 19390 7140 19440
rect 6890 19350 6985 19390
rect 6915 19330 6985 19350
rect 7045 19350 7140 19390
rect 7045 19330 7115 19350
rect 6830 19315 6886 19321
rect 6830 19255 6834 19315
rect 6915 19305 7115 19330
rect 7170 19321 7200 19509
rect 7144 19315 7200 19321
rect 6886 19255 7144 19275
rect 7196 19255 7200 19315
rect 6830 19245 7200 19255
rect 7230 19575 7600 19585
rect 7230 19515 7234 19575
rect 7286 19555 7544 19575
rect 7230 19509 7286 19515
rect 7230 19321 7260 19509
rect 7315 19500 7515 19525
rect 7596 19515 7600 19575
rect 7544 19509 7600 19515
rect 7315 19480 7385 19500
rect 7290 19440 7385 19480
rect 7445 19480 7515 19500
rect 7445 19440 7540 19480
rect 7290 19390 7540 19440
rect 7290 19350 7385 19390
rect 7315 19330 7385 19350
rect 7445 19350 7540 19390
rect 7445 19330 7515 19350
rect 7230 19315 7286 19321
rect 7230 19255 7234 19315
rect 7315 19305 7515 19330
rect 7570 19321 7600 19509
rect 7544 19315 7600 19321
rect 7286 19255 7544 19275
rect 7596 19255 7600 19315
rect 7230 19245 7600 19255
rect 7630 19575 8000 19585
rect 7630 19515 7634 19575
rect 7686 19555 7944 19575
rect 7630 19509 7686 19515
rect 7630 19321 7660 19509
rect 7715 19500 7915 19525
rect 7996 19515 8000 19575
rect 7944 19509 8000 19515
rect 7715 19480 7785 19500
rect 7690 19440 7785 19480
rect 7845 19480 7915 19500
rect 7845 19440 7940 19480
rect 7690 19390 7940 19440
rect 7690 19350 7785 19390
rect 7715 19330 7785 19350
rect 7845 19350 7940 19390
rect 7845 19330 7915 19350
rect 7630 19315 7686 19321
rect 7630 19255 7634 19315
rect 7715 19305 7915 19330
rect 7970 19321 8000 19509
rect 7944 19315 8000 19321
rect 7686 19255 7944 19275
rect 7996 19255 8000 19315
rect 7630 19245 8000 19255
rect 8030 19575 8400 19585
rect 8030 19515 8034 19575
rect 8086 19555 8344 19575
rect 8030 19509 8086 19515
rect 8030 19321 8060 19509
rect 8115 19500 8315 19525
rect 8396 19515 8400 19575
rect 8344 19509 8400 19515
rect 8115 19480 8185 19500
rect 8090 19440 8185 19480
rect 8245 19480 8315 19500
rect 8245 19440 8340 19480
rect 8090 19390 8340 19440
rect 8090 19350 8185 19390
rect 8115 19330 8185 19350
rect 8245 19350 8340 19390
rect 8245 19330 8315 19350
rect 8030 19315 8086 19321
rect 8030 19255 8034 19315
rect 8115 19305 8315 19330
rect 8370 19321 8400 19509
rect 8344 19315 8400 19321
rect 8086 19255 8344 19275
rect 8396 19255 8400 19315
rect 8030 19245 8400 19255
rect 8430 19575 8800 19585
rect 8430 19515 8434 19575
rect 8486 19555 8744 19575
rect 8430 19509 8486 19515
rect 8430 19321 8460 19509
rect 8515 19500 8715 19525
rect 8796 19515 8800 19575
rect 8744 19509 8800 19515
rect 8515 19480 8585 19500
rect 8490 19440 8585 19480
rect 8645 19480 8715 19500
rect 8645 19440 8740 19480
rect 8490 19390 8740 19440
rect 8490 19350 8585 19390
rect 8515 19330 8585 19350
rect 8645 19350 8740 19390
rect 8645 19330 8715 19350
rect 8430 19315 8486 19321
rect 8430 19255 8434 19315
rect 8515 19305 8715 19330
rect 8770 19321 8800 19509
rect 8744 19315 8800 19321
rect 8486 19255 8744 19275
rect 8796 19255 8800 19315
rect 8430 19245 8800 19255
rect 8830 19575 9200 19585
rect 8830 19515 8834 19575
rect 8886 19555 9144 19575
rect 8830 19509 8886 19515
rect 8830 19321 8860 19509
rect 8915 19500 9115 19525
rect 9196 19515 9200 19575
rect 9144 19509 9200 19515
rect 8915 19480 8985 19500
rect 8890 19440 8985 19480
rect 9045 19480 9115 19500
rect 9045 19440 9140 19480
rect 8890 19390 9140 19440
rect 8890 19350 8985 19390
rect 8915 19330 8985 19350
rect 9045 19350 9140 19390
rect 9045 19330 9115 19350
rect 8830 19315 8886 19321
rect 8830 19255 8834 19315
rect 8915 19305 9115 19330
rect 9170 19321 9200 19509
rect 9144 19315 9200 19321
rect 8886 19255 9144 19275
rect 9196 19255 9200 19315
rect 8830 19245 9200 19255
rect 9230 19575 9600 19585
rect 9230 19515 9234 19575
rect 9286 19555 9544 19575
rect 9230 19509 9286 19515
rect 9230 19321 9260 19509
rect 9315 19500 9515 19525
rect 9596 19515 9600 19575
rect 9544 19509 9600 19515
rect 9315 19480 9385 19500
rect 9290 19440 9385 19480
rect 9445 19480 9515 19500
rect 9445 19440 9540 19480
rect 9290 19390 9540 19440
rect 9290 19350 9385 19390
rect 9315 19330 9385 19350
rect 9445 19350 9540 19390
rect 9445 19330 9515 19350
rect 9230 19315 9286 19321
rect 9230 19255 9234 19315
rect 9315 19305 9515 19330
rect 9570 19321 9600 19509
rect 9544 19315 9600 19321
rect 9286 19255 9544 19275
rect 9596 19255 9600 19315
rect 9230 19245 9600 19255
rect 9630 19575 10000 19585
rect 9630 19515 9634 19575
rect 9686 19555 9944 19575
rect 9630 19509 9686 19515
rect 9630 19321 9660 19509
rect 9715 19500 9915 19525
rect 9996 19515 10000 19575
rect 9944 19509 10000 19515
rect 9715 19480 9785 19500
rect 9690 19440 9785 19480
rect 9845 19480 9915 19500
rect 9845 19440 9940 19480
rect 9690 19390 9940 19440
rect 9690 19350 9785 19390
rect 9715 19330 9785 19350
rect 9845 19350 9940 19390
rect 9845 19330 9915 19350
rect 9630 19315 9686 19321
rect 9630 19255 9634 19315
rect 9715 19305 9915 19330
rect 9970 19321 10000 19509
rect 9944 19315 10000 19321
rect 9686 19255 9944 19275
rect 9996 19255 10000 19315
rect 9630 19245 10000 19255
rect 10030 19575 10400 19585
rect 10030 19515 10034 19575
rect 10086 19555 10344 19575
rect 10030 19509 10086 19515
rect 10030 19321 10060 19509
rect 10115 19500 10315 19525
rect 10396 19515 10400 19575
rect 10344 19509 10400 19515
rect 10115 19480 10185 19500
rect 10090 19440 10185 19480
rect 10245 19480 10315 19500
rect 10245 19440 10340 19480
rect 10090 19390 10340 19440
rect 10090 19350 10185 19390
rect 10115 19330 10185 19350
rect 10245 19350 10340 19390
rect 10245 19330 10315 19350
rect 10030 19315 10086 19321
rect 10030 19255 10034 19315
rect 10115 19305 10315 19330
rect 10370 19321 10400 19509
rect 10344 19315 10400 19321
rect 10086 19255 10344 19275
rect 10396 19255 10400 19315
rect 10030 19245 10400 19255
rect 10430 19575 10800 19585
rect 10430 19515 10434 19575
rect 10486 19555 10744 19575
rect 10430 19509 10486 19515
rect 10430 19321 10460 19509
rect 10515 19500 10715 19525
rect 10796 19515 10800 19575
rect 10744 19509 10800 19515
rect 10515 19480 10585 19500
rect 10490 19440 10585 19480
rect 10645 19480 10715 19500
rect 10645 19440 10740 19480
rect 10490 19390 10740 19440
rect 10490 19350 10585 19390
rect 10515 19330 10585 19350
rect 10645 19350 10740 19390
rect 10645 19330 10715 19350
rect 10430 19315 10486 19321
rect 10430 19255 10434 19315
rect 10515 19305 10715 19330
rect 10770 19321 10800 19509
rect 10744 19315 10800 19321
rect 10486 19255 10744 19275
rect 10796 19255 10800 19315
rect 10430 19245 10800 19255
rect 10830 19575 11200 19585
rect 10830 19515 10834 19575
rect 10886 19555 11144 19575
rect 10830 19509 10886 19515
rect 10830 19321 10860 19509
rect 10915 19500 11115 19525
rect 11196 19515 11200 19575
rect 11144 19509 11200 19515
rect 10915 19480 10985 19500
rect 10890 19440 10985 19480
rect 11045 19480 11115 19500
rect 11045 19440 11140 19480
rect 10890 19390 11140 19440
rect 10890 19350 10985 19390
rect 10915 19330 10985 19350
rect 11045 19350 11140 19390
rect 11045 19330 11115 19350
rect 10830 19315 10886 19321
rect 10830 19255 10834 19315
rect 10915 19305 11115 19330
rect 11170 19321 11200 19509
rect 11144 19315 11200 19321
rect 10886 19255 11144 19275
rect 11196 19255 11200 19315
rect 10830 19245 11200 19255
rect 11230 19575 11600 19585
rect 11230 19515 11234 19575
rect 11286 19555 11544 19575
rect 11230 19509 11286 19515
rect 11230 19321 11260 19509
rect 11315 19500 11515 19525
rect 11596 19515 11600 19575
rect 11544 19509 11600 19515
rect 11315 19480 11385 19500
rect 11290 19440 11385 19480
rect 11445 19480 11515 19500
rect 11445 19440 11540 19480
rect 11290 19390 11540 19440
rect 11290 19350 11385 19390
rect 11315 19330 11385 19350
rect 11445 19350 11540 19390
rect 11445 19330 11515 19350
rect 11230 19315 11286 19321
rect 11230 19255 11234 19315
rect 11315 19305 11515 19330
rect 11570 19321 11600 19509
rect 11544 19315 11600 19321
rect 11286 19255 11544 19275
rect 11596 19255 11600 19315
rect 11230 19245 11600 19255
rect 11630 19575 12000 19585
rect 11630 19515 11634 19575
rect 11686 19555 11944 19575
rect 11630 19509 11686 19515
rect 11630 19321 11660 19509
rect 11715 19500 11915 19525
rect 11996 19515 12000 19575
rect 11944 19509 12000 19515
rect 11715 19480 11785 19500
rect 11690 19440 11785 19480
rect 11845 19480 11915 19500
rect 11845 19440 11940 19480
rect 11690 19390 11940 19440
rect 11690 19350 11785 19390
rect 11715 19330 11785 19350
rect 11845 19350 11940 19390
rect 11845 19330 11915 19350
rect 11630 19315 11686 19321
rect 11630 19255 11634 19315
rect 11715 19305 11915 19330
rect 11970 19321 12000 19509
rect 11944 19315 12000 19321
rect 11686 19255 11944 19275
rect 11996 19255 12000 19315
rect 11630 19245 12000 19255
rect 12030 19575 12400 19585
rect 12030 19515 12034 19575
rect 12086 19555 12344 19575
rect 12030 19509 12086 19515
rect 12030 19321 12060 19509
rect 12115 19500 12315 19525
rect 12396 19515 12400 19575
rect 12344 19509 12400 19515
rect 12115 19480 12185 19500
rect 12090 19440 12185 19480
rect 12245 19480 12315 19500
rect 12245 19440 12340 19480
rect 12090 19390 12340 19440
rect 12090 19350 12185 19390
rect 12115 19330 12185 19350
rect 12245 19350 12340 19390
rect 12245 19330 12315 19350
rect 12030 19315 12086 19321
rect 12030 19255 12034 19315
rect 12115 19305 12315 19330
rect 12370 19321 12400 19509
rect 12344 19315 12400 19321
rect 12086 19255 12344 19275
rect 12396 19255 12400 19315
rect 12030 19245 12400 19255
rect 12430 19575 12800 19585
rect 12430 19515 12434 19575
rect 12486 19555 12744 19575
rect 12430 19509 12486 19515
rect 12430 19321 12460 19509
rect 12515 19500 12715 19525
rect 12796 19515 12800 19575
rect 12744 19509 12800 19515
rect 12515 19480 12585 19500
rect 12490 19440 12585 19480
rect 12645 19480 12715 19500
rect 12645 19440 12740 19480
rect 12490 19390 12740 19440
rect 12490 19350 12585 19390
rect 12515 19330 12585 19350
rect 12645 19350 12740 19390
rect 12645 19330 12715 19350
rect 12430 19315 12486 19321
rect 12430 19255 12434 19315
rect 12515 19305 12715 19330
rect 12770 19321 12800 19509
rect 12744 19315 12800 19321
rect 12486 19255 12744 19275
rect 12796 19255 12800 19315
rect 12430 19245 12800 19255
rect 12830 19575 13200 19585
rect 12830 19515 12834 19575
rect 12886 19555 13144 19575
rect 12830 19509 12886 19515
rect 12830 19321 12860 19509
rect 12915 19500 13115 19525
rect 13196 19515 13200 19575
rect 13144 19509 13200 19515
rect 12915 19480 12985 19500
rect 12890 19440 12985 19480
rect 13045 19480 13115 19500
rect 13045 19440 13140 19480
rect 12890 19390 13140 19440
rect 12890 19350 12985 19390
rect 12915 19330 12985 19350
rect 13045 19350 13140 19390
rect 13045 19330 13115 19350
rect 12830 19315 12886 19321
rect 12830 19255 12834 19315
rect 12915 19305 13115 19330
rect 13170 19321 13200 19509
rect 13144 19315 13200 19321
rect 12886 19255 13144 19275
rect 13196 19255 13200 19315
rect 12830 19245 13200 19255
rect -370 19205 0 19215
rect -370 19145 -366 19205
rect -314 19185 -56 19205
rect -370 19139 -314 19145
rect -370 18951 -340 19139
rect -285 19130 -85 19155
rect -4 19145 0 19205
rect -56 19139 0 19145
rect -285 19110 -215 19130
rect -310 19070 -215 19110
rect -155 19110 -85 19130
rect -155 19070 -60 19110
rect -310 19020 -60 19070
rect -310 18980 -215 19020
rect -285 18960 -215 18980
rect -155 18980 -60 19020
rect -155 18960 -85 18980
rect -370 18945 -314 18951
rect -370 18885 -366 18945
rect -285 18935 -85 18960
rect -30 18951 0 19139
rect -56 18945 0 18951
rect -314 18885 -56 18905
rect -4 18885 0 18945
rect -370 18875 0 18885
rect 30 19205 400 19215
rect 30 19145 34 19205
rect 86 19185 344 19205
rect 30 19139 86 19145
rect 30 18951 60 19139
rect 115 19130 315 19155
rect 396 19145 400 19205
rect 344 19139 400 19145
rect 115 19110 185 19130
rect 90 19070 185 19110
rect 245 19110 315 19130
rect 245 19070 340 19110
rect 90 19020 340 19070
rect 90 18980 185 19020
rect 115 18960 185 18980
rect 245 18980 340 19020
rect 245 18960 315 18980
rect 30 18945 86 18951
rect 30 18885 34 18945
rect 115 18935 315 18960
rect 370 18951 400 19139
rect 344 18945 400 18951
rect 86 18885 344 18905
rect 396 18885 400 18945
rect 30 18875 400 18885
rect 430 19205 800 19215
rect 430 19145 434 19205
rect 486 19185 744 19205
rect 430 19139 486 19145
rect 430 18951 460 19139
rect 515 19130 715 19155
rect 796 19145 800 19205
rect 744 19139 800 19145
rect 515 19110 585 19130
rect 490 19070 585 19110
rect 645 19110 715 19130
rect 645 19070 740 19110
rect 490 19020 740 19070
rect 490 18980 585 19020
rect 515 18960 585 18980
rect 645 18980 740 19020
rect 645 18960 715 18980
rect 430 18945 486 18951
rect 430 18885 434 18945
rect 515 18935 715 18960
rect 770 18951 800 19139
rect 744 18945 800 18951
rect 486 18885 744 18905
rect 796 18885 800 18945
rect 430 18875 800 18885
rect 830 19205 1200 19215
rect 830 19145 834 19205
rect 886 19185 1144 19205
rect 830 19139 886 19145
rect 830 18951 860 19139
rect 915 19130 1115 19155
rect 1196 19145 1200 19205
rect 1144 19139 1200 19145
rect 915 19110 985 19130
rect 890 19070 985 19110
rect 1045 19110 1115 19130
rect 1045 19070 1140 19110
rect 890 19020 1140 19070
rect 890 18980 985 19020
rect 915 18960 985 18980
rect 1045 18980 1140 19020
rect 1045 18960 1115 18980
rect 830 18945 886 18951
rect 830 18885 834 18945
rect 915 18935 1115 18960
rect 1170 18951 1200 19139
rect 1144 18945 1200 18951
rect 886 18885 1144 18905
rect 1196 18885 1200 18945
rect 830 18875 1200 18885
rect 1230 19205 1600 19215
rect 1230 19145 1234 19205
rect 1286 19185 1544 19205
rect 1230 19139 1286 19145
rect 1230 18951 1260 19139
rect 1315 19130 1515 19155
rect 1596 19145 1600 19205
rect 1544 19139 1600 19145
rect 1315 19110 1385 19130
rect 1290 19070 1385 19110
rect 1445 19110 1515 19130
rect 1445 19070 1540 19110
rect 1290 19020 1540 19070
rect 1290 18980 1385 19020
rect 1315 18960 1385 18980
rect 1445 18980 1540 19020
rect 1445 18960 1515 18980
rect 1230 18945 1286 18951
rect 1230 18885 1234 18945
rect 1315 18935 1515 18960
rect 1570 18951 1600 19139
rect 1544 18945 1600 18951
rect 1286 18885 1544 18905
rect 1596 18885 1600 18945
rect 1230 18875 1600 18885
rect 1630 19205 2000 19215
rect 1630 19145 1634 19205
rect 1686 19185 1944 19205
rect 1630 19139 1686 19145
rect 1630 18951 1660 19139
rect 1715 19130 1915 19155
rect 1996 19145 2000 19205
rect 1944 19139 2000 19145
rect 1715 19110 1785 19130
rect 1690 19070 1785 19110
rect 1845 19110 1915 19130
rect 1845 19070 1940 19110
rect 1690 19020 1940 19070
rect 1690 18980 1785 19020
rect 1715 18960 1785 18980
rect 1845 18980 1940 19020
rect 1845 18960 1915 18980
rect 1630 18945 1686 18951
rect 1630 18885 1634 18945
rect 1715 18935 1915 18960
rect 1970 18951 2000 19139
rect 1944 18945 2000 18951
rect 1686 18885 1944 18905
rect 1996 18885 2000 18945
rect 1630 18875 2000 18885
rect 2030 19205 2400 19215
rect 2030 19145 2034 19205
rect 2086 19185 2344 19205
rect 2030 19139 2086 19145
rect 2030 18951 2060 19139
rect 2115 19130 2315 19155
rect 2396 19145 2400 19205
rect 2344 19139 2400 19145
rect 2115 19110 2185 19130
rect 2090 19070 2185 19110
rect 2245 19110 2315 19130
rect 2245 19070 2340 19110
rect 2090 19020 2340 19070
rect 2090 18980 2185 19020
rect 2115 18960 2185 18980
rect 2245 18980 2340 19020
rect 2245 18960 2315 18980
rect 2030 18945 2086 18951
rect 2030 18885 2034 18945
rect 2115 18935 2315 18960
rect 2370 18951 2400 19139
rect 2344 18945 2400 18951
rect 2086 18885 2344 18905
rect 2396 18885 2400 18945
rect 2030 18875 2400 18885
rect 2430 19205 2800 19215
rect 2430 19145 2434 19205
rect 2486 19185 2744 19205
rect 2430 19139 2486 19145
rect 2430 18951 2460 19139
rect 2515 19130 2715 19155
rect 2796 19145 2800 19205
rect 2744 19139 2800 19145
rect 2515 19110 2585 19130
rect 2490 19070 2585 19110
rect 2645 19110 2715 19130
rect 2645 19070 2740 19110
rect 2490 19020 2740 19070
rect 2490 18980 2585 19020
rect 2515 18960 2585 18980
rect 2645 18980 2740 19020
rect 2645 18960 2715 18980
rect 2430 18945 2486 18951
rect 2430 18885 2434 18945
rect 2515 18935 2715 18960
rect 2770 18951 2800 19139
rect 2744 18945 2800 18951
rect 2486 18885 2744 18905
rect 2796 18885 2800 18945
rect 2430 18875 2800 18885
rect 2830 19205 3200 19215
rect 2830 19145 2834 19205
rect 2886 19185 3144 19205
rect 2830 19139 2886 19145
rect 2830 18951 2860 19139
rect 2915 19130 3115 19155
rect 3196 19145 3200 19205
rect 3144 19139 3200 19145
rect 2915 19110 2985 19130
rect 2890 19070 2985 19110
rect 3045 19110 3115 19130
rect 3045 19070 3140 19110
rect 2890 19020 3140 19070
rect 2890 18980 2985 19020
rect 2915 18960 2985 18980
rect 3045 18980 3140 19020
rect 3045 18960 3115 18980
rect 2830 18945 2886 18951
rect 2830 18885 2834 18945
rect 2915 18935 3115 18960
rect 3170 18951 3200 19139
rect 3144 18945 3200 18951
rect 2886 18885 3144 18905
rect 3196 18885 3200 18945
rect 2830 18875 3200 18885
rect 3230 19205 3600 19215
rect 3230 19145 3234 19205
rect 3286 19185 3544 19205
rect 3230 19139 3286 19145
rect 3230 18951 3260 19139
rect 3315 19130 3515 19155
rect 3596 19145 3600 19205
rect 3544 19139 3600 19145
rect 3315 19110 3385 19130
rect 3290 19070 3385 19110
rect 3445 19110 3515 19130
rect 3445 19070 3540 19110
rect 3290 19020 3540 19070
rect 3290 18980 3385 19020
rect 3315 18960 3385 18980
rect 3445 18980 3540 19020
rect 3445 18960 3515 18980
rect 3230 18945 3286 18951
rect 3230 18885 3234 18945
rect 3315 18935 3515 18960
rect 3570 18951 3600 19139
rect 3544 18945 3600 18951
rect 3286 18885 3544 18905
rect 3596 18885 3600 18945
rect 3230 18875 3600 18885
rect 3630 19205 4000 19215
rect 3630 19145 3634 19205
rect 3686 19185 3944 19205
rect 3630 19139 3686 19145
rect 3630 18951 3660 19139
rect 3715 19130 3915 19155
rect 3996 19145 4000 19205
rect 3944 19139 4000 19145
rect 3715 19110 3785 19130
rect 3690 19070 3785 19110
rect 3845 19110 3915 19130
rect 3845 19070 3940 19110
rect 3690 19020 3940 19070
rect 3690 18980 3785 19020
rect 3715 18960 3785 18980
rect 3845 18980 3940 19020
rect 3845 18960 3915 18980
rect 3630 18945 3686 18951
rect 3630 18885 3634 18945
rect 3715 18935 3915 18960
rect 3970 18951 4000 19139
rect 3944 18945 4000 18951
rect 3686 18885 3944 18905
rect 3996 18885 4000 18945
rect 3630 18875 4000 18885
rect 4030 19205 4400 19215
rect 4030 19145 4034 19205
rect 4086 19185 4344 19205
rect 4030 19139 4086 19145
rect 4030 18951 4060 19139
rect 4115 19130 4315 19155
rect 4396 19145 4400 19205
rect 4344 19139 4400 19145
rect 4115 19110 4185 19130
rect 4090 19070 4185 19110
rect 4245 19110 4315 19130
rect 4245 19070 4340 19110
rect 4090 19020 4340 19070
rect 4090 18980 4185 19020
rect 4115 18960 4185 18980
rect 4245 18980 4340 19020
rect 4245 18960 4315 18980
rect 4030 18945 4086 18951
rect 4030 18885 4034 18945
rect 4115 18935 4315 18960
rect 4370 18951 4400 19139
rect 4344 18945 4400 18951
rect 4086 18885 4344 18905
rect 4396 18885 4400 18945
rect 4030 18875 4400 18885
rect 4430 19205 4800 19215
rect 4430 19145 4434 19205
rect 4486 19185 4744 19205
rect 4430 19139 4486 19145
rect 4430 18951 4460 19139
rect 4515 19130 4715 19155
rect 4796 19145 4800 19205
rect 4744 19139 4800 19145
rect 4515 19110 4585 19130
rect 4490 19070 4585 19110
rect 4645 19110 4715 19130
rect 4645 19070 4740 19110
rect 4490 19020 4740 19070
rect 4490 18980 4585 19020
rect 4515 18960 4585 18980
rect 4645 18980 4740 19020
rect 4645 18960 4715 18980
rect 4430 18945 4486 18951
rect 4430 18885 4434 18945
rect 4515 18935 4715 18960
rect 4770 18951 4800 19139
rect 4744 18945 4800 18951
rect 4486 18885 4744 18905
rect 4796 18885 4800 18945
rect 4430 18875 4800 18885
rect 4830 19205 5200 19215
rect 4830 19145 4834 19205
rect 4886 19185 5144 19205
rect 4830 19139 4886 19145
rect 4830 18951 4860 19139
rect 4915 19130 5115 19155
rect 5196 19145 5200 19205
rect 5144 19139 5200 19145
rect 4915 19110 4985 19130
rect 4890 19070 4985 19110
rect 5045 19110 5115 19130
rect 5045 19070 5140 19110
rect 4890 19020 5140 19070
rect 4890 18980 4985 19020
rect 4915 18960 4985 18980
rect 5045 18980 5140 19020
rect 5045 18960 5115 18980
rect 4830 18945 4886 18951
rect 4830 18885 4834 18945
rect 4915 18935 5115 18960
rect 5170 18951 5200 19139
rect 5144 18945 5200 18951
rect 4886 18885 5144 18905
rect 5196 18885 5200 18945
rect 4830 18875 5200 18885
rect 5230 19205 5600 19215
rect 5230 19145 5234 19205
rect 5286 19185 5544 19205
rect 5230 19139 5286 19145
rect 5230 18951 5260 19139
rect 5315 19130 5515 19155
rect 5596 19145 5600 19205
rect 5544 19139 5600 19145
rect 5315 19110 5385 19130
rect 5290 19070 5385 19110
rect 5445 19110 5515 19130
rect 5445 19070 5540 19110
rect 5290 19020 5540 19070
rect 5290 18980 5385 19020
rect 5315 18960 5385 18980
rect 5445 18980 5540 19020
rect 5445 18960 5515 18980
rect 5230 18945 5286 18951
rect 5230 18885 5234 18945
rect 5315 18935 5515 18960
rect 5570 18951 5600 19139
rect 5544 18945 5600 18951
rect 5286 18885 5544 18905
rect 5596 18885 5600 18945
rect 5230 18875 5600 18885
rect 5630 19205 6000 19215
rect 5630 19145 5634 19205
rect 5686 19185 5944 19205
rect 5630 19139 5686 19145
rect 5630 18951 5660 19139
rect 5715 19130 5915 19155
rect 5996 19145 6000 19205
rect 5944 19139 6000 19145
rect 5715 19110 5785 19130
rect 5690 19070 5785 19110
rect 5845 19110 5915 19130
rect 5845 19070 5940 19110
rect 5690 19020 5940 19070
rect 5690 18980 5785 19020
rect 5715 18960 5785 18980
rect 5845 18980 5940 19020
rect 5845 18960 5915 18980
rect 5630 18945 5686 18951
rect 5630 18885 5634 18945
rect 5715 18935 5915 18960
rect 5970 18951 6000 19139
rect 5944 18945 6000 18951
rect 5686 18885 5944 18905
rect 5996 18885 6000 18945
rect 5630 18875 6000 18885
rect 6030 19205 6400 19215
rect 6030 19145 6034 19205
rect 6086 19185 6344 19205
rect 6030 19139 6086 19145
rect 6030 18951 6060 19139
rect 6115 19130 6315 19155
rect 6396 19145 6400 19205
rect 6344 19139 6400 19145
rect 6115 19110 6185 19130
rect 6090 19070 6185 19110
rect 6245 19110 6315 19130
rect 6245 19070 6340 19110
rect 6090 19020 6340 19070
rect 6090 18980 6185 19020
rect 6115 18960 6185 18980
rect 6245 18980 6340 19020
rect 6245 18960 6315 18980
rect 6030 18945 6086 18951
rect 6030 18885 6034 18945
rect 6115 18935 6315 18960
rect 6370 18951 6400 19139
rect 6344 18945 6400 18951
rect 6086 18885 6344 18905
rect 6396 18885 6400 18945
rect 6030 18875 6400 18885
rect 6430 19205 6800 19215
rect 6430 19145 6434 19205
rect 6486 19185 6744 19205
rect 6430 19139 6486 19145
rect 6430 18951 6460 19139
rect 6515 19130 6715 19155
rect 6796 19145 6800 19205
rect 6744 19139 6800 19145
rect 6515 19110 6585 19130
rect 6490 19070 6585 19110
rect 6645 19110 6715 19130
rect 6645 19070 6740 19110
rect 6490 19020 6740 19070
rect 6490 18980 6585 19020
rect 6515 18960 6585 18980
rect 6645 18980 6740 19020
rect 6645 18960 6715 18980
rect 6430 18945 6486 18951
rect 6430 18885 6434 18945
rect 6515 18935 6715 18960
rect 6770 18951 6800 19139
rect 6744 18945 6800 18951
rect 6486 18885 6744 18905
rect 6796 18885 6800 18945
rect 6430 18875 6800 18885
rect 6830 19205 7200 19215
rect 6830 19145 6834 19205
rect 6886 19185 7144 19205
rect 6830 19139 6886 19145
rect 6830 18951 6860 19139
rect 6915 19130 7115 19155
rect 7196 19145 7200 19205
rect 7144 19139 7200 19145
rect 6915 19110 6985 19130
rect 6890 19070 6985 19110
rect 7045 19110 7115 19130
rect 7045 19070 7140 19110
rect 6890 19020 7140 19070
rect 6890 18980 6985 19020
rect 6915 18960 6985 18980
rect 7045 18980 7140 19020
rect 7045 18960 7115 18980
rect 6830 18945 6886 18951
rect 6830 18885 6834 18945
rect 6915 18935 7115 18960
rect 7170 18951 7200 19139
rect 7144 18945 7200 18951
rect 6886 18885 7144 18905
rect 7196 18885 7200 18945
rect 6830 18875 7200 18885
rect 7230 19205 7600 19215
rect 7230 19145 7234 19205
rect 7286 19185 7544 19205
rect 7230 19139 7286 19145
rect 7230 18951 7260 19139
rect 7315 19130 7515 19155
rect 7596 19145 7600 19205
rect 7544 19139 7600 19145
rect 7315 19110 7385 19130
rect 7290 19070 7385 19110
rect 7445 19110 7515 19130
rect 7445 19070 7540 19110
rect 7290 19020 7540 19070
rect 7290 18980 7385 19020
rect 7315 18960 7385 18980
rect 7445 18980 7540 19020
rect 7445 18960 7515 18980
rect 7230 18945 7286 18951
rect 7230 18885 7234 18945
rect 7315 18935 7515 18960
rect 7570 18951 7600 19139
rect 7544 18945 7600 18951
rect 7286 18885 7544 18905
rect 7596 18885 7600 18945
rect 7230 18875 7600 18885
rect 7630 19205 8000 19215
rect 7630 19145 7634 19205
rect 7686 19185 7944 19205
rect 7630 19139 7686 19145
rect 7630 18951 7660 19139
rect 7715 19130 7915 19155
rect 7996 19145 8000 19205
rect 7944 19139 8000 19145
rect 7715 19110 7785 19130
rect 7690 19070 7785 19110
rect 7845 19110 7915 19130
rect 7845 19070 7940 19110
rect 7690 19020 7940 19070
rect 7690 18980 7785 19020
rect 7715 18960 7785 18980
rect 7845 18980 7940 19020
rect 7845 18960 7915 18980
rect 7630 18945 7686 18951
rect 7630 18885 7634 18945
rect 7715 18935 7915 18960
rect 7970 18951 8000 19139
rect 7944 18945 8000 18951
rect 7686 18885 7944 18905
rect 7996 18885 8000 18945
rect 7630 18875 8000 18885
rect 8030 19205 8400 19215
rect 8030 19145 8034 19205
rect 8086 19185 8344 19205
rect 8030 19139 8086 19145
rect 8030 18951 8060 19139
rect 8115 19130 8315 19155
rect 8396 19145 8400 19205
rect 8344 19139 8400 19145
rect 8115 19110 8185 19130
rect 8090 19070 8185 19110
rect 8245 19110 8315 19130
rect 8245 19070 8340 19110
rect 8090 19020 8340 19070
rect 8090 18980 8185 19020
rect 8115 18960 8185 18980
rect 8245 18980 8340 19020
rect 8245 18960 8315 18980
rect 8030 18945 8086 18951
rect 8030 18885 8034 18945
rect 8115 18935 8315 18960
rect 8370 18951 8400 19139
rect 8344 18945 8400 18951
rect 8086 18885 8344 18905
rect 8396 18885 8400 18945
rect 8030 18875 8400 18885
rect 8430 19205 8800 19215
rect 8430 19145 8434 19205
rect 8486 19185 8744 19205
rect 8430 19139 8486 19145
rect 8430 18951 8460 19139
rect 8515 19130 8715 19155
rect 8796 19145 8800 19205
rect 8744 19139 8800 19145
rect 8515 19110 8585 19130
rect 8490 19070 8585 19110
rect 8645 19110 8715 19130
rect 8645 19070 8740 19110
rect 8490 19020 8740 19070
rect 8490 18980 8585 19020
rect 8515 18960 8585 18980
rect 8645 18980 8740 19020
rect 8645 18960 8715 18980
rect 8430 18945 8486 18951
rect 8430 18885 8434 18945
rect 8515 18935 8715 18960
rect 8770 18951 8800 19139
rect 8744 18945 8800 18951
rect 8486 18885 8744 18905
rect 8796 18885 8800 18945
rect 8430 18875 8800 18885
rect 8830 19205 9200 19215
rect 8830 19145 8834 19205
rect 8886 19185 9144 19205
rect 8830 19139 8886 19145
rect 8830 18951 8860 19139
rect 8915 19130 9115 19155
rect 9196 19145 9200 19205
rect 9144 19139 9200 19145
rect 8915 19110 8985 19130
rect 8890 19070 8985 19110
rect 9045 19110 9115 19130
rect 9045 19070 9140 19110
rect 8890 19020 9140 19070
rect 8890 18980 8985 19020
rect 8915 18960 8985 18980
rect 9045 18980 9140 19020
rect 9045 18960 9115 18980
rect 8830 18945 8886 18951
rect 8830 18885 8834 18945
rect 8915 18935 9115 18960
rect 9170 18951 9200 19139
rect 9144 18945 9200 18951
rect 8886 18885 9144 18905
rect 9196 18885 9200 18945
rect 8830 18875 9200 18885
rect 9230 19205 9600 19215
rect 9230 19145 9234 19205
rect 9286 19185 9544 19205
rect 9230 19139 9286 19145
rect 9230 18951 9260 19139
rect 9315 19130 9515 19155
rect 9596 19145 9600 19205
rect 9544 19139 9600 19145
rect 9315 19110 9385 19130
rect 9290 19070 9385 19110
rect 9445 19110 9515 19130
rect 9445 19070 9540 19110
rect 9290 19020 9540 19070
rect 9290 18980 9385 19020
rect 9315 18960 9385 18980
rect 9445 18980 9540 19020
rect 9445 18960 9515 18980
rect 9230 18945 9286 18951
rect 9230 18885 9234 18945
rect 9315 18935 9515 18960
rect 9570 18951 9600 19139
rect 9544 18945 9600 18951
rect 9286 18885 9544 18905
rect 9596 18885 9600 18945
rect 9230 18875 9600 18885
rect 9630 19205 10000 19215
rect 9630 19145 9634 19205
rect 9686 19185 9944 19205
rect 9630 19139 9686 19145
rect 9630 18951 9660 19139
rect 9715 19130 9915 19155
rect 9996 19145 10000 19205
rect 9944 19139 10000 19145
rect 9715 19110 9785 19130
rect 9690 19070 9785 19110
rect 9845 19110 9915 19130
rect 9845 19070 9940 19110
rect 9690 19020 9940 19070
rect 9690 18980 9785 19020
rect 9715 18960 9785 18980
rect 9845 18980 9940 19020
rect 9845 18960 9915 18980
rect 9630 18945 9686 18951
rect 9630 18885 9634 18945
rect 9715 18935 9915 18960
rect 9970 18951 10000 19139
rect 9944 18945 10000 18951
rect 9686 18885 9944 18905
rect 9996 18885 10000 18945
rect 9630 18875 10000 18885
rect 10030 19205 10400 19215
rect 10030 19145 10034 19205
rect 10086 19185 10344 19205
rect 10030 19139 10086 19145
rect 10030 18951 10060 19139
rect 10115 19130 10315 19155
rect 10396 19145 10400 19205
rect 10344 19139 10400 19145
rect 10115 19110 10185 19130
rect 10090 19070 10185 19110
rect 10245 19110 10315 19130
rect 10245 19070 10340 19110
rect 10090 19020 10340 19070
rect 10090 18980 10185 19020
rect 10115 18960 10185 18980
rect 10245 18980 10340 19020
rect 10245 18960 10315 18980
rect 10030 18945 10086 18951
rect 10030 18885 10034 18945
rect 10115 18935 10315 18960
rect 10370 18951 10400 19139
rect 10344 18945 10400 18951
rect 10086 18885 10344 18905
rect 10396 18885 10400 18945
rect 10030 18875 10400 18885
rect 10430 19205 10800 19215
rect 10430 19145 10434 19205
rect 10486 19185 10744 19205
rect 10430 19139 10486 19145
rect 10430 18951 10460 19139
rect 10515 19130 10715 19155
rect 10796 19145 10800 19205
rect 10744 19139 10800 19145
rect 10515 19110 10585 19130
rect 10490 19070 10585 19110
rect 10645 19110 10715 19130
rect 10645 19070 10740 19110
rect 10490 19020 10740 19070
rect 10490 18980 10585 19020
rect 10515 18960 10585 18980
rect 10645 18980 10740 19020
rect 10645 18960 10715 18980
rect 10430 18945 10486 18951
rect 10430 18885 10434 18945
rect 10515 18935 10715 18960
rect 10770 18951 10800 19139
rect 10744 18945 10800 18951
rect 10486 18885 10744 18905
rect 10796 18885 10800 18945
rect 10430 18875 10800 18885
rect 10830 19205 11200 19215
rect 10830 19145 10834 19205
rect 10886 19185 11144 19205
rect 10830 19139 10886 19145
rect 10830 18951 10860 19139
rect 10915 19130 11115 19155
rect 11196 19145 11200 19205
rect 11144 19139 11200 19145
rect 10915 19110 10985 19130
rect 10890 19070 10985 19110
rect 11045 19110 11115 19130
rect 11045 19070 11140 19110
rect 10890 19020 11140 19070
rect 10890 18980 10985 19020
rect 10915 18960 10985 18980
rect 11045 18980 11140 19020
rect 11045 18960 11115 18980
rect 10830 18945 10886 18951
rect 10830 18885 10834 18945
rect 10915 18935 11115 18960
rect 11170 18951 11200 19139
rect 11144 18945 11200 18951
rect 10886 18885 11144 18905
rect 11196 18885 11200 18945
rect 10830 18875 11200 18885
rect 11230 19205 11600 19215
rect 11230 19145 11234 19205
rect 11286 19185 11544 19205
rect 11230 19139 11286 19145
rect 11230 18951 11260 19139
rect 11315 19130 11515 19155
rect 11596 19145 11600 19205
rect 11544 19139 11600 19145
rect 11315 19110 11385 19130
rect 11290 19070 11385 19110
rect 11445 19110 11515 19130
rect 11445 19070 11540 19110
rect 11290 19020 11540 19070
rect 11290 18980 11385 19020
rect 11315 18960 11385 18980
rect 11445 18980 11540 19020
rect 11445 18960 11515 18980
rect 11230 18945 11286 18951
rect 11230 18885 11234 18945
rect 11315 18935 11515 18960
rect 11570 18951 11600 19139
rect 11544 18945 11600 18951
rect 11286 18885 11544 18905
rect 11596 18885 11600 18945
rect 11230 18875 11600 18885
rect 11630 19205 12000 19215
rect 11630 19145 11634 19205
rect 11686 19185 11944 19205
rect 11630 19139 11686 19145
rect 11630 18951 11660 19139
rect 11715 19130 11915 19155
rect 11996 19145 12000 19205
rect 11944 19139 12000 19145
rect 11715 19110 11785 19130
rect 11690 19070 11785 19110
rect 11845 19110 11915 19130
rect 11845 19070 11940 19110
rect 11690 19020 11940 19070
rect 11690 18980 11785 19020
rect 11715 18960 11785 18980
rect 11845 18980 11940 19020
rect 11845 18960 11915 18980
rect 11630 18945 11686 18951
rect 11630 18885 11634 18945
rect 11715 18935 11915 18960
rect 11970 18951 12000 19139
rect 11944 18945 12000 18951
rect 11686 18885 11944 18905
rect 11996 18885 12000 18945
rect 11630 18875 12000 18885
rect 12030 19205 12400 19215
rect 12030 19145 12034 19205
rect 12086 19185 12344 19205
rect 12030 19139 12086 19145
rect 12030 18951 12060 19139
rect 12115 19130 12315 19155
rect 12396 19145 12400 19205
rect 12344 19139 12400 19145
rect 12115 19110 12185 19130
rect 12090 19070 12185 19110
rect 12245 19110 12315 19130
rect 12245 19070 12340 19110
rect 12090 19020 12340 19070
rect 12090 18980 12185 19020
rect 12115 18960 12185 18980
rect 12245 18980 12340 19020
rect 12245 18960 12315 18980
rect 12030 18945 12086 18951
rect 12030 18885 12034 18945
rect 12115 18935 12315 18960
rect 12370 18951 12400 19139
rect 12344 18945 12400 18951
rect 12086 18885 12344 18905
rect 12396 18885 12400 18945
rect 12030 18875 12400 18885
rect 12430 19205 12800 19215
rect 12430 19145 12434 19205
rect 12486 19185 12744 19205
rect 12430 19139 12486 19145
rect 12430 18951 12460 19139
rect 12515 19130 12715 19155
rect 12796 19145 12800 19205
rect 12744 19139 12800 19145
rect 12515 19110 12585 19130
rect 12490 19070 12585 19110
rect 12645 19110 12715 19130
rect 12645 19070 12740 19110
rect 12490 19020 12740 19070
rect 12490 18980 12585 19020
rect 12515 18960 12585 18980
rect 12645 18980 12740 19020
rect 12645 18960 12715 18980
rect 12430 18945 12486 18951
rect 12430 18885 12434 18945
rect 12515 18935 12715 18960
rect 12770 18951 12800 19139
rect 12744 18945 12800 18951
rect 12486 18885 12744 18905
rect 12796 18885 12800 18945
rect 12430 18875 12800 18885
rect 12830 19205 13200 19215
rect 12830 19145 12834 19205
rect 12886 19185 13144 19205
rect 12830 19139 12886 19145
rect 12830 18951 12860 19139
rect 12915 19130 13115 19155
rect 13196 19145 13200 19205
rect 13144 19139 13200 19145
rect 12915 19110 12985 19130
rect 12890 19070 12985 19110
rect 13045 19110 13115 19130
rect 13045 19070 13140 19110
rect 12890 19020 13140 19070
rect 12890 18980 12985 19020
rect 12915 18960 12985 18980
rect 13045 18980 13140 19020
rect 13045 18960 13115 18980
rect 12830 18945 12886 18951
rect 12830 18885 12834 18945
rect 12915 18935 13115 18960
rect 13170 18951 13200 19139
rect 13144 18945 13200 18951
rect 12886 18885 13144 18905
rect 13196 18885 13200 18945
rect 12830 18875 13200 18885
rect -370 18835 0 18845
rect -370 18775 -366 18835
rect -314 18815 -56 18835
rect -370 18769 -314 18775
rect -370 18581 -340 18769
rect -285 18760 -85 18785
rect -4 18775 0 18835
rect -56 18769 0 18775
rect -285 18740 -215 18760
rect -310 18700 -215 18740
rect -155 18740 -85 18760
rect -155 18700 -60 18740
rect -310 18650 -60 18700
rect -310 18610 -215 18650
rect -285 18590 -215 18610
rect -155 18610 -60 18650
rect -155 18590 -85 18610
rect -370 18575 -314 18581
rect -370 18515 -366 18575
rect -285 18565 -85 18590
rect -30 18581 0 18769
rect -56 18575 0 18581
rect -314 18515 -56 18535
rect -4 18515 0 18575
rect -370 18505 0 18515
rect 30 18835 400 18845
rect 30 18775 34 18835
rect 86 18815 344 18835
rect 30 18769 86 18775
rect 30 18581 60 18769
rect 115 18760 315 18785
rect 396 18775 400 18835
rect 344 18769 400 18775
rect 115 18740 185 18760
rect 90 18700 185 18740
rect 245 18740 315 18760
rect 245 18700 340 18740
rect 90 18650 340 18700
rect 90 18610 185 18650
rect 115 18590 185 18610
rect 245 18610 340 18650
rect 245 18590 315 18610
rect 30 18575 86 18581
rect 30 18515 34 18575
rect 115 18565 315 18590
rect 370 18581 400 18769
rect 344 18575 400 18581
rect 86 18515 344 18535
rect 396 18515 400 18575
rect 30 18505 400 18515
rect 430 18835 800 18845
rect 430 18775 434 18835
rect 486 18815 744 18835
rect 430 18769 486 18775
rect 430 18581 460 18769
rect 515 18760 715 18785
rect 796 18775 800 18835
rect 744 18769 800 18775
rect 515 18740 585 18760
rect 490 18700 585 18740
rect 645 18740 715 18760
rect 645 18700 740 18740
rect 490 18650 740 18700
rect 490 18610 585 18650
rect 515 18590 585 18610
rect 645 18610 740 18650
rect 645 18590 715 18610
rect 430 18575 486 18581
rect 430 18515 434 18575
rect 515 18565 715 18590
rect 770 18581 800 18769
rect 744 18575 800 18581
rect 486 18515 744 18535
rect 796 18515 800 18575
rect 430 18505 800 18515
rect 830 18835 1200 18845
rect 830 18775 834 18835
rect 886 18815 1144 18835
rect 830 18769 886 18775
rect 830 18581 860 18769
rect 915 18760 1115 18785
rect 1196 18775 1200 18835
rect 1144 18769 1200 18775
rect 915 18740 985 18760
rect 890 18700 985 18740
rect 1045 18740 1115 18760
rect 1045 18700 1140 18740
rect 890 18650 1140 18700
rect 890 18610 985 18650
rect 915 18590 985 18610
rect 1045 18610 1140 18650
rect 1045 18590 1115 18610
rect 830 18575 886 18581
rect 830 18515 834 18575
rect 915 18565 1115 18590
rect 1170 18581 1200 18769
rect 1144 18575 1200 18581
rect 886 18515 1144 18535
rect 1196 18515 1200 18575
rect 830 18505 1200 18515
rect 1230 18835 1600 18845
rect 1230 18775 1234 18835
rect 1286 18815 1544 18835
rect 1230 18769 1286 18775
rect 1230 18581 1260 18769
rect 1315 18760 1515 18785
rect 1596 18775 1600 18835
rect 1544 18769 1600 18775
rect 1315 18740 1385 18760
rect 1290 18700 1385 18740
rect 1445 18740 1515 18760
rect 1445 18700 1540 18740
rect 1290 18650 1540 18700
rect 1290 18610 1385 18650
rect 1315 18590 1385 18610
rect 1445 18610 1540 18650
rect 1445 18590 1515 18610
rect 1230 18575 1286 18581
rect 1230 18515 1234 18575
rect 1315 18565 1515 18590
rect 1570 18581 1600 18769
rect 1544 18575 1600 18581
rect 1286 18515 1544 18535
rect 1596 18515 1600 18575
rect 1230 18505 1600 18515
rect 1630 18835 2000 18845
rect 1630 18775 1634 18835
rect 1686 18815 1944 18835
rect 1630 18769 1686 18775
rect 1630 18581 1660 18769
rect 1715 18760 1915 18785
rect 1996 18775 2000 18835
rect 1944 18769 2000 18775
rect 1715 18740 1785 18760
rect 1690 18700 1785 18740
rect 1845 18740 1915 18760
rect 1845 18700 1940 18740
rect 1690 18650 1940 18700
rect 1690 18610 1785 18650
rect 1715 18590 1785 18610
rect 1845 18610 1940 18650
rect 1845 18590 1915 18610
rect 1630 18575 1686 18581
rect 1630 18515 1634 18575
rect 1715 18565 1915 18590
rect 1970 18581 2000 18769
rect 1944 18575 2000 18581
rect 1686 18515 1944 18535
rect 1996 18515 2000 18575
rect 1630 18505 2000 18515
rect 2030 18835 2400 18845
rect 2030 18775 2034 18835
rect 2086 18815 2344 18835
rect 2030 18769 2086 18775
rect 2030 18581 2060 18769
rect 2115 18760 2315 18785
rect 2396 18775 2400 18835
rect 2344 18769 2400 18775
rect 2115 18740 2185 18760
rect 2090 18700 2185 18740
rect 2245 18740 2315 18760
rect 2245 18700 2340 18740
rect 2090 18650 2340 18700
rect 2090 18610 2185 18650
rect 2115 18590 2185 18610
rect 2245 18610 2340 18650
rect 2245 18590 2315 18610
rect 2030 18575 2086 18581
rect 2030 18515 2034 18575
rect 2115 18565 2315 18590
rect 2370 18581 2400 18769
rect 2344 18575 2400 18581
rect 2086 18515 2344 18535
rect 2396 18515 2400 18575
rect 2030 18505 2400 18515
rect 2430 18835 2800 18845
rect 2430 18775 2434 18835
rect 2486 18815 2744 18835
rect 2430 18769 2486 18775
rect 2430 18581 2460 18769
rect 2515 18760 2715 18785
rect 2796 18775 2800 18835
rect 2744 18769 2800 18775
rect 2515 18740 2585 18760
rect 2490 18700 2585 18740
rect 2645 18740 2715 18760
rect 2645 18700 2740 18740
rect 2490 18650 2740 18700
rect 2490 18610 2585 18650
rect 2515 18590 2585 18610
rect 2645 18610 2740 18650
rect 2645 18590 2715 18610
rect 2430 18575 2486 18581
rect 2430 18515 2434 18575
rect 2515 18565 2715 18590
rect 2770 18581 2800 18769
rect 2744 18575 2800 18581
rect 2486 18515 2744 18535
rect 2796 18515 2800 18575
rect 2430 18505 2800 18515
rect 2830 18835 3200 18845
rect 2830 18775 2834 18835
rect 2886 18815 3144 18835
rect 2830 18769 2886 18775
rect 2830 18581 2860 18769
rect 2915 18760 3115 18785
rect 3196 18775 3200 18835
rect 3144 18769 3200 18775
rect 2915 18740 2985 18760
rect 2890 18700 2985 18740
rect 3045 18740 3115 18760
rect 3045 18700 3140 18740
rect 2890 18650 3140 18700
rect 2890 18610 2985 18650
rect 2915 18590 2985 18610
rect 3045 18610 3140 18650
rect 3045 18590 3115 18610
rect 2830 18575 2886 18581
rect 2830 18515 2834 18575
rect 2915 18565 3115 18590
rect 3170 18581 3200 18769
rect 3144 18575 3200 18581
rect 2886 18515 3144 18535
rect 3196 18515 3200 18575
rect 2830 18505 3200 18515
rect 3230 18835 3600 18845
rect 3230 18775 3234 18835
rect 3286 18815 3544 18835
rect 3230 18769 3286 18775
rect 3230 18581 3260 18769
rect 3315 18760 3515 18785
rect 3596 18775 3600 18835
rect 3544 18769 3600 18775
rect 3315 18740 3385 18760
rect 3290 18700 3385 18740
rect 3445 18740 3515 18760
rect 3445 18700 3540 18740
rect 3290 18650 3540 18700
rect 3290 18610 3385 18650
rect 3315 18590 3385 18610
rect 3445 18610 3540 18650
rect 3445 18590 3515 18610
rect 3230 18575 3286 18581
rect 3230 18515 3234 18575
rect 3315 18565 3515 18590
rect 3570 18581 3600 18769
rect 3544 18575 3600 18581
rect 3286 18515 3544 18535
rect 3596 18515 3600 18575
rect 3230 18505 3600 18515
rect 3630 18835 4000 18845
rect 3630 18775 3634 18835
rect 3686 18815 3944 18835
rect 3630 18769 3686 18775
rect 3630 18581 3660 18769
rect 3715 18760 3915 18785
rect 3996 18775 4000 18835
rect 3944 18769 4000 18775
rect 3715 18740 3785 18760
rect 3690 18700 3785 18740
rect 3845 18740 3915 18760
rect 3845 18700 3940 18740
rect 3690 18650 3940 18700
rect 3690 18610 3785 18650
rect 3715 18590 3785 18610
rect 3845 18610 3940 18650
rect 3845 18590 3915 18610
rect 3630 18575 3686 18581
rect 3630 18515 3634 18575
rect 3715 18565 3915 18590
rect 3970 18581 4000 18769
rect 3944 18575 4000 18581
rect 3686 18515 3944 18535
rect 3996 18515 4000 18575
rect 3630 18505 4000 18515
rect 4030 18835 4400 18845
rect 4030 18775 4034 18835
rect 4086 18815 4344 18835
rect 4030 18769 4086 18775
rect 4030 18581 4060 18769
rect 4115 18760 4315 18785
rect 4396 18775 4400 18835
rect 4344 18769 4400 18775
rect 4115 18740 4185 18760
rect 4090 18700 4185 18740
rect 4245 18740 4315 18760
rect 4245 18700 4340 18740
rect 4090 18650 4340 18700
rect 4090 18610 4185 18650
rect 4115 18590 4185 18610
rect 4245 18610 4340 18650
rect 4245 18590 4315 18610
rect 4030 18575 4086 18581
rect 4030 18515 4034 18575
rect 4115 18565 4315 18590
rect 4370 18581 4400 18769
rect 4344 18575 4400 18581
rect 4086 18515 4344 18535
rect 4396 18515 4400 18575
rect 4030 18505 4400 18515
rect 4430 18835 4800 18845
rect 4430 18775 4434 18835
rect 4486 18815 4744 18835
rect 4430 18769 4486 18775
rect 4430 18581 4460 18769
rect 4515 18760 4715 18785
rect 4796 18775 4800 18835
rect 4744 18769 4800 18775
rect 4515 18740 4585 18760
rect 4490 18700 4585 18740
rect 4645 18740 4715 18760
rect 4645 18700 4740 18740
rect 4490 18650 4740 18700
rect 4490 18610 4585 18650
rect 4515 18590 4585 18610
rect 4645 18610 4740 18650
rect 4645 18590 4715 18610
rect 4430 18575 4486 18581
rect 4430 18515 4434 18575
rect 4515 18565 4715 18590
rect 4770 18581 4800 18769
rect 4744 18575 4800 18581
rect 4486 18515 4744 18535
rect 4796 18515 4800 18575
rect 4430 18505 4800 18515
rect 4830 18835 5200 18845
rect 4830 18775 4834 18835
rect 4886 18815 5144 18835
rect 4830 18769 4886 18775
rect 4830 18581 4860 18769
rect 4915 18760 5115 18785
rect 5196 18775 5200 18835
rect 5144 18769 5200 18775
rect 4915 18740 4985 18760
rect 4890 18700 4985 18740
rect 5045 18740 5115 18760
rect 5045 18700 5140 18740
rect 4890 18650 5140 18700
rect 4890 18610 4985 18650
rect 4915 18590 4985 18610
rect 5045 18610 5140 18650
rect 5045 18590 5115 18610
rect 4830 18575 4886 18581
rect 4830 18515 4834 18575
rect 4915 18565 5115 18590
rect 5170 18581 5200 18769
rect 5144 18575 5200 18581
rect 4886 18515 5144 18535
rect 5196 18515 5200 18575
rect 4830 18505 5200 18515
rect 5230 18835 5600 18845
rect 5230 18775 5234 18835
rect 5286 18815 5544 18835
rect 5230 18769 5286 18775
rect 5230 18581 5260 18769
rect 5315 18760 5515 18785
rect 5596 18775 5600 18835
rect 5544 18769 5600 18775
rect 5315 18740 5385 18760
rect 5290 18700 5385 18740
rect 5445 18740 5515 18760
rect 5445 18700 5540 18740
rect 5290 18650 5540 18700
rect 5290 18610 5385 18650
rect 5315 18590 5385 18610
rect 5445 18610 5540 18650
rect 5445 18590 5515 18610
rect 5230 18575 5286 18581
rect 5230 18515 5234 18575
rect 5315 18565 5515 18590
rect 5570 18581 5600 18769
rect 5544 18575 5600 18581
rect 5286 18515 5544 18535
rect 5596 18515 5600 18575
rect 5230 18505 5600 18515
rect 5630 18835 6000 18845
rect 5630 18775 5634 18835
rect 5686 18815 5944 18835
rect 5630 18769 5686 18775
rect 5630 18581 5660 18769
rect 5715 18760 5915 18785
rect 5996 18775 6000 18835
rect 5944 18769 6000 18775
rect 5715 18740 5785 18760
rect 5690 18700 5785 18740
rect 5845 18740 5915 18760
rect 5845 18700 5940 18740
rect 5690 18650 5940 18700
rect 5690 18610 5785 18650
rect 5715 18590 5785 18610
rect 5845 18610 5940 18650
rect 5845 18590 5915 18610
rect 5630 18575 5686 18581
rect 5630 18515 5634 18575
rect 5715 18565 5915 18590
rect 5970 18581 6000 18769
rect 5944 18575 6000 18581
rect 5686 18515 5944 18535
rect 5996 18515 6000 18575
rect 5630 18505 6000 18515
rect 6030 18835 6400 18845
rect 6030 18775 6034 18835
rect 6086 18815 6344 18835
rect 6030 18769 6086 18775
rect 6030 18581 6060 18769
rect 6115 18760 6315 18785
rect 6396 18775 6400 18835
rect 6344 18769 6400 18775
rect 6115 18740 6185 18760
rect 6090 18700 6185 18740
rect 6245 18740 6315 18760
rect 6245 18700 6340 18740
rect 6090 18650 6340 18700
rect 6090 18610 6185 18650
rect 6115 18590 6185 18610
rect 6245 18610 6340 18650
rect 6245 18590 6315 18610
rect 6030 18575 6086 18581
rect 6030 18515 6034 18575
rect 6115 18565 6315 18590
rect 6370 18581 6400 18769
rect 6344 18575 6400 18581
rect 6086 18515 6344 18535
rect 6396 18515 6400 18575
rect 6030 18505 6400 18515
rect 6430 18835 6800 18845
rect 6430 18775 6434 18835
rect 6486 18815 6744 18835
rect 6430 18769 6486 18775
rect 6430 18581 6460 18769
rect 6515 18760 6715 18785
rect 6796 18775 6800 18835
rect 6744 18769 6800 18775
rect 6515 18740 6585 18760
rect 6490 18700 6585 18740
rect 6645 18740 6715 18760
rect 6645 18700 6740 18740
rect 6490 18650 6740 18700
rect 6490 18610 6585 18650
rect 6515 18590 6585 18610
rect 6645 18610 6740 18650
rect 6645 18590 6715 18610
rect 6430 18575 6486 18581
rect 6430 18515 6434 18575
rect 6515 18565 6715 18590
rect 6770 18581 6800 18769
rect 6744 18575 6800 18581
rect 6486 18515 6744 18535
rect 6796 18515 6800 18575
rect 6430 18505 6800 18515
rect 6830 18835 7200 18845
rect 6830 18775 6834 18835
rect 6886 18815 7144 18835
rect 6830 18769 6886 18775
rect 6830 18581 6860 18769
rect 6915 18760 7115 18785
rect 7196 18775 7200 18835
rect 7144 18769 7200 18775
rect 6915 18740 6985 18760
rect 6890 18700 6985 18740
rect 7045 18740 7115 18760
rect 7045 18700 7140 18740
rect 6890 18650 7140 18700
rect 6890 18610 6985 18650
rect 6915 18590 6985 18610
rect 7045 18610 7140 18650
rect 7045 18590 7115 18610
rect 6830 18575 6886 18581
rect 6830 18515 6834 18575
rect 6915 18565 7115 18590
rect 7170 18581 7200 18769
rect 7144 18575 7200 18581
rect 6886 18515 7144 18535
rect 7196 18515 7200 18575
rect 6830 18505 7200 18515
rect 7230 18835 7600 18845
rect 7230 18775 7234 18835
rect 7286 18815 7544 18835
rect 7230 18769 7286 18775
rect 7230 18581 7260 18769
rect 7315 18760 7515 18785
rect 7596 18775 7600 18835
rect 7544 18769 7600 18775
rect 7315 18740 7385 18760
rect 7290 18700 7385 18740
rect 7445 18740 7515 18760
rect 7445 18700 7540 18740
rect 7290 18650 7540 18700
rect 7290 18610 7385 18650
rect 7315 18590 7385 18610
rect 7445 18610 7540 18650
rect 7445 18590 7515 18610
rect 7230 18575 7286 18581
rect 7230 18515 7234 18575
rect 7315 18565 7515 18590
rect 7570 18581 7600 18769
rect 7544 18575 7600 18581
rect 7286 18515 7544 18535
rect 7596 18515 7600 18575
rect 7230 18505 7600 18515
rect 7630 18835 8000 18845
rect 7630 18775 7634 18835
rect 7686 18815 7944 18835
rect 7630 18769 7686 18775
rect 7630 18581 7660 18769
rect 7715 18760 7915 18785
rect 7996 18775 8000 18835
rect 7944 18769 8000 18775
rect 7715 18740 7785 18760
rect 7690 18700 7785 18740
rect 7845 18740 7915 18760
rect 7845 18700 7940 18740
rect 7690 18650 7940 18700
rect 7690 18610 7785 18650
rect 7715 18590 7785 18610
rect 7845 18610 7940 18650
rect 7845 18590 7915 18610
rect 7630 18575 7686 18581
rect 7630 18515 7634 18575
rect 7715 18565 7915 18590
rect 7970 18581 8000 18769
rect 7944 18575 8000 18581
rect 7686 18515 7944 18535
rect 7996 18515 8000 18575
rect 7630 18505 8000 18515
rect 8030 18835 8400 18845
rect 8030 18775 8034 18835
rect 8086 18815 8344 18835
rect 8030 18769 8086 18775
rect 8030 18581 8060 18769
rect 8115 18760 8315 18785
rect 8396 18775 8400 18835
rect 8344 18769 8400 18775
rect 8115 18740 8185 18760
rect 8090 18700 8185 18740
rect 8245 18740 8315 18760
rect 8245 18700 8340 18740
rect 8090 18650 8340 18700
rect 8090 18610 8185 18650
rect 8115 18590 8185 18610
rect 8245 18610 8340 18650
rect 8245 18590 8315 18610
rect 8030 18575 8086 18581
rect 8030 18515 8034 18575
rect 8115 18565 8315 18590
rect 8370 18581 8400 18769
rect 8344 18575 8400 18581
rect 8086 18515 8344 18535
rect 8396 18515 8400 18575
rect 8030 18505 8400 18515
rect 8430 18835 8800 18845
rect 8430 18775 8434 18835
rect 8486 18815 8744 18835
rect 8430 18769 8486 18775
rect 8430 18581 8460 18769
rect 8515 18760 8715 18785
rect 8796 18775 8800 18835
rect 8744 18769 8800 18775
rect 8515 18740 8585 18760
rect 8490 18700 8585 18740
rect 8645 18740 8715 18760
rect 8645 18700 8740 18740
rect 8490 18650 8740 18700
rect 8490 18610 8585 18650
rect 8515 18590 8585 18610
rect 8645 18610 8740 18650
rect 8645 18590 8715 18610
rect 8430 18575 8486 18581
rect 8430 18515 8434 18575
rect 8515 18565 8715 18590
rect 8770 18581 8800 18769
rect 8744 18575 8800 18581
rect 8486 18515 8744 18535
rect 8796 18515 8800 18575
rect 8430 18505 8800 18515
rect 8830 18835 9200 18845
rect 8830 18775 8834 18835
rect 8886 18815 9144 18835
rect 8830 18769 8886 18775
rect 8830 18581 8860 18769
rect 8915 18760 9115 18785
rect 9196 18775 9200 18835
rect 9144 18769 9200 18775
rect 8915 18740 8985 18760
rect 8890 18700 8985 18740
rect 9045 18740 9115 18760
rect 9045 18700 9140 18740
rect 8890 18650 9140 18700
rect 8890 18610 8985 18650
rect 8915 18590 8985 18610
rect 9045 18610 9140 18650
rect 9045 18590 9115 18610
rect 8830 18575 8886 18581
rect 8830 18515 8834 18575
rect 8915 18565 9115 18590
rect 9170 18581 9200 18769
rect 9144 18575 9200 18581
rect 8886 18515 9144 18535
rect 9196 18515 9200 18575
rect 8830 18505 9200 18515
rect 9230 18835 9600 18845
rect 9230 18775 9234 18835
rect 9286 18815 9544 18835
rect 9230 18769 9286 18775
rect 9230 18581 9260 18769
rect 9315 18760 9515 18785
rect 9596 18775 9600 18835
rect 9544 18769 9600 18775
rect 9315 18740 9385 18760
rect 9290 18700 9385 18740
rect 9445 18740 9515 18760
rect 9445 18700 9540 18740
rect 9290 18650 9540 18700
rect 9290 18610 9385 18650
rect 9315 18590 9385 18610
rect 9445 18610 9540 18650
rect 9445 18590 9515 18610
rect 9230 18575 9286 18581
rect 9230 18515 9234 18575
rect 9315 18565 9515 18590
rect 9570 18581 9600 18769
rect 9544 18575 9600 18581
rect 9286 18515 9544 18535
rect 9596 18515 9600 18575
rect 9230 18505 9600 18515
rect 9630 18835 10000 18845
rect 9630 18775 9634 18835
rect 9686 18815 9944 18835
rect 9630 18769 9686 18775
rect 9630 18581 9660 18769
rect 9715 18760 9915 18785
rect 9996 18775 10000 18835
rect 9944 18769 10000 18775
rect 9715 18740 9785 18760
rect 9690 18700 9785 18740
rect 9845 18740 9915 18760
rect 9845 18700 9940 18740
rect 9690 18650 9940 18700
rect 9690 18610 9785 18650
rect 9715 18590 9785 18610
rect 9845 18610 9940 18650
rect 9845 18590 9915 18610
rect 9630 18575 9686 18581
rect 9630 18515 9634 18575
rect 9715 18565 9915 18590
rect 9970 18581 10000 18769
rect 9944 18575 10000 18581
rect 9686 18515 9944 18535
rect 9996 18515 10000 18575
rect 9630 18505 10000 18515
rect 10030 18835 10400 18845
rect 10030 18775 10034 18835
rect 10086 18815 10344 18835
rect 10030 18769 10086 18775
rect 10030 18581 10060 18769
rect 10115 18760 10315 18785
rect 10396 18775 10400 18835
rect 10344 18769 10400 18775
rect 10115 18740 10185 18760
rect 10090 18700 10185 18740
rect 10245 18740 10315 18760
rect 10245 18700 10340 18740
rect 10090 18650 10340 18700
rect 10090 18610 10185 18650
rect 10115 18590 10185 18610
rect 10245 18610 10340 18650
rect 10245 18590 10315 18610
rect 10030 18575 10086 18581
rect 10030 18515 10034 18575
rect 10115 18565 10315 18590
rect 10370 18581 10400 18769
rect 10344 18575 10400 18581
rect 10086 18515 10344 18535
rect 10396 18515 10400 18575
rect 10030 18505 10400 18515
rect 10430 18835 10800 18845
rect 10430 18775 10434 18835
rect 10486 18815 10744 18835
rect 10430 18769 10486 18775
rect 10430 18581 10460 18769
rect 10515 18760 10715 18785
rect 10796 18775 10800 18835
rect 10744 18769 10800 18775
rect 10515 18740 10585 18760
rect 10490 18700 10585 18740
rect 10645 18740 10715 18760
rect 10645 18700 10740 18740
rect 10490 18650 10740 18700
rect 10490 18610 10585 18650
rect 10515 18590 10585 18610
rect 10645 18610 10740 18650
rect 10645 18590 10715 18610
rect 10430 18575 10486 18581
rect 10430 18515 10434 18575
rect 10515 18565 10715 18590
rect 10770 18581 10800 18769
rect 10744 18575 10800 18581
rect 10486 18515 10744 18535
rect 10796 18515 10800 18575
rect 10430 18505 10800 18515
rect 10830 18835 11200 18845
rect 10830 18775 10834 18835
rect 10886 18815 11144 18835
rect 10830 18769 10886 18775
rect 10830 18581 10860 18769
rect 10915 18760 11115 18785
rect 11196 18775 11200 18835
rect 11144 18769 11200 18775
rect 10915 18740 10985 18760
rect 10890 18700 10985 18740
rect 11045 18740 11115 18760
rect 11045 18700 11140 18740
rect 10890 18650 11140 18700
rect 10890 18610 10985 18650
rect 10915 18590 10985 18610
rect 11045 18610 11140 18650
rect 11045 18590 11115 18610
rect 10830 18575 10886 18581
rect 10830 18515 10834 18575
rect 10915 18565 11115 18590
rect 11170 18581 11200 18769
rect 11144 18575 11200 18581
rect 10886 18515 11144 18535
rect 11196 18515 11200 18575
rect 10830 18505 11200 18515
rect 11230 18835 11600 18845
rect 11230 18775 11234 18835
rect 11286 18815 11544 18835
rect 11230 18769 11286 18775
rect 11230 18581 11260 18769
rect 11315 18760 11515 18785
rect 11596 18775 11600 18835
rect 11544 18769 11600 18775
rect 11315 18740 11385 18760
rect 11290 18700 11385 18740
rect 11445 18740 11515 18760
rect 11445 18700 11540 18740
rect 11290 18650 11540 18700
rect 11290 18610 11385 18650
rect 11315 18590 11385 18610
rect 11445 18610 11540 18650
rect 11445 18590 11515 18610
rect 11230 18575 11286 18581
rect 11230 18515 11234 18575
rect 11315 18565 11515 18590
rect 11570 18581 11600 18769
rect 11544 18575 11600 18581
rect 11286 18515 11544 18535
rect 11596 18515 11600 18575
rect 11230 18505 11600 18515
rect 11630 18835 12000 18845
rect 11630 18775 11634 18835
rect 11686 18815 11944 18835
rect 11630 18769 11686 18775
rect 11630 18581 11660 18769
rect 11715 18760 11915 18785
rect 11996 18775 12000 18835
rect 11944 18769 12000 18775
rect 11715 18740 11785 18760
rect 11690 18700 11785 18740
rect 11845 18740 11915 18760
rect 11845 18700 11940 18740
rect 11690 18650 11940 18700
rect 11690 18610 11785 18650
rect 11715 18590 11785 18610
rect 11845 18610 11940 18650
rect 11845 18590 11915 18610
rect 11630 18575 11686 18581
rect 11630 18515 11634 18575
rect 11715 18565 11915 18590
rect 11970 18581 12000 18769
rect 11944 18575 12000 18581
rect 11686 18515 11944 18535
rect 11996 18515 12000 18575
rect 11630 18505 12000 18515
rect 12030 18835 12400 18845
rect 12030 18775 12034 18835
rect 12086 18815 12344 18835
rect 12030 18769 12086 18775
rect 12030 18581 12060 18769
rect 12115 18760 12315 18785
rect 12396 18775 12400 18835
rect 12344 18769 12400 18775
rect 12115 18740 12185 18760
rect 12090 18700 12185 18740
rect 12245 18740 12315 18760
rect 12245 18700 12340 18740
rect 12090 18650 12340 18700
rect 12090 18610 12185 18650
rect 12115 18590 12185 18610
rect 12245 18610 12340 18650
rect 12245 18590 12315 18610
rect 12030 18575 12086 18581
rect 12030 18515 12034 18575
rect 12115 18565 12315 18590
rect 12370 18581 12400 18769
rect 12344 18575 12400 18581
rect 12086 18515 12344 18535
rect 12396 18515 12400 18575
rect 12030 18505 12400 18515
rect 12430 18835 12800 18845
rect 12430 18775 12434 18835
rect 12486 18815 12744 18835
rect 12430 18769 12486 18775
rect 12430 18581 12460 18769
rect 12515 18760 12715 18785
rect 12796 18775 12800 18835
rect 12744 18769 12800 18775
rect 12515 18740 12585 18760
rect 12490 18700 12585 18740
rect 12645 18740 12715 18760
rect 12645 18700 12740 18740
rect 12490 18650 12740 18700
rect 12490 18610 12585 18650
rect 12515 18590 12585 18610
rect 12645 18610 12740 18650
rect 12645 18590 12715 18610
rect 12430 18575 12486 18581
rect 12430 18515 12434 18575
rect 12515 18565 12715 18590
rect 12770 18581 12800 18769
rect 12744 18575 12800 18581
rect 12486 18515 12744 18535
rect 12796 18515 12800 18575
rect 12430 18505 12800 18515
rect 12830 18835 13200 18845
rect 12830 18775 12834 18835
rect 12886 18815 13144 18835
rect 12830 18769 12886 18775
rect 12830 18581 12860 18769
rect 12915 18760 13115 18785
rect 13196 18775 13200 18835
rect 13144 18769 13200 18775
rect 12915 18740 12985 18760
rect 12890 18700 12985 18740
rect 13045 18740 13115 18760
rect 13045 18700 13140 18740
rect 12890 18650 13140 18700
rect 12890 18610 12985 18650
rect 12915 18590 12985 18610
rect 13045 18610 13140 18650
rect 13045 18590 13115 18610
rect 12830 18575 12886 18581
rect 12830 18515 12834 18575
rect 12915 18565 13115 18590
rect 13170 18581 13200 18769
rect 13144 18575 13200 18581
rect 12886 18515 13144 18535
rect 13196 18515 13200 18575
rect 12830 18505 13200 18515
rect -370 18465 0 18475
rect -370 18405 -366 18465
rect -314 18445 -56 18465
rect -370 18399 -314 18405
rect -370 18211 -340 18399
rect -285 18390 -85 18415
rect -4 18405 0 18465
rect -56 18399 0 18405
rect -285 18370 -215 18390
rect -310 18330 -215 18370
rect -155 18370 -85 18390
rect -155 18330 -60 18370
rect -310 18280 -60 18330
rect -310 18240 -215 18280
rect -285 18220 -215 18240
rect -155 18240 -60 18280
rect -155 18220 -85 18240
rect -370 18205 -314 18211
rect -370 18145 -366 18205
rect -285 18195 -85 18220
rect -30 18211 0 18399
rect -56 18205 0 18211
rect -314 18145 -56 18165
rect -4 18145 0 18205
rect -370 18135 0 18145
rect 30 18465 400 18475
rect 30 18405 34 18465
rect 86 18445 344 18465
rect 30 18399 86 18405
rect 30 18211 60 18399
rect 115 18390 315 18415
rect 396 18405 400 18465
rect 344 18399 400 18405
rect 115 18370 185 18390
rect 90 18330 185 18370
rect 245 18370 315 18390
rect 245 18330 340 18370
rect 90 18280 340 18330
rect 90 18240 185 18280
rect 115 18220 185 18240
rect 245 18240 340 18280
rect 245 18220 315 18240
rect 30 18205 86 18211
rect 30 18145 34 18205
rect 115 18195 315 18220
rect 370 18211 400 18399
rect 344 18205 400 18211
rect 86 18145 344 18165
rect 396 18145 400 18205
rect 30 18135 400 18145
rect 430 18465 800 18475
rect 430 18405 434 18465
rect 486 18445 744 18465
rect 430 18399 486 18405
rect 430 18211 460 18399
rect 515 18390 715 18415
rect 796 18405 800 18465
rect 744 18399 800 18405
rect 515 18370 585 18390
rect 490 18330 585 18370
rect 645 18370 715 18390
rect 645 18330 740 18370
rect 490 18280 740 18330
rect 490 18240 585 18280
rect 515 18220 585 18240
rect 645 18240 740 18280
rect 645 18220 715 18240
rect 430 18205 486 18211
rect 430 18145 434 18205
rect 515 18195 715 18220
rect 770 18211 800 18399
rect 744 18205 800 18211
rect 486 18145 744 18165
rect 796 18145 800 18205
rect 430 18135 800 18145
rect 830 18465 1200 18475
rect 830 18405 834 18465
rect 886 18445 1144 18465
rect 830 18399 886 18405
rect 830 18211 860 18399
rect 915 18390 1115 18415
rect 1196 18405 1200 18465
rect 1144 18399 1200 18405
rect 915 18370 985 18390
rect 890 18330 985 18370
rect 1045 18370 1115 18390
rect 1045 18330 1140 18370
rect 890 18280 1140 18330
rect 890 18240 985 18280
rect 915 18220 985 18240
rect 1045 18240 1140 18280
rect 1045 18220 1115 18240
rect 830 18205 886 18211
rect 830 18145 834 18205
rect 915 18195 1115 18220
rect 1170 18211 1200 18399
rect 1144 18205 1200 18211
rect 886 18145 1144 18165
rect 1196 18145 1200 18205
rect 830 18135 1200 18145
rect 1230 18465 1600 18475
rect 1230 18405 1234 18465
rect 1286 18445 1544 18465
rect 1230 18399 1286 18405
rect 1230 18211 1260 18399
rect 1315 18390 1515 18415
rect 1596 18405 1600 18465
rect 1544 18399 1600 18405
rect 1315 18370 1385 18390
rect 1290 18330 1385 18370
rect 1445 18370 1515 18390
rect 1445 18330 1540 18370
rect 1290 18280 1540 18330
rect 1290 18240 1385 18280
rect 1315 18220 1385 18240
rect 1445 18240 1540 18280
rect 1445 18220 1515 18240
rect 1230 18205 1286 18211
rect 1230 18145 1234 18205
rect 1315 18195 1515 18220
rect 1570 18211 1600 18399
rect 1544 18205 1600 18211
rect 1286 18145 1544 18165
rect 1596 18145 1600 18205
rect 1230 18135 1600 18145
rect 1630 18465 2000 18475
rect 1630 18405 1634 18465
rect 1686 18445 1944 18465
rect 1630 18399 1686 18405
rect 1630 18211 1660 18399
rect 1715 18390 1915 18415
rect 1996 18405 2000 18465
rect 1944 18399 2000 18405
rect 1715 18370 1785 18390
rect 1690 18330 1785 18370
rect 1845 18370 1915 18390
rect 1845 18330 1940 18370
rect 1690 18280 1940 18330
rect 1690 18240 1785 18280
rect 1715 18220 1785 18240
rect 1845 18240 1940 18280
rect 1845 18220 1915 18240
rect 1630 18205 1686 18211
rect 1630 18145 1634 18205
rect 1715 18195 1915 18220
rect 1970 18211 2000 18399
rect 1944 18205 2000 18211
rect 1686 18145 1944 18165
rect 1996 18145 2000 18205
rect 1630 18135 2000 18145
rect 2030 18465 2400 18475
rect 2030 18405 2034 18465
rect 2086 18445 2344 18465
rect 2030 18399 2086 18405
rect 2030 18211 2060 18399
rect 2115 18390 2315 18415
rect 2396 18405 2400 18465
rect 2344 18399 2400 18405
rect 2115 18370 2185 18390
rect 2090 18330 2185 18370
rect 2245 18370 2315 18390
rect 2245 18330 2340 18370
rect 2090 18280 2340 18330
rect 2090 18240 2185 18280
rect 2115 18220 2185 18240
rect 2245 18240 2340 18280
rect 2245 18220 2315 18240
rect 2030 18205 2086 18211
rect 2030 18145 2034 18205
rect 2115 18195 2315 18220
rect 2370 18211 2400 18399
rect 2344 18205 2400 18211
rect 2086 18145 2344 18165
rect 2396 18145 2400 18205
rect 2030 18135 2400 18145
rect 2430 18465 2800 18475
rect 2430 18405 2434 18465
rect 2486 18445 2744 18465
rect 2430 18399 2486 18405
rect 2430 18211 2460 18399
rect 2515 18390 2715 18415
rect 2796 18405 2800 18465
rect 2744 18399 2800 18405
rect 2515 18370 2585 18390
rect 2490 18330 2585 18370
rect 2645 18370 2715 18390
rect 2645 18330 2740 18370
rect 2490 18280 2740 18330
rect 2490 18240 2585 18280
rect 2515 18220 2585 18240
rect 2645 18240 2740 18280
rect 2645 18220 2715 18240
rect 2430 18205 2486 18211
rect 2430 18145 2434 18205
rect 2515 18195 2715 18220
rect 2770 18211 2800 18399
rect 2744 18205 2800 18211
rect 2486 18145 2744 18165
rect 2796 18145 2800 18205
rect 2430 18135 2800 18145
rect 2830 18465 3200 18475
rect 2830 18405 2834 18465
rect 2886 18445 3144 18465
rect 2830 18399 2886 18405
rect 2830 18211 2860 18399
rect 2915 18390 3115 18415
rect 3196 18405 3200 18465
rect 3144 18399 3200 18405
rect 2915 18370 2985 18390
rect 2890 18330 2985 18370
rect 3045 18370 3115 18390
rect 3045 18330 3140 18370
rect 2890 18280 3140 18330
rect 2890 18240 2985 18280
rect 2915 18220 2985 18240
rect 3045 18240 3140 18280
rect 3045 18220 3115 18240
rect 2830 18205 2886 18211
rect 2830 18145 2834 18205
rect 2915 18195 3115 18220
rect 3170 18211 3200 18399
rect 3144 18205 3200 18211
rect 2886 18145 3144 18165
rect 3196 18145 3200 18205
rect 2830 18135 3200 18145
rect 3230 18465 3600 18475
rect 3230 18405 3234 18465
rect 3286 18445 3544 18465
rect 3230 18399 3286 18405
rect 3230 18211 3260 18399
rect 3315 18390 3515 18415
rect 3596 18405 3600 18465
rect 3544 18399 3600 18405
rect 3315 18370 3385 18390
rect 3290 18330 3385 18370
rect 3445 18370 3515 18390
rect 3445 18330 3540 18370
rect 3290 18280 3540 18330
rect 3290 18240 3385 18280
rect 3315 18220 3385 18240
rect 3445 18240 3540 18280
rect 3445 18220 3515 18240
rect 3230 18205 3286 18211
rect 3230 18145 3234 18205
rect 3315 18195 3515 18220
rect 3570 18211 3600 18399
rect 3544 18205 3600 18211
rect 3286 18145 3544 18165
rect 3596 18145 3600 18205
rect 3230 18135 3600 18145
rect 3630 18465 4000 18475
rect 3630 18405 3634 18465
rect 3686 18445 3944 18465
rect 3630 18399 3686 18405
rect 3630 18211 3660 18399
rect 3715 18390 3915 18415
rect 3996 18405 4000 18465
rect 3944 18399 4000 18405
rect 3715 18370 3785 18390
rect 3690 18330 3785 18370
rect 3845 18370 3915 18390
rect 3845 18330 3940 18370
rect 3690 18280 3940 18330
rect 3690 18240 3785 18280
rect 3715 18220 3785 18240
rect 3845 18240 3940 18280
rect 3845 18220 3915 18240
rect 3630 18205 3686 18211
rect 3630 18145 3634 18205
rect 3715 18195 3915 18220
rect 3970 18211 4000 18399
rect 3944 18205 4000 18211
rect 3686 18145 3944 18165
rect 3996 18145 4000 18205
rect 3630 18135 4000 18145
rect 4030 18465 4400 18475
rect 4030 18405 4034 18465
rect 4086 18445 4344 18465
rect 4030 18399 4086 18405
rect 4030 18211 4060 18399
rect 4115 18390 4315 18415
rect 4396 18405 4400 18465
rect 4344 18399 4400 18405
rect 4115 18370 4185 18390
rect 4090 18330 4185 18370
rect 4245 18370 4315 18390
rect 4245 18330 4340 18370
rect 4090 18280 4340 18330
rect 4090 18240 4185 18280
rect 4115 18220 4185 18240
rect 4245 18240 4340 18280
rect 4245 18220 4315 18240
rect 4030 18205 4086 18211
rect 4030 18145 4034 18205
rect 4115 18195 4315 18220
rect 4370 18211 4400 18399
rect 4344 18205 4400 18211
rect 4086 18145 4344 18165
rect 4396 18145 4400 18205
rect 4030 18135 4400 18145
rect 4430 18465 4800 18475
rect 4430 18405 4434 18465
rect 4486 18445 4744 18465
rect 4430 18399 4486 18405
rect 4430 18211 4460 18399
rect 4515 18390 4715 18415
rect 4796 18405 4800 18465
rect 4744 18399 4800 18405
rect 4515 18370 4585 18390
rect 4490 18330 4585 18370
rect 4645 18370 4715 18390
rect 4645 18330 4740 18370
rect 4490 18280 4740 18330
rect 4490 18240 4585 18280
rect 4515 18220 4585 18240
rect 4645 18240 4740 18280
rect 4645 18220 4715 18240
rect 4430 18205 4486 18211
rect 4430 18145 4434 18205
rect 4515 18195 4715 18220
rect 4770 18211 4800 18399
rect 4744 18205 4800 18211
rect 4486 18145 4744 18165
rect 4796 18145 4800 18205
rect 4430 18135 4800 18145
rect 4830 18465 5200 18475
rect 4830 18405 4834 18465
rect 4886 18445 5144 18465
rect 4830 18399 4886 18405
rect 4830 18211 4860 18399
rect 4915 18390 5115 18415
rect 5196 18405 5200 18465
rect 5144 18399 5200 18405
rect 4915 18370 4985 18390
rect 4890 18330 4985 18370
rect 5045 18370 5115 18390
rect 5045 18330 5140 18370
rect 4890 18280 5140 18330
rect 4890 18240 4985 18280
rect 4915 18220 4985 18240
rect 5045 18240 5140 18280
rect 5045 18220 5115 18240
rect 4830 18205 4886 18211
rect 4830 18145 4834 18205
rect 4915 18195 5115 18220
rect 5170 18211 5200 18399
rect 5144 18205 5200 18211
rect 4886 18145 5144 18165
rect 5196 18145 5200 18205
rect 4830 18135 5200 18145
rect 5230 18465 5600 18475
rect 5230 18405 5234 18465
rect 5286 18445 5544 18465
rect 5230 18399 5286 18405
rect 5230 18211 5260 18399
rect 5315 18390 5515 18415
rect 5596 18405 5600 18465
rect 5544 18399 5600 18405
rect 5315 18370 5385 18390
rect 5290 18330 5385 18370
rect 5445 18370 5515 18390
rect 5445 18330 5540 18370
rect 5290 18280 5540 18330
rect 5290 18240 5385 18280
rect 5315 18220 5385 18240
rect 5445 18240 5540 18280
rect 5445 18220 5515 18240
rect 5230 18205 5286 18211
rect 5230 18145 5234 18205
rect 5315 18195 5515 18220
rect 5570 18211 5600 18399
rect 5544 18205 5600 18211
rect 5286 18145 5544 18165
rect 5596 18145 5600 18205
rect 5230 18135 5600 18145
rect 5630 18465 6000 18475
rect 5630 18405 5634 18465
rect 5686 18445 5944 18465
rect 5630 18399 5686 18405
rect 5630 18211 5660 18399
rect 5715 18390 5915 18415
rect 5996 18405 6000 18465
rect 5944 18399 6000 18405
rect 5715 18370 5785 18390
rect 5690 18330 5785 18370
rect 5845 18370 5915 18390
rect 5845 18330 5940 18370
rect 5690 18280 5940 18330
rect 5690 18240 5785 18280
rect 5715 18220 5785 18240
rect 5845 18240 5940 18280
rect 5845 18220 5915 18240
rect 5630 18205 5686 18211
rect 5630 18145 5634 18205
rect 5715 18195 5915 18220
rect 5970 18211 6000 18399
rect 5944 18205 6000 18211
rect 5686 18145 5944 18165
rect 5996 18145 6000 18205
rect 5630 18135 6000 18145
rect 6030 18465 6400 18475
rect 6030 18405 6034 18465
rect 6086 18445 6344 18465
rect 6030 18399 6086 18405
rect 6030 18211 6060 18399
rect 6115 18390 6315 18415
rect 6396 18405 6400 18465
rect 6344 18399 6400 18405
rect 6115 18370 6185 18390
rect 6090 18330 6185 18370
rect 6245 18370 6315 18390
rect 6245 18330 6340 18370
rect 6090 18280 6340 18330
rect 6090 18240 6185 18280
rect 6115 18220 6185 18240
rect 6245 18240 6340 18280
rect 6245 18220 6315 18240
rect 6030 18205 6086 18211
rect 6030 18145 6034 18205
rect 6115 18195 6315 18220
rect 6370 18211 6400 18399
rect 6344 18205 6400 18211
rect 6086 18145 6344 18165
rect 6396 18145 6400 18205
rect 6030 18135 6400 18145
rect 6430 18465 6800 18475
rect 6430 18405 6434 18465
rect 6486 18445 6744 18465
rect 6430 18399 6486 18405
rect 6430 18211 6460 18399
rect 6515 18390 6715 18415
rect 6796 18405 6800 18465
rect 6744 18399 6800 18405
rect 6515 18370 6585 18390
rect 6490 18330 6585 18370
rect 6645 18370 6715 18390
rect 6645 18330 6740 18370
rect 6490 18280 6740 18330
rect 6490 18240 6585 18280
rect 6515 18220 6585 18240
rect 6645 18240 6740 18280
rect 6645 18220 6715 18240
rect 6430 18205 6486 18211
rect 6430 18145 6434 18205
rect 6515 18195 6715 18220
rect 6770 18211 6800 18399
rect 6744 18205 6800 18211
rect 6486 18145 6744 18165
rect 6796 18145 6800 18205
rect 6430 18135 6800 18145
rect 6830 18465 7200 18475
rect 6830 18405 6834 18465
rect 6886 18445 7144 18465
rect 6830 18399 6886 18405
rect 6830 18211 6860 18399
rect 6915 18390 7115 18415
rect 7196 18405 7200 18465
rect 7144 18399 7200 18405
rect 6915 18370 6985 18390
rect 6890 18330 6985 18370
rect 7045 18370 7115 18390
rect 7045 18330 7140 18370
rect 6890 18280 7140 18330
rect 6890 18240 6985 18280
rect 6915 18220 6985 18240
rect 7045 18240 7140 18280
rect 7045 18220 7115 18240
rect 6830 18205 6886 18211
rect 6830 18145 6834 18205
rect 6915 18195 7115 18220
rect 7170 18211 7200 18399
rect 7144 18205 7200 18211
rect 6886 18145 7144 18165
rect 7196 18145 7200 18205
rect 6830 18135 7200 18145
rect 7230 18465 7600 18475
rect 7230 18405 7234 18465
rect 7286 18445 7544 18465
rect 7230 18399 7286 18405
rect 7230 18211 7260 18399
rect 7315 18390 7515 18415
rect 7596 18405 7600 18465
rect 7544 18399 7600 18405
rect 7315 18370 7385 18390
rect 7290 18330 7385 18370
rect 7445 18370 7515 18390
rect 7445 18330 7540 18370
rect 7290 18280 7540 18330
rect 7290 18240 7385 18280
rect 7315 18220 7385 18240
rect 7445 18240 7540 18280
rect 7445 18220 7515 18240
rect 7230 18205 7286 18211
rect 7230 18145 7234 18205
rect 7315 18195 7515 18220
rect 7570 18211 7600 18399
rect 7544 18205 7600 18211
rect 7286 18145 7544 18165
rect 7596 18145 7600 18205
rect 7230 18135 7600 18145
rect 7630 18465 8000 18475
rect 7630 18405 7634 18465
rect 7686 18445 7944 18465
rect 7630 18399 7686 18405
rect 7630 18211 7660 18399
rect 7715 18390 7915 18415
rect 7996 18405 8000 18465
rect 7944 18399 8000 18405
rect 7715 18370 7785 18390
rect 7690 18330 7785 18370
rect 7845 18370 7915 18390
rect 7845 18330 7940 18370
rect 7690 18280 7940 18330
rect 7690 18240 7785 18280
rect 7715 18220 7785 18240
rect 7845 18240 7940 18280
rect 7845 18220 7915 18240
rect 7630 18205 7686 18211
rect 7630 18145 7634 18205
rect 7715 18195 7915 18220
rect 7970 18211 8000 18399
rect 7944 18205 8000 18211
rect 7686 18145 7944 18165
rect 7996 18145 8000 18205
rect 7630 18135 8000 18145
rect 8030 18465 8400 18475
rect 8030 18405 8034 18465
rect 8086 18445 8344 18465
rect 8030 18399 8086 18405
rect 8030 18211 8060 18399
rect 8115 18390 8315 18415
rect 8396 18405 8400 18465
rect 8344 18399 8400 18405
rect 8115 18370 8185 18390
rect 8090 18330 8185 18370
rect 8245 18370 8315 18390
rect 8245 18330 8340 18370
rect 8090 18280 8340 18330
rect 8090 18240 8185 18280
rect 8115 18220 8185 18240
rect 8245 18240 8340 18280
rect 8245 18220 8315 18240
rect 8030 18205 8086 18211
rect 8030 18145 8034 18205
rect 8115 18195 8315 18220
rect 8370 18211 8400 18399
rect 8344 18205 8400 18211
rect 8086 18145 8344 18165
rect 8396 18145 8400 18205
rect 8030 18135 8400 18145
rect 8430 18465 8800 18475
rect 8430 18405 8434 18465
rect 8486 18445 8744 18465
rect 8430 18399 8486 18405
rect 8430 18211 8460 18399
rect 8515 18390 8715 18415
rect 8796 18405 8800 18465
rect 8744 18399 8800 18405
rect 8515 18370 8585 18390
rect 8490 18330 8585 18370
rect 8645 18370 8715 18390
rect 8645 18330 8740 18370
rect 8490 18280 8740 18330
rect 8490 18240 8585 18280
rect 8515 18220 8585 18240
rect 8645 18240 8740 18280
rect 8645 18220 8715 18240
rect 8430 18205 8486 18211
rect 8430 18145 8434 18205
rect 8515 18195 8715 18220
rect 8770 18211 8800 18399
rect 8744 18205 8800 18211
rect 8486 18145 8744 18165
rect 8796 18145 8800 18205
rect 8430 18135 8800 18145
rect 8830 18465 9200 18475
rect 8830 18405 8834 18465
rect 8886 18445 9144 18465
rect 8830 18399 8886 18405
rect 8830 18211 8860 18399
rect 8915 18390 9115 18415
rect 9196 18405 9200 18465
rect 9144 18399 9200 18405
rect 8915 18370 8985 18390
rect 8890 18330 8985 18370
rect 9045 18370 9115 18390
rect 9045 18330 9140 18370
rect 8890 18280 9140 18330
rect 8890 18240 8985 18280
rect 8915 18220 8985 18240
rect 9045 18240 9140 18280
rect 9045 18220 9115 18240
rect 8830 18205 8886 18211
rect 8830 18145 8834 18205
rect 8915 18195 9115 18220
rect 9170 18211 9200 18399
rect 9144 18205 9200 18211
rect 8886 18145 9144 18165
rect 9196 18145 9200 18205
rect 8830 18135 9200 18145
rect 9230 18465 9600 18475
rect 9230 18405 9234 18465
rect 9286 18445 9544 18465
rect 9230 18399 9286 18405
rect 9230 18211 9260 18399
rect 9315 18390 9515 18415
rect 9596 18405 9600 18465
rect 9544 18399 9600 18405
rect 9315 18370 9385 18390
rect 9290 18330 9385 18370
rect 9445 18370 9515 18390
rect 9445 18330 9540 18370
rect 9290 18280 9540 18330
rect 9290 18240 9385 18280
rect 9315 18220 9385 18240
rect 9445 18240 9540 18280
rect 9445 18220 9515 18240
rect 9230 18205 9286 18211
rect 9230 18145 9234 18205
rect 9315 18195 9515 18220
rect 9570 18211 9600 18399
rect 9544 18205 9600 18211
rect 9286 18145 9544 18165
rect 9596 18145 9600 18205
rect 9230 18135 9600 18145
rect 9630 18465 10000 18475
rect 9630 18405 9634 18465
rect 9686 18445 9944 18465
rect 9630 18399 9686 18405
rect 9630 18211 9660 18399
rect 9715 18390 9915 18415
rect 9996 18405 10000 18465
rect 9944 18399 10000 18405
rect 9715 18370 9785 18390
rect 9690 18330 9785 18370
rect 9845 18370 9915 18390
rect 9845 18330 9940 18370
rect 9690 18280 9940 18330
rect 9690 18240 9785 18280
rect 9715 18220 9785 18240
rect 9845 18240 9940 18280
rect 9845 18220 9915 18240
rect 9630 18205 9686 18211
rect 9630 18145 9634 18205
rect 9715 18195 9915 18220
rect 9970 18211 10000 18399
rect 9944 18205 10000 18211
rect 9686 18145 9944 18165
rect 9996 18145 10000 18205
rect 9630 18135 10000 18145
rect 10030 18465 10400 18475
rect 10030 18405 10034 18465
rect 10086 18445 10344 18465
rect 10030 18399 10086 18405
rect 10030 18211 10060 18399
rect 10115 18390 10315 18415
rect 10396 18405 10400 18465
rect 10344 18399 10400 18405
rect 10115 18370 10185 18390
rect 10090 18330 10185 18370
rect 10245 18370 10315 18390
rect 10245 18330 10340 18370
rect 10090 18280 10340 18330
rect 10090 18240 10185 18280
rect 10115 18220 10185 18240
rect 10245 18240 10340 18280
rect 10245 18220 10315 18240
rect 10030 18205 10086 18211
rect 10030 18145 10034 18205
rect 10115 18195 10315 18220
rect 10370 18211 10400 18399
rect 10344 18205 10400 18211
rect 10086 18145 10344 18165
rect 10396 18145 10400 18205
rect 10030 18135 10400 18145
rect 10430 18465 10800 18475
rect 10430 18405 10434 18465
rect 10486 18445 10744 18465
rect 10430 18399 10486 18405
rect 10430 18211 10460 18399
rect 10515 18390 10715 18415
rect 10796 18405 10800 18465
rect 10744 18399 10800 18405
rect 10515 18370 10585 18390
rect 10490 18330 10585 18370
rect 10645 18370 10715 18390
rect 10645 18330 10740 18370
rect 10490 18280 10740 18330
rect 10490 18240 10585 18280
rect 10515 18220 10585 18240
rect 10645 18240 10740 18280
rect 10645 18220 10715 18240
rect 10430 18205 10486 18211
rect 10430 18145 10434 18205
rect 10515 18195 10715 18220
rect 10770 18211 10800 18399
rect 10744 18205 10800 18211
rect 10486 18145 10744 18165
rect 10796 18145 10800 18205
rect 10430 18135 10800 18145
rect 10830 18465 11200 18475
rect 10830 18405 10834 18465
rect 10886 18445 11144 18465
rect 10830 18399 10886 18405
rect 10830 18211 10860 18399
rect 10915 18390 11115 18415
rect 11196 18405 11200 18465
rect 11144 18399 11200 18405
rect 10915 18370 10985 18390
rect 10890 18330 10985 18370
rect 11045 18370 11115 18390
rect 11045 18330 11140 18370
rect 10890 18280 11140 18330
rect 10890 18240 10985 18280
rect 10915 18220 10985 18240
rect 11045 18240 11140 18280
rect 11045 18220 11115 18240
rect 10830 18205 10886 18211
rect 10830 18145 10834 18205
rect 10915 18195 11115 18220
rect 11170 18211 11200 18399
rect 11144 18205 11200 18211
rect 10886 18145 11144 18165
rect 11196 18145 11200 18205
rect 10830 18135 11200 18145
rect 11230 18465 11600 18475
rect 11230 18405 11234 18465
rect 11286 18445 11544 18465
rect 11230 18399 11286 18405
rect 11230 18211 11260 18399
rect 11315 18390 11515 18415
rect 11596 18405 11600 18465
rect 11544 18399 11600 18405
rect 11315 18370 11385 18390
rect 11290 18330 11385 18370
rect 11445 18370 11515 18390
rect 11445 18330 11540 18370
rect 11290 18280 11540 18330
rect 11290 18240 11385 18280
rect 11315 18220 11385 18240
rect 11445 18240 11540 18280
rect 11445 18220 11515 18240
rect 11230 18205 11286 18211
rect 11230 18145 11234 18205
rect 11315 18195 11515 18220
rect 11570 18211 11600 18399
rect 11544 18205 11600 18211
rect 11286 18145 11544 18165
rect 11596 18145 11600 18205
rect 11230 18135 11600 18145
rect 11630 18465 12000 18475
rect 11630 18405 11634 18465
rect 11686 18445 11944 18465
rect 11630 18399 11686 18405
rect 11630 18211 11660 18399
rect 11715 18390 11915 18415
rect 11996 18405 12000 18465
rect 11944 18399 12000 18405
rect 11715 18370 11785 18390
rect 11690 18330 11785 18370
rect 11845 18370 11915 18390
rect 11845 18330 11940 18370
rect 11690 18280 11940 18330
rect 11690 18240 11785 18280
rect 11715 18220 11785 18240
rect 11845 18240 11940 18280
rect 11845 18220 11915 18240
rect 11630 18205 11686 18211
rect 11630 18145 11634 18205
rect 11715 18195 11915 18220
rect 11970 18211 12000 18399
rect 11944 18205 12000 18211
rect 11686 18145 11944 18165
rect 11996 18145 12000 18205
rect 11630 18135 12000 18145
rect 12030 18465 12400 18475
rect 12030 18405 12034 18465
rect 12086 18445 12344 18465
rect 12030 18399 12086 18405
rect 12030 18211 12060 18399
rect 12115 18390 12315 18415
rect 12396 18405 12400 18465
rect 12344 18399 12400 18405
rect 12115 18370 12185 18390
rect 12090 18330 12185 18370
rect 12245 18370 12315 18390
rect 12245 18330 12340 18370
rect 12090 18280 12340 18330
rect 12090 18240 12185 18280
rect 12115 18220 12185 18240
rect 12245 18240 12340 18280
rect 12245 18220 12315 18240
rect 12030 18205 12086 18211
rect 12030 18145 12034 18205
rect 12115 18195 12315 18220
rect 12370 18211 12400 18399
rect 12344 18205 12400 18211
rect 12086 18145 12344 18165
rect 12396 18145 12400 18205
rect 12030 18135 12400 18145
rect 12430 18465 12800 18475
rect 12430 18405 12434 18465
rect 12486 18445 12744 18465
rect 12430 18399 12486 18405
rect 12430 18211 12460 18399
rect 12515 18390 12715 18415
rect 12796 18405 12800 18465
rect 12744 18399 12800 18405
rect 12515 18370 12585 18390
rect 12490 18330 12585 18370
rect 12645 18370 12715 18390
rect 12645 18330 12740 18370
rect 12490 18280 12740 18330
rect 12490 18240 12585 18280
rect 12515 18220 12585 18240
rect 12645 18240 12740 18280
rect 12645 18220 12715 18240
rect 12430 18205 12486 18211
rect 12430 18145 12434 18205
rect 12515 18195 12715 18220
rect 12770 18211 12800 18399
rect 12744 18205 12800 18211
rect 12486 18145 12744 18165
rect 12796 18145 12800 18205
rect 12430 18135 12800 18145
rect 12830 18465 13200 18475
rect 12830 18405 12834 18465
rect 12886 18445 13144 18465
rect 12830 18399 12886 18405
rect 12830 18211 12860 18399
rect 12915 18390 13115 18415
rect 13196 18405 13200 18465
rect 13144 18399 13200 18405
rect 12915 18370 12985 18390
rect 12890 18330 12985 18370
rect 13045 18370 13115 18390
rect 13045 18330 13140 18370
rect 12890 18280 13140 18330
rect 12890 18240 12985 18280
rect 12915 18220 12985 18240
rect 13045 18240 13140 18280
rect 13045 18220 13115 18240
rect 12830 18205 12886 18211
rect 12830 18145 12834 18205
rect 12915 18195 13115 18220
rect 13170 18211 13200 18399
rect 13144 18205 13200 18211
rect 12886 18145 13144 18165
rect 13196 18145 13200 18205
rect 12830 18135 13200 18145
rect -370 18095 0 18105
rect -370 18035 -366 18095
rect -314 18075 -56 18095
rect -370 18029 -314 18035
rect -370 17841 -340 18029
rect -285 18020 -85 18045
rect -4 18035 0 18095
rect -56 18029 0 18035
rect -285 18000 -215 18020
rect -310 17960 -215 18000
rect -155 18000 -85 18020
rect -155 17960 -60 18000
rect -310 17910 -60 17960
rect -310 17870 -215 17910
rect -285 17850 -215 17870
rect -155 17870 -60 17910
rect -155 17850 -85 17870
rect -370 17835 -314 17841
rect -370 17775 -366 17835
rect -285 17825 -85 17850
rect -30 17841 0 18029
rect -56 17835 0 17841
rect -314 17775 -56 17795
rect -4 17775 0 17835
rect -370 17765 0 17775
rect 30 18095 400 18105
rect 30 18035 34 18095
rect 86 18075 344 18095
rect 30 18029 86 18035
rect 30 17841 60 18029
rect 115 18020 315 18045
rect 396 18035 400 18095
rect 344 18029 400 18035
rect 115 18000 185 18020
rect 90 17960 185 18000
rect 245 18000 315 18020
rect 245 17960 340 18000
rect 90 17910 340 17960
rect 90 17870 185 17910
rect 115 17850 185 17870
rect 245 17870 340 17910
rect 245 17850 315 17870
rect 30 17835 86 17841
rect 30 17775 34 17835
rect 115 17825 315 17850
rect 370 17841 400 18029
rect 344 17835 400 17841
rect 86 17775 344 17795
rect 396 17775 400 17835
rect 30 17765 400 17775
rect 430 18095 800 18105
rect 430 18035 434 18095
rect 486 18075 744 18095
rect 430 18029 486 18035
rect 430 17841 460 18029
rect 515 18020 715 18045
rect 796 18035 800 18095
rect 744 18029 800 18035
rect 515 18000 585 18020
rect 490 17960 585 18000
rect 645 18000 715 18020
rect 645 17960 740 18000
rect 490 17910 740 17960
rect 490 17870 585 17910
rect 515 17850 585 17870
rect 645 17870 740 17910
rect 645 17850 715 17870
rect 430 17835 486 17841
rect 430 17775 434 17835
rect 515 17825 715 17850
rect 770 17841 800 18029
rect 744 17835 800 17841
rect 486 17775 744 17795
rect 796 17775 800 17835
rect 430 17765 800 17775
rect 830 18095 1200 18105
rect 830 18035 834 18095
rect 886 18075 1144 18095
rect 830 18029 886 18035
rect 830 17841 860 18029
rect 915 18020 1115 18045
rect 1196 18035 1200 18095
rect 1144 18029 1200 18035
rect 915 18000 985 18020
rect 890 17960 985 18000
rect 1045 18000 1115 18020
rect 1045 17960 1140 18000
rect 890 17910 1140 17960
rect 890 17870 985 17910
rect 915 17850 985 17870
rect 1045 17870 1140 17910
rect 1045 17850 1115 17870
rect 830 17835 886 17841
rect 830 17775 834 17835
rect 915 17825 1115 17850
rect 1170 17841 1200 18029
rect 1144 17835 1200 17841
rect 886 17775 1144 17795
rect 1196 17775 1200 17835
rect 830 17765 1200 17775
rect 1230 18095 1600 18105
rect 1230 18035 1234 18095
rect 1286 18075 1544 18095
rect 1230 18029 1286 18035
rect 1230 17841 1260 18029
rect 1315 18020 1515 18045
rect 1596 18035 1600 18095
rect 1544 18029 1600 18035
rect 1315 18000 1385 18020
rect 1290 17960 1385 18000
rect 1445 18000 1515 18020
rect 1445 17960 1540 18000
rect 1290 17910 1540 17960
rect 1290 17870 1385 17910
rect 1315 17850 1385 17870
rect 1445 17870 1540 17910
rect 1445 17850 1515 17870
rect 1230 17835 1286 17841
rect 1230 17775 1234 17835
rect 1315 17825 1515 17850
rect 1570 17841 1600 18029
rect 1544 17835 1600 17841
rect 1286 17775 1544 17795
rect 1596 17775 1600 17835
rect 1230 17765 1600 17775
rect 1630 18095 2000 18105
rect 1630 18035 1634 18095
rect 1686 18075 1944 18095
rect 1630 18029 1686 18035
rect 1630 17841 1660 18029
rect 1715 18020 1915 18045
rect 1996 18035 2000 18095
rect 1944 18029 2000 18035
rect 1715 18000 1785 18020
rect 1690 17960 1785 18000
rect 1845 18000 1915 18020
rect 1845 17960 1940 18000
rect 1690 17910 1940 17960
rect 1690 17870 1785 17910
rect 1715 17850 1785 17870
rect 1845 17870 1940 17910
rect 1845 17850 1915 17870
rect 1630 17835 1686 17841
rect 1630 17775 1634 17835
rect 1715 17825 1915 17850
rect 1970 17841 2000 18029
rect 1944 17835 2000 17841
rect 1686 17775 1944 17795
rect 1996 17775 2000 17835
rect 1630 17765 2000 17775
rect 2030 18095 2400 18105
rect 2030 18035 2034 18095
rect 2086 18075 2344 18095
rect 2030 18029 2086 18035
rect 2030 17841 2060 18029
rect 2115 18020 2315 18045
rect 2396 18035 2400 18095
rect 2344 18029 2400 18035
rect 2115 18000 2185 18020
rect 2090 17960 2185 18000
rect 2245 18000 2315 18020
rect 2245 17960 2340 18000
rect 2090 17910 2340 17960
rect 2090 17870 2185 17910
rect 2115 17850 2185 17870
rect 2245 17870 2340 17910
rect 2245 17850 2315 17870
rect 2030 17835 2086 17841
rect 2030 17775 2034 17835
rect 2115 17825 2315 17850
rect 2370 17841 2400 18029
rect 2344 17835 2400 17841
rect 2086 17775 2344 17795
rect 2396 17775 2400 17835
rect 2030 17765 2400 17775
rect 2430 18095 2800 18105
rect 2430 18035 2434 18095
rect 2486 18075 2744 18095
rect 2430 18029 2486 18035
rect 2430 17841 2460 18029
rect 2515 18020 2715 18045
rect 2796 18035 2800 18095
rect 2744 18029 2800 18035
rect 2515 18000 2585 18020
rect 2490 17960 2585 18000
rect 2645 18000 2715 18020
rect 2645 17960 2740 18000
rect 2490 17910 2740 17960
rect 2490 17870 2585 17910
rect 2515 17850 2585 17870
rect 2645 17870 2740 17910
rect 2645 17850 2715 17870
rect 2430 17835 2486 17841
rect 2430 17775 2434 17835
rect 2515 17825 2715 17850
rect 2770 17841 2800 18029
rect 2744 17835 2800 17841
rect 2486 17775 2744 17795
rect 2796 17775 2800 17835
rect 2430 17765 2800 17775
rect 2830 18095 3200 18105
rect 2830 18035 2834 18095
rect 2886 18075 3144 18095
rect 2830 18029 2886 18035
rect 2830 17841 2860 18029
rect 2915 18020 3115 18045
rect 3196 18035 3200 18095
rect 3144 18029 3200 18035
rect 2915 18000 2985 18020
rect 2890 17960 2985 18000
rect 3045 18000 3115 18020
rect 3045 17960 3140 18000
rect 2890 17910 3140 17960
rect 2890 17870 2985 17910
rect 2915 17850 2985 17870
rect 3045 17870 3140 17910
rect 3045 17850 3115 17870
rect 2830 17835 2886 17841
rect 2830 17775 2834 17835
rect 2915 17825 3115 17850
rect 3170 17841 3200 18029
rect 3144 17835 3200 17841
rect 2886 17775 3144 17795
rect 3196 17775 3200 17835
rect 2830 17765 3200 17775
rect 3230 18095 3600 18105
rect 3230 18035 3234 18095
rect 3286 18075 3544 18095
rect 3230 18029 3286 18035
rect 3230 17841 3260 18029
rect 3315 18020 3515 18045
rect 3596 18035 3600 18095
rect 3544 18029 3600 18035
rect 3315 18000 3385 18020
rect 3290 17960 3385 18000
rect 3445 18000 3515 18020
rect 3445 17960 3540 18000
rect 3290 17910 3540 17960
rect 3290 17870 3385 17910
rect 3315 17850 3385 17870
rect 3445 17870 3540 17910
rect 3445 17850 3515 17870
rect 3230 17835 3286 17841
rect 3230 17775 3234 17835
rect 3315 17825 3515 17850
rect 3570 17841 3600 18029
rect 3544 17835 3600 17841
rect 3286 17775 3544 17795
rect 3596 17775 3600 17835
rect 3230 17765 3600 17775
rect 3630 18095 4000 18105
rect 3630 18035 3634 18095
rect 3686 18075 3944 18095
rect 3630 18029 3686 18035
rect 3630 17841 3660 18029
rect 3715 18020 3915 18045
rect 3996 18035 4000 18095
rect 3944 18029 4000 18035
rect 3715 18000 3785 18020
rect 3690 17960 3785 18000
rect 3845 18000 3915 18020
rect 3845 17960 3940 18000
rect 3690 17910 3940 17960
rect 3690 17870 3785 17910
rect 3715 17850 3785 17870
rect 3845 17870 3940 17910
rect 3845 17850 3915 17870
rect 3630 17835 3686 17841
rect 3630 17775 3634 17835
rect 3715 17825 3915 17850
rect 3970 17841 4000 18029
rect 3944 17835 4000 17841
rect 3686 17775 3944 17795
rect 3996 17775 4000 17835
rect 3630 17765 4000 17775
rect 4030 18095 4400 18105
rect 4030 18035 4034 18095
rect 4086 18075 4344 18095
rect 4030 18029 4086 18035
rect 4030 17841 4060 18029
rect 4115 18020 4315 18045
rect 4396 18035 4400 18095
rect 4344 18029 4400 18035
rect 4115 18000 4185 18020
rect 4090 17960 4185 18000
rect 4245 18000 4315 18020
rect 4245 17960 4340 18000
rect 4090 17910 4340 17960
rect 4090 17870 4185 17910
rect 4115 17850 4185 17870
rect 4245 17870 4340 17910
rect 4245 17850 4315 17870
rect 4030 17835 4086 17841
rect 4030 17775 4034 17835
rect 4115 17825 4315 17850
rect 4370 17841 4400 18029
rect 4344 17835 4400 17841
rect 4086 17775 4344 17795
rect 4396 17775 4400 17835
rect 4030 17765 4400 17775
rect 4430 18095 4800 18105
rect 4430 18035 4434 18095
rect 4486 18075 4744 18095
rect 4430 18029 4486 18035
rect 4430 17841 4460 18029
rect 4515 18020 4715 18045
rect 4796 18035 4800 18095
rect 4744 18029 4800 18035
rect 4515 18000 4585 18020
rect 4490 17960 4585 18000
rect 4645 18000 4715 18020
rect 4645 17960 4740 18000
rect 4490 17910 4740 17960
rect 4490 17870 4585 17910
rect 4515 17850 4585 17870
rect 4645 17870 4740 17910
rect 4645 17850 4715 17870
rect 4430 17835 4486 17841
rect 4430 17775 4434 17835
rect 4515 17825 4715 17850
rect 4770 17841 4800 18029
rect 4744 17835 4800 17841
rect 4486 17775 4744 17795
rect 4796 17775 4800 17835
rect 4430 17765 4800 17775
rect 4830 18095 5200 18105
rect 4830 18035 4834 18095
rect 4886 18075 5144 18095
rect 4830 18029 4886 18035
rect 4830 17841 4860 18029
rect 4915 18020 5115 18045
rect 5196 18035 5200 18095
rect 5144 18029 5200 18035
rect 4915 18000 4985 18020
rect 4890 17960 4985 18000
rect 5045 18000 5115 18020
rect 5045 17960 5140 18000
rect 4890 17910 5140 17960
rect 4890 17870 4985 17910
rect 4915 17850 4985 17870
rect 5045 17870 5140 17910
rect 5045 17850 5115 17870
rect 4830 17835 4886 17841
rect 4830 17775 4834 17835
rect 4915 17825 5115 17850
rect 5170 17841 5200 18029
rect 5144 17835 5200 17841
rect 4886 17775 5144 17795
rect 5196 17775 5200 17835
rect 4830 17765 5200 17775
rect 5230 18095 5600 18105
rect 5230 18035 5234 18095
rect 5286 18075 5544 18095
rect 5230 18029 5286 18035
rect 5230 17841 5260 18029
rect 5315 18020 5515 18045
rect 5596 18035 5600 18095
rect 5544 18029 5600 18035
rect 5315 18000 5385 18020
rect 5290 17960 5385 18000
rect 5445 18000 5515 18020
rect 5445 17960 5540 18000
rect 5290 17910 5540 17960
rect 5290 17870 5385 17910
rect 5315 17850 5385 17870
rect 5445 17870 5540 17910
rect 5445 17850 5515 17870
rect 5230 17835 5286 17841
rect 5230 17775 5234 17835
rect 5315 17825 5515 17850
rect 5570 17841 5600 18029
rect 5544 17835 5600 17841
rect 5286 17775 5544 17795
rect 5596 17775 5600 17835
rect 5230 17765 5600 17775
rect 5630 18095 6000 18105
rect 5630 18035 5634 18095
rect 5686 18075 5944 18095
rect 5630 18029 5686 18035
rect 5630 17841 5660 18029
rect 5715 18020 5915 18045
rect 5996 18035 6000 18095
rect 5944 18029 6000 18035
rect 5715 18000 5785 18020
rect 5690 17960 5785 18000
rect 5845 18000 5915 18020
rect 5845 17960 5940 18000
rect 5690 17910 5940 17960
rect 5690 17870 5785 17910
rect 5715 17850 5785 17870
rect 5845 17870 5940 17910
rect 5845 17850 5915 17870
rect 5630 17835 5686 17841
rect 5630 17775 5634 17835
rect 5715 17825 5915 17850
rect 5970 17841 6000 18029
rect 5944 17835 6000 17841
rect 5686 17775 5944 17795
rect 5996 17775 6000 17835
rect 5630 17765 6000 17775
rect 6030 18095 6400 18105
rect 6030 18035 6034 18095
rect 6086 18075 6344 18095
rect 6030 18029 6086 18035
rect 6030 17841 6060 18029
rect 6115 18020 6315 18045
rect 6396 18035 6400 18095
rect 6344 18029 6400 18035
rect 6115 18000 6185 18020
rect 6090 17960 6185 18000
rect 6245 18000 6315 18020
rect 6245 17960 6340 18000
rect 6090 17910 6340 17960
rect 6090 17870 6185 17910
rect 6115 17850 6185 17870
rect 6245 17870 6340 17910
rect 6245 17850 6315 17870
rect 6030 17835 6086 17841
rect 6030 17775 6034 17835
rect 6115 17825 6315 17850
rect 6370 17841 6400 18029
rect 6344 17835 6400 17841
rect 6086 17775 6344 17795
rect 6396 17775 6400 17835
rect 6030 17765 6400 17775
rect 6430 18095 6800 18105
rect 6430 18035 6434 18095
rect 6486 18075 6744 18095
rect 6430 18029 6486 18035
rect 6430 17841 6460 18029
rect 6515 18020 6715 18045
rect 6796 18035 6800 18095
rect 6744 18029 6800 18035
rect 6515 18000 6585 18020
rect 6490 17960 6585 18000
rect 6645 18000 6715 18020
rect 6645 17960 6740 18000
rect 6490 17910 6740 17960
rect 6490 17870 6585 17910
rect 6515 17850 6585 17870
rect 6645 17870 6740 17910
rect 6645 17850 6715 17870
rect 6430 17835 6486 17841
rect 6430 17775 6434 17835
rect 6515 17825 6715 17850
rect 6770 17841 6800 18029
rect 6744 17835 6800 17841
rect 6486 17775 6744 17795
rect 6796 17775 6800 17835
rect 6430 17765 6800 17775
rect 6830 18095 7200 18105
rect 6830 18035 6834 18095
rect 6886 18075 7144 18095
rect 6830 18029 6886 18035
rect 6830 17841 6860 18029
rect 6915 18020 7115 18045
rect 7196 18035 7200 18095
rect 7144 18029 7200 18035
rect 6915 18000 6985 18020
rect 6890 17960 6985 18000
rect 7045 18000 7115 18020
rect 7045 17960 7140 18000
rect 6890 17910 7140 17960
rect 6890 17870 6985 17910
rect 6915 17850 6985 17870
rect 7045 17870 7140 17910
rect 7045 17850 7115 17870
rect 6830 17835 6886 17841
rect 6830 17775 6834 17835
rect 6915 17825 7115 17850
rect 7170 17841 7200 18029
rect 7144 17835 7200 17841
rect 6886 17775 7144 17795
rect 7196 17775 7200 17835
rect 6830 17765 7200 17775
rect 7230 18095 7600 18105
rect 7230 18035 7234 18095
rect 7286 18075 7544 18095
rect 7230 18029 7286 18035
rect 7230 17841 7260 18029
rect 7315 18020 7515 18045
rect 7596 18035 7600 18095
rect 7544 18029 7600 18035
rect 7315 18000 7385 18020
rect 7290 17960 7385 18000
rect 7445 18000 7515 18020
rect 7445 17960 7540 18000
rect 7290 17910 7540 17960
rect 7290 17870 7385 17910
rect 7315 17850 7385 17870
rect 7445 17870 7540 17910
rect 7445 17850 7515 17870
rect 7230 17835 7286 17841
rect 7230 17775 7234 17835
rect 7315 17825 7515 17850
rect 7570 17841 7600 18029
rect 7544 17835 7600 17841
rect 7286 17775 7544 17795
rect 7596 17775 7600 17835
rect 7230 17765 7600 17775
rect 7630 18095 8000 18105
rect 7630 18035 7634 18095
rect 7686 18075 7944 18095
rect 7630 18029 7686 18035
rect 7630 17841 7660 18029
rect 7715 18020 7915 18045
rect 7996 18035 8000 18095
rect 7944 18029 8000 18035
rect 7715 18000 7785 18020
rect 7690 17960 7785 18000
rect 7845 18000 7915 18020
rect 7845 17960 7940 18000
rect 7690 17910 7940 17960
rect 7690 17870 7785 17910
rect 7715 17850 7785 17870
rect 7845 17870 7940 17910
rect 7845 17850 7915 17870
rect 7630 17835 7686 17841
rect 7630 17775 7634 17835
rect 7715 17825 7915 17850
rect 7970 17841 8000 18029
rect 7944 17835 8000 17841
rect 7686 17775 7944 17795
rect 7996 17775 8000 17835
rect 7630 17765 8000 17775
rect 8030 18095 8400 18105
rect 8030 18035 8034 18095
rect 8086 18075 8344 18095
rect 8030 18029 8086 18035
rect 8030 17841 8060 18029
rect 8115 18020 8315 18045
rect 8396 18035 8400 18095
rect 8344 18029 8400 18035
rect 8115 18000 8185 18020
rect 8090 17960 8185 18000
rect 8245 18000 8315 18020
rect 8245 17960 8340 18000
rect 8090 17910 8340 17960
rect 8090 17870 8185 17910
rect 8115 17850 8185 17870
rect 8245 17870 8340 17910
rect 8245 17850 8315 17870
rect 8030 17835 8086 17841
rect 8030 17775 8034 17835
rect 8115 17825 8315 17850
rect 8370 17841 8400 18029
rect 8344 17835 8400 17841
rect 8086 17775 8344 17795
rect 8396 17775 8400 17835
rect 8030 17765 8400 17775
rect 8430 18095 8800 18105
rect 8430 18035 8434 18095
rect 8486 18075 8744 18095
rect 8430 18029 8486 18035
rect 8430 17841 8460 18029
rect 8515 18020 8715 18045
rect 8796 18035 8800 18095
rect 8744 18029 8800 18035
rect 8515 18000 8585 18020
rect 8490 17960 8585 18000
rect 8645 18000 8715 18020
rect 8645 17960 8740 18000
rect 8490 17910 8740 17960
rect 8490 17870 8585 17910
rect 8515 17850 8585 17870
rect 8645 17870 8740 17910
rect 8645 17850 8715 17870
rect 8430 17835 8486 17841
rect 8430 17775 8434 17835
rect 8515 17825 8715 17850
rect 8770 17841 8800 18029
rect 8744 17835 8800 17841
rect 8486 17775 8744 17795
rect 8796 17775 8800 17835
rect 8430 17765 8800 17775
rect 8830 18095 9200 18105
rect 8830 18035 8834 18095
rect 8886 18075 9144 18095
rect 8830 18029 8886 18035
rect 8830 17841 8860 18029
rect 8915 18020 9115 18045
rect 9196 18035 9200 18095
rect 9144 18029 9200 18035
rect 8915 18000 8985 18020
rect 8890 17960 8985 18000
rect 9045 18000 9115 18020
rect 9045 17960 9140 18000
rect 8890 17910 9140 17960
rect 8890 17870 8985 17910
rect 8915 17850 8985 17870
rect 9045 17870 9140 17910
rect 9045 17850 9115 17870
rect 8830 17835 8886 17841
rect 8830 17775 8834 17835
rect 8915 17825 9115 17850
rect 9170 17841 9200 18029
rect 9144 17835 9200 17841
rect 8886 17775 9144 17795
rect 9196 17775 9200 17835
rect 8830 17765 9200 17775
rect 9230 18095 9600 18105
rect 9230 18035 9234 18095
rect 9286 18075 9544 18095
rect 9230 18029 9286 18035
rect 9230 17841 9260 18029
rect 9315 18020 9515 18045
rect 9596 18035 9600 18095
rect 9544 18029 9600 18035
rect 9315 18000 9385 18020
rect 9290 17960 9385 18000
rect 9445 18000 9515 18020
rect 9445 17960 9540 18000
rect 9290 17910 9540 17960
rect 9290 17870 9385 17910
rect 9315 17850 9385 17870
rect 9445 17870 9540 17910
rect 9445 17850 9515 17870
rect 9230 17835 9286 17841
rect 9230 17775 9234 17835
rect 9315 17825 9515 17850
rect 9570 17841 9600 18029
rect 9544 17835 9600 17841
rect 9286 17775 9544 17795
rect 9596 17775 9600 17835
rect 9230 17765 9600 17775
rect 9630 18095 10000 18105
rect 9630 18035 9634 18095
rect 9686 18075 9944 18095
rect 9630 18029 9686 18035
rect 9630 17841 9660 18029
rect 9715 18020 9915 18045
rect 9996 18035 10000 18095
rect 9944 18029 10000 18035
rect 9715 18000 9785 18020
rect 9690 17960 9785 18000
rect 9845 18000 9915 18020
rect 9845 17960 9940 18000
rect 9690 17910 9940 17960
rect 9690 17870 9785 17910
rect 9715 17850 9785 17870
rect 9845 17870 9940 17910
rect 9845 17850 9915 17870
rect 9630 17835 9686 17841
rect 9630 17775 9634 17835
rect 9715 17825 9915 17850
rect 9970 17841 10000 18029
rect 9944 17835 10000 17841
rect 9686 17775 9944 17795
rect 9996 17775 10000 17835
rect 9630 17765 10000 17775
rect 10030 18095 10400 18105
rect 10030 18035 10034 18095
rect 10086 18075 10344 18095
rect 10030 18029 10086 18035
rect 10030 17841 10060 18029
rect 10115 18020 10315 18045
rect 10396 18035 10400 18095
rect 10344 18029 10400 18035
rect 10115 18000 10185 18020
rect 10090 17960 10185 18000
rect 10245 18000 10315 18020
rect 10245 17960 10340 18000
rect 10090 17910 10340 17960
rect 10090 17870 10185 17910
rect 10115 17850 10185 17870
rect 10245 17870 10340 17910
rect 10245 17850 10315 17870
rect 10030 17835 10086 17841
rect 10030 17775 10034 17835
rect 10115 17825 10315 17850
rect 10370 17841 10400 18029
rect 10344 17835 10400 17841
rect 10086 17775 10344 17795
rect 10396 17775 10400 17835
rect 10030 17765 10400 17775
rect 10430 18095 10800 18105
rect 10430 18035 10434 18095
rect 10486 18075 10744 18095
rect 10430 18029 10486 18035
rect 10430 17841 10460 18029
rect 10515 18020 10715 18045
rect 10796 18035 10800 18095
rect 10744 18029 10800 18035
rect 10515 18000 10585 18020
rect 10490 17960 10585 18000
rect 10645 18000 10715 18020
rect 10645 17960 10740 18000
rect 10490 17910 10740 17960
rect 10490 17870 10585 17910
rect 10515 17850 10585 17870
rect 10645 17870 10740 17910
rect 10645 17850 10715 17870
rect 10430 17835 10486 17841
rect 10430 17775 10434 17835
rect 10515 17825 10715 17850
rect 10770 17841 10800 18029
rect 10744 17835 10800 17841
rect 10486 17775 10744 17795
rect 10796 17775 10800 17835
rect 10430 17765 10800 17775
rect 10830 18095 11200 18105
rect 10830 18035 10834 18095
rect 10886 18075 11144 18095
rect 10830 18029 10886 18035
rect 10830 17841 10860 18029
rect 10915 18020 11115 18045
rect 11196 18035 11200 18095
rect 11144 18029 11200 18035
rect 10915 18000 10985 18020
rect 10890 17960 10985 18000
rect 11045 18000 11115 18020
rect 11045 17960 11140 18000
rect 10890 17910 11140 17960
rect 10890 17870 10985 17910
rect 10915 17850 10985 17870
rect 11045 17870 11140 17910
rect 11045 17850 11115 17870
rect 10830 17835 10886 17841
rect 10830 17775 10834 17835
rect 10915 17825 11115 17850
rect 11170 17841 11200 18029
rect 11144 17835 11200 17841
rect 10886 17775 11144 17795
rect 11196 17775 11200 17835
rect 10830 17765 11200 17775
rect 11230 18095 11600 18105
rect 11230 18035 11234 18095
rect 11286 18075 11544 18095
rect 11230 18029 11286 18035
rect 11230 17841 11260 18029
rect 11315 18020 11515 18045
rect 11596 18035 11600 18095
rect 11544 18029 11600 18035
rect 11315 18000 11385 18020
rect 11290 17960 11385 18000
rect 11445 18000 11515 18020
rect 11445 17960 11540 18000
rect 11290 17910 11540 17960
rect 11290 17870 11385 17910
rect 11315 17850 11385 17870
rect 11445 17870 11540 17910
rect 11445 17850 11515 17870
rect 11230 17835 11286 17841
rect 11230 17775 11234 17835
rect 11315 17825 11515 17850
rect 11570 17841 11600 18029
rect 11544 17835 11600 17841
rect 11286 17775 11544 17795
rect 11596 17775 11600 17835
rect 11230 17765 11600 17775
rect 11630 18095 12000 18105
rect 11630 18035 11634 18095
rect 11686 18075 11944 18095
rect 11630 18029 11686 18035
rect 11630 17841 11660 18029
rect 11715 18020 11915 18045
rect 11996 18035 12000 18095
rect 11944 18029 12000 18035
rect 11715 18000 11785 18020
rect 11690 17960 11785 18000
rect 11845 18000 11915 18020
rect 11845 17960 11940 18000
rect 11690 17910 11940 17960
rect 11690 17870 11785 17910
rect 11715 17850 11785 17870
rect 11845 17870 11940 17910
rect 11845 17850 11915 17870
rect 11630 17835 11686 17841
rect 11630 17775 11634 17835
rect 11715 17825 11915 17850
rect 11970 17841 12000 18029
rect 11944 17835 12000 17841
rect 11686 17775 11944 17795
rect 11996 17775 12000 17835
rect 11630 17765 12000 17775
rect 12030 18095 12400 18105
rect 12030 18035 12034 18095
rect 12086 18075 12344 18095
rect 12030 18029 12086 18035
rect 12030 17841 12060 18029
rect 12115 18020 12315 18045
rect 12396 18035 12400 18095
rect 12344 18029 12400 18035
rect 12115 18000 12185 18020
rect 12090 17960 12185 18000
rect 12245 18000 12315 18020
rect 12245 17960 12340 18000
rect 12090 17910 12340 17960
rect 12090 17870 12185 17910
rect 12115 17850 12185 17870
rect 12245 17870 12340 17910
rect 12245 17850 12315 17870
rect 12030 17835 12086 17841
rect 12030 17775 12034 17835
rect 12115 17825 12315 17850
rect 12370 17841 12400 18029
rect 12344 17835 12400 17841
rect 12086 17775 12344 17795
rect 12396 17775 12400 17835
rect 12030 17765 12400 17775
rect 12430 18095 12800 18105
rect 12430 18035 12434 18095
rect 12486 18075 12744 18095
rect 12430 18029 12486 18035
rect 12430 17841 12460 18029
rect 12515 18020 12715 18045
rect 12796 18035 12800 18095
rect 12744 18029 12800 18035
rect 12515 18000 12585 18020
rect 12490 17960 12585 18000
rect 12645 18000 12715 18020
rect 12645 17960 12740 18000
rect 12490 17910 12740 17960
rect 12490 17870 12585 17910
rect 12515 17850 12585 17870
rect 12645 17870 12740 17910
rect 12645 17850 12715 17870
rect 12430 17835 12486 17841
rect 12430 17775 12434 17835
rect 12515 17825 12715 17850
rect 12770 17841 12800 18029
rect 12744 17835 12800 17841
rect 12486 17775 12744 17795
rect 12796 17775 12800 17835
rect 12430 17765 12800 17775
rect 12830 18095 13200 18105
rect 12830 18035 12834 18095
rect 12886 18075 13144 18095
rect 12830 18029 12886 18035
rect 12830 17841 12860 18029
rect 12915 18020 13115 18045
rect 13196 18035 13200 18095
rect 13144 18029 13200 18035
rect 12915 18000 12985 18020
rect 12890 17960 12985 18000
rect 13045 18000 13115 18020
rect 13045 17960 13140 18000
rect 12890 17910 13140 17960
rect 12890 17870 12985 17910
rect 12915 17850 12985 17870
rect 13045 17870 13140 17910
rect 13045 17850 13115 17870
rect 12830 17835 12886 17841
rect 12830 17775 12834 17835
rect 12915 17825 13115 17850
rect 13170 17841 13200 18029
rect 13144 17835 13200 17841
rect 12886 17775 13144 17795
rect 13196 17775 13200 17835
rect 12830 17765 13200 17775
rect -370 17725 0 17735
rect -370 17665 -366 17725
rect -314 17705 -56 17725
rect -370 17659 -314 17665
rect -370 17471 -340 17659
rect -285 17650 -85 17675
rect -4 17665 0 17725
rect -56 17659 0 17665
rect -285 17630 -215 17650
rect -310 17590 -215 17630
rect -155 17630 -85 17650
rect -155 17590 -60 17630
rect -310 17540 -60 17590
rect -310 17500 -215 17540
rect -285 17480 -215 17500
rect -155 17500 -60 17540
rect -155 17480 -85 17500
rect -370 17465 -314 17471
rect -370 17405 -366 17465
rect -285 17455 -85 17480
rect -30 17471 0 17659
rect -56 17465 0 17471
rect -314 17405 -56 17425
rect -4 17405 0 17465
rect -370 17395 0 17405
rect 30 17725 400 17735
rect 30 17665 34 17725
rect 86 17705 344 17725
rect 30 17659 86 17665
rect 30 17471 60 17659
rect 115 17650 315 17675
rect 396 17665 400 17725
rect 344 17659 400 17665
rect 115 17630 185 17650
rect 90 17590 185 17630
rect 245 17630 315 17650
rect 245 17590 340 17630
rect 90 17540 340 17590
rect 90 17500 185 17540
rect 115 17480 185 17500
rect 245 17500 340 17540
rect 245 17480 315 17500
rect 30 17465 86 17471
rect 30 17405 34 17465
rect 115 17455 315 17480
rect 370 17471 400 17659
rect 344 17465 400 17471
rect 86 17405 344 17425
rect 396 17405 400 17465
rect 30 17395 400 17405
rect 430 17725 800 17735
rect 430 17665 434 17725
rect 486 17705 744 17725
rect 430 17659 486 17665
rect 430 17471 460 17659
rect 515 17650 715 17675
rect 796 17665 800 17725
rect 744 17659 800 17665
rect 515 17630 585 17650
rect 490 17590 585 17630
rect 645 17630 715 17650
rect 645 17590 740 17630
rect 490 17540 740 17590
rect 490 17500 585 17540
rect 515 17480 585 17500
rect 645 17500 740 17540
rect 645 17480 715 17500
rect 430 17465 486 17471
rect 430 17405 434 17465
rect 515 17455 715 17480
rect 770 17471 800 17659
rect 744 17465 800 17471
rect 486 17405 744 17425
rect 796 17405 800 17465
rect 430 17395 800 17405
rect 830 17725 1200 17735
rect 830 17665 834 17725
rect 886 17705 1144 17725
rect 830 17659 886 17665
rect 830 17471 860 17659
rect 915 17650 1115 17675
rect 1196 17665 1200 17725
rect 1144 17659 1200 17665
rect 915 17630 985 17650
rect 890 17590 985 17630
rect 1045 17630 1115 17650
rect 1045 17590 1140 17630
rect 890 17540 1140 17590
rect 890 17500 985 17540
rect 915 17480 985 17500
rect 1045 17500 1140 17540
rect 1045 17480 1115 17500
rect 830 17465 886 17471
rect 830 17405 834 17465
rect 915 17455 1115 17480
rect 1170 17471 1200 17659
rect 1144 17465 1200 17471
rect 886 17405 1144 17425
rect 1196 17405 1200 17465
rect 830 17395 1200 17405
rect 1230 17725 1600 17735
rect 1230 17665 1234 17725
rect 1286 17705 1544 17725
rect 1230 17659 1286 17665
rect 1230 17471 1260 17659
rect 1315 17650 1515 17675
rect 1596 17665 1600 17725
rect 1544 17659 1600 17665
rect 1315 17630 1385 17650
rect 1290 17590 1385 17630
rect 1445 17630 1515 17650
rect 1445 17590 1540 17630
rect 1290 17540 1540 17590
rect 1290 17500 1385 17540
rect 1315 17480 1385 17500
rect 1445 17500 1540 17540
rect 1445 17480 1515 17500
rect 1230 17465 1286 17471
rect 1230 17405 1234 17465
rect 1315 17455 1515 17480
rect 1570 17471 1600 17659
rect 1544 17465 1600 17471
rect 1286 17405 1544 17425
rect 1596 17405 1600 17465
rect 1230 17395 1600 17405
rect 1630 17725 2000 17735
rect 1630 17665 1634 17725
rect 1686 17705 1944 17725
rect 1630 17659 1686 17665
rect 1630 17471 1660 17659
rect 1715 17650 1915 17675
rect 1996 17665 2000 17725
rect 1944 17659 2000 17665
rect 1715 17630 1785 17650
rect 1690 17590 1785 17630
rect 1845 17630 1915 17650
rect 1845 17590 1940 17630
rect 1690 17540 1940 17590
rect 1690 17500 1785 17540
rect 1715 17480 1785 17500
rect 1845 17500 1940 17540
rect 1845 17480 1915 17500
rect 1630 17465 1686 17471
rect 1630 17405 1634 17465
rect 1715 17455 1915 17480
rect 1970 17471 2000 17659
rect 1944 17465 2000 17471
rect 1686 17405 1944 17425
rect 1996 17405 2000 17465
rect 1630 17395 2000 17405
rect 2030 17725 2400 17735
rect 2030 17665 2034 17725
rect 2086 17705 2344 17725
rect 2030 17659 2086 17665
rect 2030 17471 2060 17659
rect 2115 17650 2315 17675
rect 2396 17665 2400 17725
rect 2344 17659 2400 17665
rect 2115 17630 2185 17650
rect 2090 17590 2185 17630
rect 2245 17630 2315 17650
rect 2245 17590 2340 17630
rect 2090 17540 2340 17590
rect 2090 17500 2185 17540
rect 2115 17480 2185 17500
rect 2245 17500 2340 17540
rect 2245 17480 2315 17500
rect 2030 17465 2086 17471
rect 2030 17405 2034 17465
rect 2115 17455 2315 17480
rect 2370 17471 2400 17659
rect 2344 17465 2400 17471
rect 2086 17405 2344 17425
rect 2396 17405 2400 17465
rect 2030 17395 2400 17405
rect 2430 17725 2800 17735
rect 2430 17665 2434 17725
rect 2486 17705 2744 17725
rect 2430 17659 2486 17665
rect 2430 17471 2460 17659
rect 2515 17650 2715 17675
rect 2796 17665 2800 17725
rect 2744 17659 2800 17665
rect 2515 17630 2585 17650
rect 2490 17590 2585 17630
rect 2645 17630 2715 17650
rect 2645 17590 2740 17630
rect 2490 17540 2740 17590
rect 2490 17500 2585 17540
rect 2515 17480 2585 17500
rect 2645 17500 2740 17540
rect 2645 17480 2715 17500
rect 2430 17465 2486 17471
rect 2430 17405 2434 17465
rect 2515 17455 2715 17480
rect 2770 17471 2800 17659
rect 2744 17465 2800 17471
rect 2486 17405 2744 17425
rect 2796 17405 2800 17465
rect 2430 17395 2800 17405
rect 2830 17725 3200 17735
rect 2830 17665 2834 17725
rect 2886 17705 3144 17725
rect 2830 17659 2886 17665
rect 2830 17471 2860 17659
rect 2915 17650 3115 17675
rect 3196 17665 3200 17725
rect 3144 17659 3200 17665
rect 2915 17630 2985 17650
rect 2890 17590 2985 17630
rect 3045 17630 3115 17650
rect 3045 17590 3140 17630
rect 2890 17540 3140 17590
rect 2890 17500 2985 17540
rect 2915 17480 2985 17500
rect 3045 17500 3140 17540
rect 3045 17480 3115 17500
rect 2830 17465 2886 17471
rect 2830 17405 2834 17465
rect 2915 17455 3115 17480
rect 3170 17471 3200 17659
rect 3144 17465 3200 17471
rect 2886 17405 3144 17425
rect 3196 17405 3200 17465
rect 2830 17395 3200 17405
rect 3230 17725 3600 17735
rect 3230 17665 3234 17725
rect 3286 17705 3544 17725
rect 3230 17659 3286 17665
rect 3230 17471 3260 17659
rect 3315 17650 3515 17675
rect 3596 17665 3600 17725
rect 3544 17659 3600 17665
rect 3315 17630 3385 17650
rect 3290 17590 3385 17630
rect 3445 17630 3515 17650
rect 3445 17590 3540 17630
rect 3290 17540 3540 17590
rect 3290 17500 3385 17540
rect 3315 17480 3385 17500
rect 3445 17500 3540 17540
rect 3445 17480 3515 17500
rect 3230 17465 3286 17471
rect 3230 17405 3234 17465
rect 3315 17455 3515 17480
rect 3570 17471 3600 17659
rect 3544 17465 3600 17471
rect 3286 17405 3544 17425
rect 3596 17405 3600 17465
rect 3230 17395 3600 17405
rect 3630 17725 4000 17735
rect 3630 17665 3634 17725
rect 3686 17705 3944 17725
rect 3630 17659 3686 17665
rect 3630 17471 3660 17659
rect 3715 17650 3915 17675
rect 3996 17665 4000 17725
rect 3944 17659 4000 17665
rect 3715 17630 3785 17650
rect 3690 17590 3785 17630
rect 3845 17630 3915 17650
rect 3845 17590 3940 17630
rect 3690 17540 3940 17590
rect 3690 17500 3785 17540
rect 3715 17480 3785 17500
rect 3845 17500 3940 17540
rect 3845 17480 3915 17500
rect 3630 17465 3686 17471
rect 3630 17405 3634 17465
rect 3715 17455 3915 17480
rect 3970 17471 4000 17659
rect 3944 17465 4000 17471
rect 3686 17405 3944 17425
rect 3996 17405 4000 17465
rect 3630 17395 4000 17405
rect 4030 17725 4400 17735
rect 4030 17665 4034 17725
rect 4086 17705 4344 17725
rect 4030 17659 4086 17665
rect 4030 17471 4060 17659
rect 4115 17650 4315 17675
rect 4396 17665 4400 17725
rect 4344 17659 4400 17665
rect 4115 17630 4185 17650
rect 4090 17590 4185 17630
rect 4245 17630 4315 17650
rect 4245 17590 4340 17630
rect 4090 17540 4340 17590
rect 4090 17500 4185 17540
rect 4115 17480 4185 17500
rect 4245 17500 4340 17540
rect 4245 17480 4315 17500
rect 4030 17465 4086 17471
rect 4030 17405 4034 17465
rect 4115 17455 4315 17480
rect 4370 17471 4400 17659
rect 4344 17465 4400 17471
rect 4086 17405 4344 17425
rect 4396 17405 4400 17465
rect 4030 17395 4400 17405
rect 4430 17725 4800 17735
rect 4430 17665 4434 17725
rect 4486 17705 4744 17725
rect 4430 17659 4486 17665
rect 4430 17471 4460 17659
rect 4515 17650 4715 17675
rect 4796 17665 4800 17725
rect 4744 17659 4800 17665
rect 4515 17630 4585 17650
rect 4490 17590 4585 17630
rect 4645 17630 4715 17650
rect 4645 17590 4740 17630
rect 4490 17540 4740 17590
rect 4490 17500 4585 17540
rect 4515 17480 4585 17500
rect 4645 17500 4740 17540
rect 4645 17480 4715 17500
rect 4430 17465 4486 17471
rect 4430 17405 4434 17465
rect 4515 17455 4715 17480
rect 4770 17471 4800 17659
rect 4744 17465 4800 17471
rect 4486 17405 4744 17425
rect 4796 17405 4800 17465
rect 4430 17395 4800 17405
rect 4830 17725 5200 17735
rect 4830 17665 4834 17725
rect 4886 17705 5144 17725
rect 4830 17659 4886 17665
rect 4830 17471 4860 17659
rect 4915 17650 5115 17675
rect 5196 17665 5200 17725
rect 5144 17659 5200 17665
rect 4915 17630 4985 17650
rect 4890 17590 4985 17630
rect 5045 17630 5115 17650
rect 5045 17590 5140 17630
rect 4890 17540 5140 17590
rect 4890 17500 4985 17540
rect 4915 17480 4985 17500
rect 5045 17500 5140 17540
rect 5045 17480 5115 17500
rect 4830 17465 4886 17471
rect 4830 17405 4834 17465
rect 4915 17455 5115 17480
rect 5170 17471 5200 17659
rect 5144 17465 5200 17471
rect 4886 17405 5144 17425
rect 5196 17405 5200 17465
rect 4830 17395 5200 17405
rect 5230 17725 5600 17735
rect 5230 17665 5234 17725
rect 5286 17705 5544 17725
rect 5230 17659 5286 17665
rect 5230 17471 5260 17659
rect 5315 17650 5515 17675
rect 5596 17665 5600 17725
rect 5544 17659 5600 17665
rect 5315 17630 5385 17650
rect 5290 17590 5385 17630
rect 5445 17630 5515 17650
rect 5445 17590 5540 17630
rect 5290 17540 5540 17590
rect 5290 17500 5385 17540
rect 5315 17480 5385 17500
rect 5445 17500 5540 17540
rect 5445 17480 5515 17500
rect 5230 17465 5286 17471
rect 5230 17405 5234 17465
rect 5315 17455 5515 17480
rect 5570 17471 5600 17659
rect 5544 17465 5600 17471
rect 5286 17405 5544 17425
rect 5596 17405 5600 17465
rect 5230 17395 5600 17405
rect 5630 17725 6000 17735
rect 5630 17665 5634 17725
rect 5686 17705 5944 17725
rect 5630 17659 5686 17665
rect 5630 17471 5660 17659
rect 5715 17650 5915 17675
rect 5996 17665 6000 17725
rect 5944 17659 6000 17665
rect 5715 17630 5785 17650
rect 5690 17590 5785 17630
rect 5845 17630 5915 17650
rect 5845 17590 5940 17630
rect 5690 17540 5940 17590
rect 5690 17500 5785 17540
rect 5715 17480 5785 17500
rect 5845 17500 5940 17540
rect 5845 17480 5915 17500
rect 5630 17465 5686 17471
rect 5630 17405 5634 17465
rect 5715 17455 5915 17480
rect 5970 17471 6000 17659
rect 5944 17465 6000 17471
rect 5686 17405 5944 17425
rect 5996 17405 6000 17465
rect 5630 17395 6000 17405
rect 6030 17725 6400 17735
rect 6030 17665 6034 17725
rect 6086 17705 6344 17725
rect 6030 17659 6086 17665
rect 6030 17471 6060 17659
rect 6115 17650 6315 17675
rect 6396 17665 6400 17725
rect 6344 17659 6400 17665
rect 6115 17630 6185 17650
rect 6090 17590 6185 17630
rect 6245 17630 6315 17650
rect 6245 17590 6340 17630
rect 6090 17540 6340 17590
rect 6090 17500 6185 17540
rect 6115 17480 6185 17500
rect 6245 17500 6340 17540
rect 6245 17480 6315 17500
rect 6030 17465 6086 17471
rect 6030 17405 6034 17465
rect 6115 17455 6315 17480
rect 6370 17471 6400 17659
rect 6344 17465 6400 17471
rect 6086 17405 6344 17425
rect 6396 17405 6400 17465
rect 6030 17395 6400 17405
rect 6430 17725 6800 17735
rect 6430 17665 6434 17725
rect 6486 17705 6744 17725
rect 6430 17659 6486 17665
rect 6430 17471 6460 17659
rect 6515 17650 6715 17675
rect 6796 17665 6800 17725
rect 6744 17659 6800 17665
rect 6515 17630 6585 17650
rect 6490 17590 6585 17630
rect 6645 17630 6715 17650
rect 6645 17590 6740 17630
rect 6490 17540 6740 17590
rect 6490 17500 6585 17540
rect 6515 17480 6585 17500
rect 6645 17500 6740 17540
rect 6645 17480 6715 17500
rect 6430 17465 6486 17471
rect 6430 17405 6434 17465
rect 6515 17455 6715 17480
rect 6770 17471 6800 17659
rect 6744 17465 6800 17471
rect 6486 17405 6744 17425
rect 6796 17405 6800 17465
rect 6430 17395 6800 17405
rect 6830 17725 7200 17735
rect 6830 17665 6834 17725
rect 6886 17705 7144 17725
rect 6830 17659 6886 17665
rect 6830 17471 6860 17659
rect 6915 17650 7115 17675
rect 7196 17665 7200 17725
rect 7144 17659 7200 17665
rect 6915 17630 6985 17650
rect 6890 17590 6985 17630
rect 7045 17630 7115 17650
rect 7045 17590 7140 17630
rect 6890 17540 7140 17590
rect 6890 17500 6985 17540
rect 6915 17480 6985 17500
rect 7045 17500 7140 17540
rect 7045 17480 7115 17500
rect 6830 17465 6886 17471
rect 6830 17405 6834 17465
rect 6915 17455 7115 17480
rect 7170 17471 7200 17659
rect 7144 17465 7200 17471
rect 6886 17405 7144 17425
rect 7196 17405 7200 17465
rect 6830 17395 7200 17405
rect 7230 17725 7600 17735
rect 7230 17665 7234 17725
rect 7286 17705 7544 17725
rect 7230 17659 7286 17665
rect 7230 17471 7260 17659
rect 7315 17650 7515 17675
rect 7596 17665 7600 17725
rect 7544 17659 7600 17665
rect 7315 17630 7385 17650
rect 7290 17590 7385 17630
rect 7445 17630 7515 17650
rect 7445 17590 7540 17630
rect 7290 17540 7540 17590
rect 7290 17500 7385 17540
rect 7315 17480 7385 17500
rect 7445 17500 7540 17540
rect 7445 17480 7515 17500
rect 7230 17465 7286 17471
rect 7230 17405 7234 17465
rect 7315 17455 7515 17480
rect 7570 17471 7600 17659
rect 7544 17465 7600 17471
rect 7286 17405 7544 17425
rect 7596 17405 7600 17465
rect 7230 17395 7600 17405
rect 7630 17725 8000 17735
rect 7630 17665 7634 17725
rect 7686 17705 7944 17725
rect 7630 17659 7686 17665
rect 7630 17471 7660 17659
rect 7715 17650 7915 17675
rect 7996 17665 8000 17725
rect 7944 17659 8000 17665
rect 7715 17630 7785 17650
rect 7690 17590 7785 17630
rect 7845 17630 7915 17650
rect 7845 17590 7940 17630
rect 7690 17540 7940 17590
rect 7690 17500 7785 17540
rect 7715 17480 7785 17500
rect 7845 17500 7940 17540
rect 7845 17480 7915 17500
rect 7630 17465 7686 17471
rect 7630 17405 7634 17465
rect 7715 17455 7915 17480
rect 7970 17471 8000 17659
rect 7944 17465 8000 17471
rect 7686 17405 7944 17425
rect 7996 17405 8000 17465
rect 7630 17395 8000 17405
rect 8030 17725 8400 17735
rect 8030 17665 8034 17725
rect 8086 17705 8344 17725
rect 8030 17659 8086 17665
rect 8030 17471 8060 17659
rect 8115 17650 8315 17675
rect 8396 17665 8400 17725
rect 8344 17659 8400 17665
rect 8115 17630 8185 17650
rect 8090 17590 8185 17630
rect 8245 17630 8315 17650
rect 8245 17590 8340 17630
rect 8090 17540 8340 17590
rect 8090 17500 8185 17540
rect 8115 17480 8185 17500
rect 8245 17500 8340 17540
rect 8245 17480 8315 17500
rect 8030 17465 8086 17471
rect 8030 17405 8034 17465
rect 8115 17455 8315 17480
rect 8370 17471 8400 17659
rect 8344 17465 8400 17471
rect 8086 17405 8344 17425
rect 8396 17405 8400 17465
rect 8030 17395 8400 17405
rect 8430 17725 8800 17735
rect 8430 17665 8434 17725
rect 8486 17705 8744 17725
rect 8430 17659 8486 17665
rect 8430 17471 8460 17659
rect 8515 17650 8715 17675
rect 8796 17665 8800 17725
rect 8744 17659 8800 17665
rect 8515 17630 8585 17650
rect 8490 17590 8585 17630
rect 8645 17630 8715 17650
rect 8645 17590 8740 17630
rect 8490 17540 8740 17590
rect 8490 17500 8585 17540
rect 8515 17480 8585 17500
rect 8645 17500 8740 17540
rect 8645 17480 8715 17500
rect 8430 17465 8486 17471
rect 8430 17405 8434 17465
rect 8515 17455 8715 17480
rect 8770 17471 8800 17659
rect 8744 17465 8800 17471
rect 8486 17405 8744 17425
rect 8796 17405 8800 17465
rect 8430 17395 8800 17405
rect 8830 17725 9200 17735
rect 8830 17665 8834 17725
rect 8886 17705 9144 17725
rect 8830 17659 8886 17665
rect 8830 17471 8860 17659
rect 8915 17650 9115 17675
rect 9196 17665 9200 17725
rect 9144 17659 9200 17665
rect 8915 17630 8985 17650
rect 8890 17590 8985 17630
rect 9045 17630 9115 17650
rect 9045 17590 9140 17630
rect 8890 17540 9140 17590
rect 8890 17500 8985 17540
rect 8915 17480 8985 17500
rect 9045 17500 9140 17540
rect 9045 17480 9115 17500
rect 8830 17465 8886 17471
rect 8830 17405 8834 17465
rect 8915 17455 9115 17480
rect 9170 17471 9200 17659
rect 9144 17465 9200 17471
rect 8886 17405 9144 17425
rect 9196 17405 9200 17465
rect 8830 17395 9200 17405
rect 9230 17725 9600 17735
rect 9230 17665 9234 17725
rect 9286 17705 9544 17725
rect 9230 17659 9286 17665
rect 9230 17471 9260 17659
rect 9315 17650 9515 17675
rect 9596 17665 9600 17725
rect 9544 17659 9600 17665
rect 9315 17630 9385 17650
rect 9290 17590 9385 17630
rect 9445 17630 9515 17650
rect 9445 17590 9540 17630
rect 9290 17540 9540 17590
rect 9290 17500 9385 17540
rect 9315 17480 9385 17500
rect 9445 17500 9540 17540
rect 9445 17480 9515 17500
rect 9230 17465 9286 17471
rect 9230 17405 9234 17465
rect 9315 17455 9515 17480
rect 9570 17471 9600 17659
rect 9544 17465 9600 17471
rect 9286 17405 9544 17425
rect 9596 17405 9600 17465
rect 9230 17395 9600 17405
rect 9630 17725 10000 17735
rect 9630 17665 9634 17725
rect 9686 17705 9944 17725
rect 9630 17659 9686 17665
rect 9630 17471 9660 17659
rect 9715 17650 9915 17675
rect 9996 17665 10000 17725
rect 9944 17659 10000 17665
rect 9715 17630 9785 17650
rect 9690 17590 9785 17630
rect 9845 17630 9915 17650
rect 9845 17590 9940 17630
rect 9690 17540 9940 17590
rect 9690 17500 9785 17540
rect 9715 17480 9785 17500
rect 9845 17500 9940 17540
rect 9845 17480 9915 17500
rect 9630 17465 9686 17471
rect 9630 17405 9634 17465
rect 9715 17455 9915 17480
rect 9970 17471 10000 17659
rect 9944 17465 10000 17471
rect 9686 17405 9944 17425
rect 9996 17405 10000 17465
rect 9630 17395 10000 17405
rect 10030 17725 10400 17735
rect 10030 17665 10034 17725
rect 10086 17705 10344 17725
rect 10030 17659 10086 17665
rect 10030 17471 10060 17659
rect 10115 17650 10315 17675
rect 10396 17665 10400 17725
rect 10344 17659 10400 17665
rect 10115 17630 10185 17650
rect 10090 17590 10185 17630
rect 10245 17630 10315 17650
rect 10245 17590 10340 17630
rect 10090 17540 10340 17590
rect 10090 17500 10185 17540
rect 10115 17480 10185 17500
rect 10245 17500 10340 17540
rect 10245 17480 10315 17500
rect 10030 17465 10086 17471
rect 10030 17405 10034 17465
rect 10115 17455 10315 17480
rect 10370 17471 10400 17659
rect 10344 17465 10400 17471
rect 10086 17405 10344 17425
rect 10396 17405 10400 17465
rect 10030 17395 10400 17405
rect 10430 17725 10800 17735
rect 10430 17665 10434 17725
rect 10486 17705 10744 17725
rect 10430 17659 10486 17665
rect 10430 17471 10460 17659
rect 10515 17650 10715 17675
rect 10796 17665 10800 17725
rect 10744 17659 10800 17665
rect 10515 17630 10585 17650
rect 10490 17590 10585 17630
rect 10645 17630 10715 17650
rect 10645 17590 10740 17630
rect 10490 17540 10740 17590
rect 10490 17500 10585 17540
rect 10515 17480 10585 17500
rect 10645 17500 10740 17540
rect 10645 17480 10715 17500
rect 10430 17465 10486 17471
rect 10430 17405 10434 17465
rect 10515 17455 10715 17480
rect 10770 17471 10800 17659
rect 10744 17465 10800 17471
rect 10486 17405 10744 17425
rect 10796 17405 10800 17465
rect 10430 17395 10800 17405
rect 10830 17725 11200 17735
rect 10830 17665 10834 17725
rect 10886 17705 11144 17725
rect 10830 17659 10886 17665
rect 10830 17471 10860 17659
rect 10915 17650 11115 17675
rect 11196 17665 11200 17725
rect 11144 17659 11200 17665
rect 10915 17630 10985 17650
rect 10890 17590 10985 17630
rect 11045 17630 11115 17650
rect 11045 17590 11140 17630
rect 10890 17540 11140 17590
rect 10890 17500 10985 17540
rect 10915 17480 10985 17500
rect 11045 17500 11140 17540
rect 11045 17480 11115 17500
rect 10830 17465 10886 17471
rect 10830 17405 10834 17465
rect 10915 17455 11115 17480
rect 11170 17471 11200 17659
rect 11144 17465 11200 17471
rect 10886 17405 11144 17425
rect 11196 17405 11200 17465
rect 10830 17395 11200 17405
rect 11230 17725 11600 17735
rect 11230 17665 11234 17725
rect 11286 17705 11544 17725
rect 11230 17659 11286 17665
rect 11230 17471 11260 17659
rect 11315 17650 11515 17675
rect 11596 17665 11600 17725
rect 11544 17659 11600 17665
rect 11315 17630 11385 17650
rect 11290 17590 11385 17630
rect 11445 17630 11515 17650
rect 11445 17590 11540 17630
rect 11290 17540 11540 17590
rect 11290 17500 11385 17540
rect 11315 17480 11385 17500
rect 11445 17500 11540 17540
rect 11445 17480 11515 17500
rect 11230 17465 11286 17471
rect 11230 17405 11234 17465
rect 11315 17455 11515 17480
rect 11570 17471 11600 17659
rect 11544 17465 11600 17471
rect 11286 17405 11544 17425
rect 11596 17405 11600 17465
rect 11230 17395 11600 17405
rect 11630 17725 12000 17735
rect 11630 17665 11634 17725
rect 11686 17705 11944 17725
rect 11630 17659 11686 17665
rect 11630 17471 11660 17659
rect 11715 17650 11915 17675
rect 11996 17665 12000 17725
rect 11944 17659 12000 17665
rect 11715 17630 11785 17650
rect 11690 17590 11785 17630
rect 11845 17630 11915 17650
rect 11845 17590 11940 17630
rect 11690 17540 11940 17590
rect 11690 17500 11785 17540
rect 11715 17480 11785 17500
rect 11845 17500 11940 17540
rect 11845 17480 11915 17500
rect 11630 17465 11686 17471
rect 11630 17405 11634 17465
rect 11715 17455 11915 17480
rect 11970 17471 12000 17659
rect 11944 17465 12000 17471
rect 11686 17405 11944 17425
rect 11996 17405 12000 17465
rect 11630 17395 12000 17405
rect 12030 17725 12400 17735
rect 12030 17665 12034 17725
rect 12086 17705 12344 17725
rect 12030 17659 12086 17665
rect 12030 17471 12060 17659
rect 12115 17650 12315 17675
rect 12396 17665 12400 17725
rect 12344 17659 12400 17665
rect 12115 17630 12185 17650
rect 12090 17590 12185 17630
rect 12245 17630 12315 17650
rect 12245 17590 12340 17630
rect 12090 17540 12340 17590
rect 12090 17500 12185 17540
rect 12115 17480 12185 17500
rect 12245 17500 12340 17540
rect 12245 17480 12315 17500
rect 12030 17465 12086 17471
rect 12030 17405 12034 17465
rect 12115 17455 12315 17480
rect 12370 17471 12400 17659
rect 12344 17465 12400 17471
rect 12086 17405 12344 17425
rect 12396 17405 12400 17465
rect 12030 17395 12400 17405
rect 12430 17725 12800 17735
rect 12430 17665 12434 17725
rect 12486 17705 12744 17725
rect 12430 17659 12486 17665
rect 12430 17471 12460 17659
rect 12515 17650 12715 17675
rect 12796 17665 12800 17725
rect 12744 17659 12800 17665
rect 12515 17630 12585 17650
rect 12490 17590 12585 17630
rect 12645 17630 12715 17650
rect 12645 17590 12740 17630
rect 12490 17540 12740 17590
rect 12490 17500 12585 17540
rect 12515 17480 12585 17500
rect 12645 17500 12740 17540
rect 12645 17480 12715 17500
rect 12430 17465 12486 17471
rect 12430 17405 12434 17465
rect 12515 17455 12715 17480
rect 12770 17471 12800 17659
rect 12744 17465 12800 17471
rect 12486 17405 12744 17425
rect 12796 17405 12800 17465
rect 12430 17395 12800 17405
rect 12830 17725 13200 17735
rect 12830 17665 12834 17725
rect 12886 17705 13144 17725
rect 12830 17659 12886 17665
rect 12830 17471 12860 17659
rect 12915 17650 13115 17675
rect 13196 17665 13200 17725
rect 13144 17659 13200 17665
rect 12915 17630 12985 17650
rect 12890 17590 12985 17630
rect 13045 17630 13115 17650
rect 13045 17590 13140 17630
rect 12890 17540 13140 17590
rect 12890 17500 12985 17540
rect 12915 17480 12985 17500
rect 13045 17500 13140 17540
rect 13045 17480 13115 17500
rect 12830 17465 12886 17471
rect 12830 17405 12834 17465
rect 12915 17455 13115 17480
rect 13170 17471 13200 17659
rect 13144 17465 13200 17471
rect 12886 17405 13144 17425
rect 13196 17405 13200 17465
rect 12830 17395 13200 17405
rect -370 17355 0 17365
rect -370 17295 -366 17355
rect -314 17335 -56 17355
rect -370 17289 -314 17295
rect -370 17101 -340 17289
rect -285 17280 -85 17305
rect -4 17295 0 17355
rect -56 17289 0 17295
rect -285 17260 -215 17280
rect -310 17220 -215 17260
rect -155 17260 -85 17280
rect -155 17220 -60 17260
rect -310 17170 -60 17220
rect -310 17130 -215 17170
rect -285 17110 -215 17130
rect -155 17130 -60 17170
rect -155 17110 -85 17130
rect -370 17095 -314 17101
rect -370 17035 -366 17095
rect -285 17085 -85 17110
rect -30 17101 0 17289
rect -56 17095 0 17101
rect -314 17035 -56 17055
rect -4 17035 0 17095
rect -370 17025 0 17035
rect 30 17355 400 17365
rect 30 17295 34 17355
rect 86 17335 344 17355
rect 30 17289 86 17295
rect 30 17101 60 17289
rect 115 17280 315 17305
rect 396 17295 400 17355
rect 344 17289 400 17295
rect 115 17260 185 17280
rect 90 17220 185 17260
rect 245 17260 315 17280
rect 245 17220 340 17260
rect 90 17170 340 17220
rect 90 17130 185 17170
rect 115 17110 185 17130
rect 245 17130 340 17170
rect 245 17110 315 17130
rect 30 17095 86 17101
rect 30 17035 34 17095
rect 115 17085 315 17110
rect 370 17101 400 17289
rect 344 17095 400 17101
rect 86 17035 344 17055
rect 396 17035 400 17095
rect 30 17025 400 17035
rect 430 17355 800 17365
rect 430 17295 434 17355
rect 486 17335 744 17355
rect 430 17289 486 17295
rect 430 17101 460 17289
rect 515 17280 715 17305
rect 796 17295 800 17355
rect 744 17289 800 17295
rect 515 17260 585 17280
rect 490 17220 585 17260
rect 645 17260 715 17280
rect 645 17220 740 17260
rect 490 17170 740 17220
rect 490 17130 585 17170
rect 515 17110 585 17130
rect 645 17130 740 17170
rect 645 17110 715 17130
rect 430 17095 486 17101
rect 430 17035 434 17095
rect 515 17085 715 17110
rect 770 17101 800 17289
rect 744 17095 800 17101
rect 486 17035 744 17055
rect 796 17035 800 17095
rect 430 17025 800 17035
rect 830 17355 1200 17365
rect 830 17295 834 17355
rect 886 17335 1144 17355
rect 830 17289 886 17295
rect 830 17101 860 17289
rect 915 17280 1115 17305
rect 1196 17295 1200 17355
rect 1144 17289 1200 17295
rect 915 17260 985 17280
rect 890 17220 985 17260
rect 1045 17260 1115 17280
rect 1045 17220 1140 17260
rect 890 17170 1140 17220
rect 890 17130 985 17170
rect 915 17110 985 17130
rect 1045 17130 1140 17170
rect 1045 17110 1115 17130
rect 830 17095 886 17101
rect 830 17035 834 17095
rect 915 17085 1115 17110
rect 1170 17101 1200 17289
rect 1144 17095 1200 17101
rect 886 17035 1144 17055
rect 1196 17035 1200 17095
rect 830 17025 1200 17035
rect 1230 17355 1600 17365
rect 1230 17295 1234 17355
rect 1286 17335 1544 17355
rect 1230 17289 1286 17295
rect 1230 17101 1260 17289
rect 1315 17280 1515 17305
rect 1596 17295 1600 17355
rect 1544 17289 1600 17295
rect 1315 17260 1385 17280
rect 1290 17220 1385 17260
rect 1445 17260 1515 17280
rect 1445 17220 1540 17260
rect 1290 17170 1540 17220
rect 1290 17130 1385 17170
rect 1315 17110 1385 17130
rect 1445 17130 1540 17170
rect 1445 17110 1515 17130
rect 1230 17095 1286 17101
rect 1230 17035 1234 17095
rect 1315 17085 1515 17110
rect 1570 17101 1600 17289
rect 1544 17095 1600 17101
rect 1286 17035 1544 17055
rect 1596 17035 1600 17095
rect 1230 17025 1600 17035
rect 1630 17355 2000 17365
rect 1630 17295 1634 17355
rect 1686 17335 1944 17355
rect 1630 17289 1686 17295
rect 1630 17101 1660 17289
rect 1715 17280 1915 17305
rect 1996 17295 2000 17355
rect 1944 17289 2000 17295
rect 1715 17260 1785 17280
rect 1690 17220 1785 17260
rect 1845 17260 1915 17280
rect 1845 17220 1940 17260
rect 1690 17170 1940 17220
rect 1690 17130 1785 17170
rect 1715 17110 1785 17130
rect 1845 17130 1940 17170
rect 1845 17110 1915 17130
rect 1630 17095 1686 17101
rect 1630 17035 1634 17095
rect 1715 17085 1915 17110
rect 1970 17101 2000 17289
rect 1944 17095 2000 17101
rect 1686 17035 1944 17055
rect 1996 17035 2000 17095
rect 1630 17025 2000 17035
rect 2030 17355 2400 17365
rect 2030 17295 2034 17355
rect 2086 17335 2344 17355
rect 2030 17289 2086 17295
rect 2030 17101 2060 17289
rect 2115 17280 2315 17305
rect 2396 17295 2400 17355
rect 2344 17289 2400 17295
rect 2115 17260 2185 17280
rect 2090 17220 2185 17260
rect 2245 17260 2315 17280
rect 2245 17220 2340 17260
rect 2090 17170 2340 17220
rect 2090 17130 2185 17170
rect 2115 17110 2185 17130
rect 2245 17130 2340 17170
rect 2245 17110 2315 17130
rect 2030 17095 2086 17101
rect 2030 17035 2034 17095
rect 2115 17085 2315 17110
rect 2370 17101 2400 17289
rect 2344 17095 2400 17101
rect 2086 17035 2344 17055
rect 2396 17035 2400 17095
rect 2030 17025 2400 17035
rect 2430 17355 2800 17365
rect 2430 17295 2434 17355
rect 2486 17335 2744 17355
rect 2430 17289 2486 17295
rect 2430 17101 2460 17289
rect 2515 17280 2715 17305
rect 2796 17295 2800 17355
rect 2744 17289 2800 17295
rect 2515 17260 2585 17280
rect 2490 17220 2585 17260
rect 2645 17260 2715 17280
rect 2645 17220 2740 17260
rect 2490 17170 2740 17220
rect 2490 17130 2585 17170
rect 2515 17110 2585 17130
rect 2645 17130 2740 17170
rect 2645 17110 2715 17130
rect 2430 17095 2486 17101
rect 2430 17035 2434 17095
rect 2515 17085 2715 17110
rect 2770 17101 2800 17289
rect 2744 17095 2800 17101
rect 2486 17035 2744 17055
rect 2796 17035 2800 17095
rect 2430 17025 2800 17035
rect 2830 17355 3200 17365
rect 2830 17295 2834 17355
rect 2886 17335 3144 17355
rect 2830 17289 2886 17295
rect 2830 17101 2860 17289
rect 2915 17280 3115 17305
rect 3196 17295 3200 17355
rect 3144 17289 3200 17295
rect 2915 17260 2985 17280
rect 2890 17220 2985 17260
rect 3045 17260 3115 17280
rect 3045 17220 3140 17260
rect 2890 17170 3140 17220
rect 2890 17130 2985 17170
rect 2915 17110 2985 17130
rect 3045 17130 3140 17170
rect 3045 17110 3115 17130
rect 2830 17095 2886 17101
rect 2830 17035 2834 17095
rect 2915 17085 3115 17110
rect 3170 17101 3200 17289
rect 3144 17095 3200 17101
rect 2886 17035 3144 17055
rect 3196 17035 3200 17095
rect 2830 17025 3200 17035
rect 3230 17355 3600 17365
rect 3230 17295 3234 17355
rect 3286 17335 3544 17355
rect 3230 17289 3286 17295
rect 3230 17101 3260 17289
rect 3315 17280 3515 17305
rect 3596 17295 3600 17355
rect 3544 17289 3600 17295
rect 3315 17260 3385 17280
rect 3290 17220 3385 17260
rect 3445 17260 3515 17280
rect 3445 17220 3540 17260
rect 3290 17170 3540 17220
rect 3290 17130 3385 17170
rect 3315 17110 3385 17130
rect 3445 17130 3540 17170
rect 3445 17110 3515 17130
rect 3230 17095 3286 17101
rect 3230 17035 3234 17095
rect 3315 17085 3515 17110
rect 3570 17101 3600 17289
rect 3544 17095 3600 17101
rect 3286 17035 3544 17055
rect 3596 17035 3600 17095
rect 3230 17025 3600 17035
rect 3630 17355 4000 17365
rect 3630 17295 3634 17355
rect 3686 17335 3944 17355
rect 3630 17289 3686 17295
rect 3630 17101 3660 17289
rect 3715 17280 3915 17305
rect 3996 17295 4000 17355
rect 3944 17289 4000 17295
rect 3715 17260 3785 17280
rect 3690 17220 3785 17260
rect 3845 17260 3915 17280
rect 3845 17220 3940 17260
rect 3690 17170 3940 17220
rect 3690 17130 3785 17170
rect 3715 17110 3785 17130
rect 3845 17130 3940 17170
rect 3845 17110 3915 17130
rect 3630 17095 3686 17101
rect 3630 17035 3634 17095
rect 3715 17085 3915 17110
rect 3970 17101 4000 17289
rect 3944 17095 4000 17101
rect 3686 17035 3944 17055
rect 3996 17035 4000 17095
rect 3630 17025 4000 17035
rect 4030 17355 4400 17365
rect 4030 17295 4034 17355
rect 4086 17335 4344 17355
rect 4030 17289 4086 17295
rect 4030 17101 4060 17289
rect 4115 17280 4315 17305
rect 4396 17295 4400 17355
rect 4344 17289 4400 17295
rect 4115 17260 4185 17280
rect 4090 17220 4185 17260
rect 4245 17260 4315 17280
rect 4245 17220 4340 17260
rect 4090 17170 4340 17220
rect 4090 17130 4185 17170
rect 4115 17110 4185 17130
rect 4245 17130 4340 17170
rect 4245 17110 4315 17130
rect 4030 17095 4086 17101
rect 4030 17035 4034 17095
rect 4115 17085 4315 17110
rect 4370 17101 4400 17289
rect 4344 17095 4400 17101
rect 4086 17035 4344 17055
rect 4396 17035 4400 17095
rect 4030 17025 4400 17035
rect 4430 17355 4800 17365
rect 4430 17295 4434 17355
rect 4486 17335 4744 17355
rect 4430 17289 4486 17295
rect 4430 17101 4460 17289
rect 4515 17280 4715 17305
rect 4796 17295 4800 17355
rect 4744 17289 4800 17295
rect 4515 17260 4585 17280
rect 4490 17220 4585 17260
rect 4645 17260 4715 17280
rect 4645 17220 4740 17260
rect 4490 17170 4740 17220
rect 4490 17130 4585 17170
rect 4515 17110 4585 17130
rect 4645 17130 4740 17170
rect 4645 17110 4715 17130
rect 4430 17095 4486 17101
rect 4430 17035 4434 17095
rect 4515 17085 4715 17110
rect 4770 17101 4800 17289
rect 4744 17095 4800 17101
rect 4486 17035 4744 17055
rect 4796 17035 4800 17095
rect 4430 17025 4800 17035
rect 4830 17355 5200 17365
rect 4830 17295 4834 17355
rect 4886 17335 5144 17355
rect 4830 17289 4886 17295
rect 4830 17101 4860 17289
rect 4915 17280 5115 17305
rect 5196 17295 5200 17355
rect 5144 17289 5200 17295
rect 4915 17260 4985 17280
rect 4890 17220 4985 17260
rect 5045 17260 5115 17280
rect 5045 17220 5140 17260
rect 4890 17170 5140 17220
rect 4890 17130 4985 17170
rect 4915 17110 4985 17130
rect 5045 17130 5140 17170
rect 5045 17110 5115 17130
rect 4830 17095 4886 17101
rect 4830 17035 4834 17095
rect 4915 17085 5115 17110
rect 5170 17101 5200 17289
rect 5144 17095 5200 17101
rect 4886 17035 5144 17055
rect 5196 17035 5200 17095
rect 4830 17025 5200 17035
rect 5230 17355 5600 17365
rect 5230 17295 5234 17355
rect 5286 17335 5544 17355
rect 5230 17289 5286 17295
rect 5230 17101 5260 17289
rect 5315 17280 5515 17305
rect 5596 17295 5600 17355
rect 5544 17289 5600 17295
rect 5315 17260 5385 17280
rect 5290 17220 5385 17260
rect 5445 17260 5515 17280
rect 5445 17220 5540 17260
rect 5290 17170 5540 17220
rect 5290 17130 5385 17170
rect 5315 17110 5385 17130
rect 5445 17130 5540 17170
rect 5445 17110 5515 17130
rect 5230 17095 5286 17101
rect 5230 17035 5234 17095
rect 5315 17085 5515 17110
rect 5570 17101 5600 17289
rect 5544 17095 5600 17101
rect 5286 17035 5544 17055
rect 5596 17035 5600 17095
rect 5230 17025 5600 17035
rect 5630 17355 6000 17365
rect 5630 17295 5634 17355
rect 5686 17335 5944 17355
rect 5630 17289 5686 17295
rect 5630 17101 5660 17289
rect 5715 17280 5915 17305
rect 5996 17295 6000 17355
rect 5944 17289 6000 17295
rect 5715 17260 5785 17280
rect 5690 17220 5785 17260
rect 5845 17260 5915 17280
rect 5845 17220 5940 17260
rect 5690 17170 5940 17220
rect 5690 17130 5785 17170
rect 5715 17110 5785 17130
rect 5845 17130 5940 17170
rect 5845 17110 5915 17130
rect 5630 17095 5686 17101
rect 5630 17035 5634 17095
rect 5715 17085 5915 17110
rect 5970 17101 6000 17289
rect 5944 17095 6000 17101
rect 5686 17035 5944 17055
rect 5996 17035 6000 17095
rect 5630 17025 6000 17035
rect 6030 17355 6400 17365
rect 6030 17295 6034 17355
rect 6086 17335 6344 17355
rect 6030 17289 6086 17295
rect 6030 17101 6060 17289
rect 6115 17280 6315 17305
rect 6396 17295 6400 17355
rect 6344 17289 6400 17295
rect 6115 17260 6185 17280
rect 6090 17220 6185 17260
rect 6245 17260 6315 17280
rect 6245 17220 6340 17260
rect 6090 17170 6340 17220
rect 6090 17130 6185 17170
rect 6115 17110 6185 17130
rect 6245 17130 6340 17170
rect 6245 17110 6315 17130
rect 6030 17095 6086 17101
rect 6030 17035 6034 17095
rect 6115 17085 6315 17110
rect 6370 17101 6400 17289
rect 6344 17095 6400 17101
rect 6086 17035 6344 17055
rect 6396 17035 6400 17095
rect 6030 17025 6400 17035
rect 6430 17355 6800 17365
rect 6430 17295 6434 17355
rect 6486 17335 6744 17355
rect 6430 17289 6486 17295
rect 6430 17101 6460 17289
rect 6515 17280 6715 17305
rect 6796 17295 6800 17355
rect 6744 17289 6800 17295
rect 6515 17260 6585 17280
rect 6490 17220 6585 17260
rect 6645 17260 6715 17280
rect 6645 17220 6740 17260
rect 6490 17170 6740 17220
rect 6490 17130 6585 17170
rect 6515 17110 6585 17130
rect 6645 17130 6740 17170
rect 6645 17110 6715 17130
rect 6430 17095 6486 17101
rect 6430 17035 6434 17095
rect 6515 17085 6715 17110
rect 6770 17101 6800 17289
rect 6744 17095 6800 17101
rect 6486 17035 6744 17055
rect 6796 17035 6800 17095
rect 6430 17025 6800 17035
rect 6830 17355 7200 17365
rect 6830 17295 6834 17355
rect 6886 17335 7144 17355
rect 6830 17289 6886 17295
rect 6830 17101 6860 17289
rect 6915 17280 7115 17305
rect 7196 17295 7200 17355
rect 7144 17289 7200 17295
rect 6915 17260 6985 17280
rect 6890 17220 6985 17260
rect 7045 17260 7115 17280
rect 7045 17220 7140 17260
rect 6890 17170 7140 17220
rect 6890 17130 6985 17170
rect 6915 17110 6985 17130
rect 7045 17130 7140 17170
rect 7045 17110 7115 17130
rect 6830 17095 6886 17101
rect 6830 17035 6834 17095
rect 6915 17085 7115 17110
rect 7170 17101 7200 17289
rect 7144 17095 7200 17101
rect 6886 17035 7144 17055
rect 7196 17035 7200 17095
rect 6830 17025 7200 17035
rect 7230 17355 7600 17365
rect 7230 17295 7234 17355
rect 7286 17335 7544 17355
rect 7230 17289 7286 17295
rect 7230 17101 7260 17289
rect 7315 17280 7515 17305
rect 7596 17295 7600 17355
rect 7544 17289 7600 17295
rect 7315 17260 7385 17280
rect 7290 17220 7385 17260
rect 7445 17260 7515 17280
rect 7445 17220 7540 17260
rect 7290 17170 7540 17220
rect 7290 17130 7385 17170
rect 7315 17110 7385 17130
rect 7445 17130 7540 17170
rect 7445 17110 7515 17130
rect 7230 17095 7286 17101
rect 7230 17035 7234 17095
rect 7315 17085 7515 17110
rect 7570 17101 7600 17289
rect 7544 17095 7600 17101
rect 7286 17035 7544 17055
rect 7596 17035 7600 17095
rect 7230 17025 7600 17035
rect 7630 17355 8000 17365
rect 7630 17295 7634 17355
rect 7686 17335 7944 17355
rect 7630 17289 7686 17295
rect 7630 17101 7660 17289
rect 7715 17280 7915 17305
rect 7996 17295 8000 17355
rect 7944 17289 8000 17295
rect 7715 17260 7785 17280
rect 7690 17220 7785 17260
rect 7845 17260 7915 17280
rect 7845 17220 7940 17260
rect 7690 17170 7940 17220
rect 7690 17130 7785 17170
rect 7715 17110 7785 17130
rect 7845 17130 7940 17170
rect 7845 17110 7915 17130
rect 7630 17095 7686 17101
rect 7630 17035 7634 17095
rect 7715 17085 7915 17110
rect 7970 17101 8000 17289
rect 7944 17095 8000 17101
rect 7686 17035 7944 17055
rect 7996 17035 8000 17095
rect 7630 17025 8000 17035
rect 8030 17355 8400 17365
rect 8030 17295 8034 17355
rect 8086 17335 8344 17355
rect 8030 17289 8086 17295
rect 8030 17101 8060 17289
rect 8115 17280 8315 17305
rect 8396 17295 8400 17355
rect 8344 17289 8400 17295
rect 8115 17260 8185 17280
rect 8090 17220 8185 17260
rect 8245 17260 8315 17280
rect 8245 17220 8340 17260
rect 8090 17170 8340 17220
rect 8090 17130 8185 17170
rect 8115 17110 8185 17130
rect 8245 17130 8340 17170
rect 8245 17110 8315 17130
rect 8030 17095 8086 17101
rect 8030 17035 8034 17095
rect 8115 17085 8315 17110
rect 8370 17101 8400 17289
rect 8344 17095 8400 17101
rect 8086 17035 8344 17055
rect 8396 17035 8400 17095
rect 8030 17025 8400 17035
rect 8430 17355 8800 17365
rect 8430 17295 8434 17355
rect 8486 17335 8744 17355
rect 8430 17289 8486 17295
rect 8430 17101 8460 17289
rect 8515 17280 8715 17305
rect 8796 17295 8800 17355
rect 8744 17289 8800 17295
rect 8515 17260 8585 17280
rect 8490 17220 8585 17260
rect 8645 17260 8715 17280
rect 8645 17220 8740 17260
rect 8490 17170 8740 17220
rect 8490 17130 8585 17170
rect 8515 17110 8585 17130
rect 8645 17130 8740 17170
rect 8645 17110 8715 17130
rect 8430 17095 8486 17101
rect 8430 17035 8434 17095
rect 8515 17085 8715 17110
rect 8770 17101 8800 17289
rect 8744 17095 8800 17101
rect 8486 17035 8744 17055
rect 8796 17035 8800 17095
rect 8430 17025 8800 17035
rect 8830 17355 9200 17365
rect 8830 17295 8834 17355
rect 8886 17335 9144 17355
rect 8830 17289 8886 17295
rect 8830 17101 8860 17289
rect 8915 17280 9115 17305
rect 9196 17295 9200 17355
rect 9144 17289 9200 17295
rect 8915 17260 8985 17280
rect 8890 17220 8985 17260
rect 9045 17260 9115 17280
rect 9045 17220 9140 17260
rect 8890 17170 9140 17220
rect 8890 17130 8985 17170
rect 8915 17110 8985 17130
rect 9045 17130 9140 17170
rect 9045 17110 9115 17130
rect 8830 17095 8886 17101
rect 8830 17035 8834 17095
rect 8915 17085 9115 17110
rect 9170 17101 9200 17289
rect 9144 17095 9200 17101
rect 8886 17035 9144 17055
rect 9196 17035 9200 17095
rect 8830 17025 9200 17035
rect 9230 17355 9600 17365
rect 9230 17295 9234 17355
rect 9286 17335 9544 17355
rect 9230 17289 9286 17295
rect 9230 17101 9260 17289
rect 9315 17280 9515 17305
rect 9596 17295 9600 17355
rect 9544 17289 9600 17295
rect 9315 17260 9385 17280
rect 9290 17220 9385 17260
rect 9445 17260 9515 17280
rect 9445 17220 9540 17260
rect 9290 17170 9540 17220
rect 9290 17130 9385 17170
rect 9315 17110 9385 17130
rect 9445 17130 9540 17170
rect 9445 17110 9515 17130
rect 9230 17095 9286 17101
rect 9230 17035 9234 17095
rect 9315 17085 9515 17110
rect 9570 17101 9600 17289
rect 9544 17095 9600 17101
rect 9286 17035 9544 17055
rect 9596 17035 9600 17095
rect 9230 17025 9600 17035
rect 9630 17355 10000 17365
rect 9630 17295 9634 17355
rect 9686 17335 9944 17355
rect 9630 17289 9686 17295
rect 9630 17101 9660 17289
rect 9715 17280 9915 17305
rect 9996 17295 10000 17355
rect 9944 17289 10000 17295
rect 9715 17260 9785 17280
rect 9690 17220 9785 17260
rect 9845 17260 9915 17280
rect 9845 17220 9940 17260
rect 9690 17170 9940 17220
rect 9690 17130 9785 17170
rect 9715 17110 9785 17130
rect 9845 17130 9940 17170
rect 9845 17110 9915 17130
rect 9630 17095 9686 17101
rect 9630 17035 9634 17095
rect 9715 17085 9915 17110
rect 9970 17101 10000 17289
rect 9944 17095 10000 17101
rect 9686 17035 9944 17055
rect 9996 17035 10000 17095
rect 9630 17025 10000 17035
rect 10030 17355 10400 17365
rect 10030 17295 10034 17355
rect 10086 17335 10344 17355
rect 10030 17289 10086 17295
rect 10030 17101 10060 17289
rect 10115 17280 10315 17305
rect 10396 17295 10400 17355
rect 10344 17289 10400 17295
rect 10115 17260 10185 17280
rect 10090 17220 10185 17260
rect 10245 17260 10315 17280
rect 10245 17220 10340 17260
rect 10090 17170 10340 17220
rect 10090 17130 10185 17170
rect 10115 17110 10185 17130
rect 10245 17130 10340 17170
rect 10245 17110 10315 17130
rect 10030 17095 10086 17101
rect 10030 17035 10034 17095
rect 10115 17085 10315 17110
rect 10370 17101 10400 17289
rect 10344 17095 10400 17101
rect 10086 17035 10344 17055
rect 10396 17035 10400 17095
rect 10030 17025 10400 17035
rect 10430 17355 10800 17365
rect 10430 17295 10434 17355
rect 10486 17335 10744 17355
rect 10430 17289 10486 17295
rect 10430 17101 10460 17289
rect 10515 17280 10715 17305
rect 10796 17295 10800 17355
rect 10744 17289 10800 17295
rect 10515 17260 10585 17280
rect 10490 17220 10585 17260
rect 10645 17260 10715 17280
rect 10645 17220 10740 17260
rect 10490 17170 10740 17220
rect 10490 17130 10585 17170
rect 10515 17110 10585 17130
rect 10645 17130 10740 17170
rect 10645 17110 10715 17130
rect 10430 17095 10486 17101
rect 10430 17035 10434 17095
rect 10515 17085 10715 17110
rect 10770 17101 10800 17289
rect 10744 17095 10800 17101
rect 10486 17035 10744 17055
rect 10796 17035 10800 17095
rect 10430 17025 10800 17035
rect 10830 17355 11200 17365
rect 10830 17295 10834 17355
rect 10886 17335 11144 17355
rect 10830 17289 10886 17295
rect 10830 17101 10860 17289
rect 10915 17280 11115 17305
rect 11196 17295 11200 17355
rect 11144 17289 11200 17295
rect 10915 17260 10985 17280
rect 10890 17220 10985 17260
rect 11045 17260 11115 17280
rect 11045 17220 11140 17260
rect 10890 17170 11140 17220
rect 10890 17130 10985 17170
rect 10915 17110 10985 17130
rect 11045 17130 11140 17170
rect 11045 17110 11115 17130
rect 10830 17095 10886 17101
rect 10830 17035 10834 17095
rect 10915 17085 11115 17110
rect 11170 17101 11200 17289
rect 11144 17095 11200 17101
rect 10886 17035 11144 17055
rect 11196 17035 11200 17095
rect 10830 17025 11200 17035
rect 11230 17355 11600 17365
rect 11230 17295 11234 17355
rect 11286 17335 11544 17355
rect 11230 17289 11286 17295
rect 11230 17101 11260 17289
rect 11315 17280 11515 17305
rect 11596 17295 11600 17355
rect 11544 17289 11600 17295
rect 11315 17260 11385 17280
rect 11290 17220 11385 17260
rect 11445 17260 11515 17280
rect 11445 17220 11540 17260
rect 11290 17170 11540 17220
rect 11290 17130 11385 17170
rect 11315 17110 11385 17130
rect 11445 17130 11540 17170
rect 11445 17110 11515 17130
rect 11230 17095 11286 17101
rect 11230 17035 11234 17095
rect 11315 17085 11515 17110
rect 11570 17101 11600 17289
rect 11544 17095 11600 17101
rect 11286 17035 11544 17055
rect 11596 17035 11600 17095
rect 11230 17025 11600 17035
rect 11630 17355 12000 17365
rect 11630 17295 11634 17355
rect 11686 17335 11944 17355
rect 11630 17289 11686 17295
rect 11630 17101 11660 17289
rect 11715 17280 11915 17305
rect 11996 17295 12000 17355
rect 11944 17289 12000 17295
rect 11715 17260 11785 17280
rect 11690 17220 11785 17260
rect 11845 17260 11915 17280
rect 11845 17220 11940 17260
rect 11690 17170 11940 17220
rect 11690 17130 11785 17170
rect 11715 17110 11785 17130
rect 11845 17130 11940 17170
rect 11845 17110 11915 17130
rect 11630 17095 11686 17101
rect 11630 17035 11634 17095
rect 11715 17085 11915 17110
rect 11970 17101 12000 17289
rect 11944 17095 12000 17101
rect 11686 17035 11944 17055
rect 11996 17035 12000 17095
rect 11630 17025 12000 17035
rect 12030 17355 12400 17365
rect 12030 17295 12034 17355
rect 12086 17335 12344 17355
rect 12030 17289 12086 17295
rect 12030 17101 12060 17289
rect 12115 17280 12315 17305
rect 12396 17295 12400 17355
rect 12344 17289 12400 17295
rect 12115 17260 12185 17280
rect 12090 17220 12185 17260
rect 12245 17260 12315 17280
rect 12245 17220 12340 17260
rect 12090 17170 12340 17220
rect 12090 17130 12185 17170
rect 12115 17110 12185 17130
rect 12245 17130 12340 17170
rect 12245 17110 12315 17130
rect 12030 17095 12086 17101
rect 12030 17035 12034 17095
rect 12115 17085 12315 17110
rect 12370 17101 12400 17289
rect 12344 17095 12400 17101
rect 12086 17035 12344 17055
rect 12396 17035 12400 17095
rect 12030 17025 12400 17035
rect 12430 17355 12800 17365
rect 12430 17295 12434 17355
rect 12486 17335 12744 17355
rect 12430 17289 12486 17295
rect 12430 17101 12460 17289
rect 12515 17280 12715 17305
rect 12796 17295 12800 17355
rect 12744 17289 12800 17295
rect 12515 17260 12585 17280
rect 12490 17220 12585 17260
rect 12645 17260 12715 17280
rect 12645 17220 12740 17260
rect 12490 17170 12740 17220
rect 12490 17130 12585 17170
rect 12515 17110 12585 17130
rect 12645 17130 12740 17170
rect 12645 17110 12715 17130
rect 12430 17095 12486 17101
rect 12430 17035 12434 17095
rect 12515 17085 12715 17110
rect 12770 17101 12800 17289
rect 12744 17095 12800 17101
rect 12486 17035 12744 17055
rect 12796 17035 12800 17095
rect 12430 17025 12800 17035
rect 12830 17355 13200 17365
rect 12830 17295 12834 17355
rect 12886 17335 13144 17355
rect 12830 17289 12886 17295
rect 12830 17101 12860 17289
rect 12915 17280 13115 17305
rect 13196 17295 13200 17355
rect 13144 17289 13200 17295
rect 12915 17260 12985 17280
rect 12890 17220 12985 17260
rect 13045 17260 13115 17280
rect 13045 17220 13140 17260
rect 12890 17170 13140 17220
rect 12890 17130 12985 17170
rect 12915 17110 12985 17130
rect 13045 17130 13140 17170
rect 13045 17110 13115 17130
rect 12830 17095 12886 17101
rect 12830 17035 12834 17095
rect 12915 17085 13115 17110
rect 13170 17101 13200 17289
rect 13144 17095 13200 17101
rect 12886 17035 13144 17055
rect 13196 17035 13200 17095
rect 12830 17025 13200 17035
rect -370 16985 0 16995
rect -370 16925 -366 16985
rect -314 16965 -56 16985
rect -370 16919 -314 16925
rect -370 16731 -340 16919
rect -285 16910 -85 16935
rect -4 16925 0 16985
rect -56 16919 0 16925
rect -285 16890 -215 16910
rect -310 16850 -215 16890
rect -155 16890 -85 16910
rect -155 16850 -60 16890
rect -310 16800 -60 16850
rect -310 16760 -215 16800
rect -285 16740 -215 16760
rect -155 16760 -60 16800
rect -155 16740 -85 16760
rect -370 16725 -314 16731
rect -370 16665 -366 16725
rect -285 16715 -85 16740
rect -30 16731 0 16919
rect -56 16725 0 16731
rect -314 16665 -56 16685
rect -4 16665 0 16725
rect -370 16655 0 16665
rect 30 16985 400 16995
rect 30 16925 34 16985
rect 86 16965 344 16985
rect 30 16919 86 16925
rect 30 16731 60 16919
rect 115 16910 315 16935
rect 396 16925 400 16985
rect 344 16919 400 16925
rect 115 16890 185 16910
rect 90 16850 185 16890
rect 245 16890 315 16910
rect 245 16850 340 16890
rect 90 16800 340 16850
rect 90 16760 185 16800
rect 115 16740 185 16760
rect 245 16760 340 16800
rect 245 16740 315 16760
rect 30 16725 86 16731
rect 30 16665 34 16725
rect 115 16715 315 16740
rect 370 16731 400 16919
rect 344 16725 400 16731
rect 86 16665 344 16685
rect 396 16665 400 16725
rect 30 16655 400 16665
rect 430 16985 800 16995
rect 430 16925 434 16985
rect 486 16965 744 16985
rect 430 16919 486 16925
rect 430 16731 460 16919
rect 515 16910 715 16935
rect 796 16925 800 16985
rect 744 16919 800 16925
rect 515 16890 585 16910
rect 490 16850 585 16890
rect 645 16890 715 16910
rect 645 16850 740 16890
rect 490 16800 740 16850
rect 490 16760 585 16800
rect 515 16740 585 16760
rect 645 16760 740 16800
rect 645 16740 715 16760
rect 430 16725 486 16731
rect 430 16665 434 16725
rect 515 16715 715 16740
rect 770 16731 800 16919
rect 744 16725 800 16731
rect 486 16665 744 16685
rect 796 16665 800 16725
rect 430 16655 800 16665
rect 830 16985 1200 16995
rect 830 16925 834 16985
rect 886 16965 1144 16985
rect 830 16919 886 16925
rect 830 16731 860 16919
rect 915 16910 1115 16935
rect 1196 16925 1200 16985
rect 1144 16919 1200 16925
rect 915 16890 985 16910
rect 890 16850 985 16890
rect 1045 16890 1115 16910
rect 1045 16850 1140 16890
rect 890 16800 1140 16850
rect 890 16760 985 16800
rect 915 16740 985 16760
rect 1045 16760 1140 16800
rect 1045 16740 1115 16760
rect 830 16725 886 16731
rect 830 16665 834 16725
rect 915 16715 1115 16740
rect 1170 16731 1200 16919
rect 1144 16725 1200 16731
rect 886 16665 1144 16685
rect 1196 16665 1200 16725
rect 830 16655 1200 16665
rect 1230 16985 1600 16995
rect 1230 16925 1234 16985
rect 1286 16965 1544 16985
rect 1230 16919 1286 16925
rect 1230 16731 1260 16919
rect 1315 16910 1515 16935
rect 1596 16925 1600 16985
rect 1544 16919 1600 16925
rect 1315 16890 1385 16910
rect 1290 16850 1385 16890
rect 1445 16890 1515 16910
rect 1445 16850 1540 16890
rect 1290 16800 1540 16850
rect 1290 16760 1385 16800
rect 1315 16740 1385 16760
rect 1445 16760 1540 16800
rect 1445 16740 1515 16760
rect 1230 16725 1286 16731
rect 1230 16665 1234 16725
rect 1315 16715 1515 16740
rect 1570 16731 1600 16919
rect 1544 16725 1600 16731
rect 1286 16665 1544 16685
rect 1596 16665 1600 16725
rect 1230 16655 1600 16665
rect 1630 16985 2000 16995
rect 1630 16925 1634 16985
rect 1686 16965 1944 16985
rect 1630 16919 1686 16925
rect 1630 16731 1660 16919
rect 1715 16910 1915 16935
rect 1996 16925 2000 16985
rect 1944 16919 2000 16925
rect 1715 16890 1785 16910
rect 1690 16850 1785 16890
rect 1845 16890 1915 16910
rect 1845 16850 1940 16890
rect 1690 16800 1940 16850
rect 1690 16760 1785 16800
rect 1715 16740 1785 16760
rect 1845 16760 1940 16800
rect 1845 16740 1915 16760
rect 1630 16725 1686 16731
rect 1630 16665 1634 16725
rect 1715 16715 1915 16740
rect 1970 16731 2000 16919
rect 1944 16725 2000 16731
rect 1686 16665 1944 16685
rect 1996 16665 2000 16725
rect 1630 16655 2000 16665
rect 2030 16985 2400 16995
rect 2030 16925 2034 16985
rect 2086 16965 2344 16985
rect 2030 16919 2086 16925
rect 2030 16731 2060 16919
rect 2115 16910 2315 16935
rect 2396 16925 2400 16985
rect 2344 16919 2400 16925
rect 2115 16890 2185 16910
rect 2090 16850 2185 16890
rect 2245 16890 2315 16910
rect 2245 16850 2340 16890
rect 2090 16800 2340 16850
rect 2090 16760 2185 16800
rect 2115 16740 2185 16760
rect 2245 16760 2340 16800
rect 2245 16740 2315 16760
rect 2030 16725 2086 16731
rect 2030 16665 2034 16725
rect 2115 16715 2315 16740
rect 2370 16731 2400 16919
rect 2344 16725 2400 16731
rect 2086 16665 2344 16685
rect 2396 16665 2400 16725
rect 2030 16655 2400 16665
rect 2430 16985 2800 16995
rect 2430 16925 2434 16985
rect 2486 16965 2744 16985
rect 2430 16919 2486 16925
rect 2430 16731 2460 16919
rect 2515 16910 2715 16935
rect 2796 16925 2800 16985
rect 2744 16919 2800 16925
rect 2515 16890 2585 16910
rect 2490 16850 2585 16890
rect 2645 16890 2715 16910
rect 2645 16850 2740 16890
rect 2490 16800 2740 16850
rect 2490 16760 2585 16800
rect 2515 16740 2585 16760
rect 2645 16760 2740 16800
rect 2645 16740 2715 16760
rect 2430 16725 2486 16731
rect 2430 16665 2434 16725
rect 2515 16715 2715 16740
rect 2770 16731 2800 16919
rect 2744 16725 2800 16731
rect 2486 16665 2744 16685
rect 2796 16665 2800 16725
rect 2430 16655 2800 16665
rect 2830 16985 3200 16995
rect 2830 16925 2834 16985
rect 2886 16965 3144 16985
rect 2830 16919 2886 16925
rect 2830 16731 2860 16919
rect 2915 16910 3115 16935
rect 3196 16925 3200 16985
rect 3144 16919 3200 16925
rect 2915 16890 2985 16910
rect 2890 16850 2985 16890
rect 3045 16890 3115 16910
rect 3045 16850 3140 16890
rect 2890 16800 3140 16850
rect 2890 16760 2985 16800
rect 2915 16740 2985 16760
rect 3045 16760 3140 16800
rect 3045 16740 3115 16760
rect 2830 16725 2886 16731
rect 2830 16665 2834 16725
rect 2915 16715 3115 16740
rect 3170 16731 3200 16919
rect 3144 16725 3200 16731
rect 2886 16665 3144 16685
rect 3196 16665 3200 16725
rect 2830 16655 3200 16665
rect 3230 16985 3600 16995
rect 3230 16925 3234 16985
rect 3286 16965 3544 16985
rect 3230 16919 3286 16925
rect 3230 16731 3260 16919
rect 3315 16910 3515 16935
rect 3596 16925 3600 16985
rect 3544 16919 3600 16925
rect 3315 16890 3385 16910
rect 3290 16850 3385 16890
rect 3445 16890 3515 16910
rect 3445 16850 3540 16890
rect 3290 16800 3540 16850
rect 3290 16760 3385 16800
rect 3315 16740 3385 16760
rect 3445 16760 3540 16800
rect 3445 16740 3515 16760
rect 3230 16725 3286 16731
rect 3230 16665 3234 16725
rect 3315 16715 3515 16740
rect 3570 16731 3600 16919
rect 3544 16725 3600 16731
rect 3286 16665 3544 16685
rect 3596 16665 3600 16725
rect 3230 16655 3600 16665
rect 3630 16985 4000 16995
rect 3630 16925 3634 16985
rect 3686 16965 3944 16985
rect 3630 16919 3686 16925
rect 3630 16731 3660 16919
rect 3715 16910 3915 16935
rect 3996 16925 4000 16985
rect 3944 16919 4000 16925
rect 3715 16890 3785 16910
rect 3690 16850 3785 16890
rect 3845 16890 3915 16910
rect 3845 16850 3940 16890
rect 3690 16800 3940 16850
rect 3690 16760 3785 16800
rect 3715 16740 3785 16760
rect 3845 16760 3940 16800
rect 3845 16740 3915 16760
rect 3630 16725 3686 16731
rect 3630 16665 3634 16725
rect 3715 16715 3915 16740
rect 3970 16731 4000 16919
rect 3944 16725 4000 16731
rect 3686 16665 3944 16685
rect 3996 16665 4000 16725
rect 3630 16655 4000 16665
rect 4030 16985 4400 16995
rect 4030 16925 4034 16985
rect 4086 16965 4344 16985
rect 4030 16919 4086 16925
rect 4030 16731 4060 16919
rect 4115 16910 4315 16935
rect 4396 16925 4400 16985
rect 4344 16919 4400 16925
rect 4115 16890 4185 16910
rect 4090 16850 4185 16890
rect 4245 16890 4315 16910
rect 4245 16850 4340 16890
rect 4090 16800 4340 16850
rect 4090 16760 4185 16800
rect 4115 16740 4185 16760
rect 4245 16760 4340 16800
rect 4245 16740 4315 16760
rect 4030 16725 4086 16731
rect 4030 16665 4034 16725
rect 4115 16715 4315 16740
rect 4370 16731 4400 16919
rect 4344 16725 4400 16731
rect 4086 16665 4344 16685
rect 4396 16665 4400 16725
rect 4030 16655 4400 16665
rect 4430 16985 4800 16995
rect 4430 16925 4434 16985
rect 4486 16965 4744 16985
rect 4430 16919 4486 16925
rect 4430 16731 4460 16919
rect 4515 16910 4715 16935
rect 4796 16925 4800 16985
rect 4744 16919 4800 16925
rect 4515 16890 4585 16910
rect 4490 16850 4585 16890
rect 4645 16890 4715 16910
rect 4645 16850 4740 16890
rect 4490 16800 4740 16850
rect 4490 16760 4585 16800
rect 4515 16740 4585 16760
rect 4645 16760 4740 16800
rect 4645 16740 4715 16760
rect 4430 16725 4486 16731
rect 4430 16665 4434 16725
rect 4515 16715 4715 16740
rect 4770 16731 4800 16919
rect 4744 16725 4800 16731
rect 4486 16665 4744 16685
rect 4796 16665 4800 16725
rect 4430 16655 4800 16665
rect 4830 16985 5200 16995
rect 4830 16925 4834 16985
rect 4886 16965 5144 16985
rect 4830 16919 4886 16925
rect 4830 16731 4860 16919
rect 4915 16910 5115 16935
rect 5196 16925 5200 16985
rect 5144 16919 5200 16925
rect 4915 16890 4985 16910
rect 4890 16850 4985 16890
rect 5045 16890 5115 16910
rect 5045 16850 5140 16890
rect 4890 16800 5140 16850
rect 4890 16760 4985 16800
rect 4915 16740 4985 16760
rect 5045 16760 5140 16800
rect 5045 16740 5115 16760
rect 4830 16725 4886 16731
rect 4830 16665 4834 16725
rect 4915 16715 5115 16740
rect 5170 16731 5200 16919
rect 5144 16725 5200 16731
rect 4886 16665 5144 16685
rect 5196 16665 5200 16725
rect 4830 16655 5200 16665
rect 5230 16985 5600 16995
rect 5230 16925 5234 16985
rect 5286 16965 5544 16985
rect 5230 16919 5286 16925
rect 5230 16731 5260 16919
rect 5315 16910 5515 16935
rect 5596 16925 5600 16985
rect 5544 16919 5600 16925
rect 5315 16890 5385 16910
rect 5290 16850 5385 16890
rect 5445 16890 5515 16910
rect 5445 16850 5540 16890
rect 5290 16800 5540 16850
rect 5290 16760 5385 16800
rect 5315 16740 5385 16760
rect 5445 16760 5540 16800
rect 5445 16740 5515 16760
rect 5230 16725 5286 16731
rect 5230 16665 5234 16725
rect 5315 16715 5515 16740
rect 5570 16731 5600 16919
rect 5544 16725 5600 16731
rect 5286 16665 5544 16685
rect 5596 16665 5600 16725
rect 5230 16655 5600 16665
rect 5630 16985 6000 16995
rect 5630 16925 5634 16985
rect 5686 16965 5944 16985
rect 5630 16919 5686 16925
rect 5630 16731 5660 16919
rect 5715 16910 5915 16935
rect 5996 16925 6000 16985
rect 5944 16919 6000 16925
rect 5715 16890 5785 16910
rect 5690 16850 5785 16890
rect 5845 16890 5915 16910
rect 5845 16850 5940 16890
rect 5690 16800 5940 16850
rect 5690 16760 5785 16800
rect 5715 16740 5785 16760
rect 5845 16760 5940 16800
rect 5845 16740 5915 16760
rect 5630 16725 5686 16731
rect 5630 16665 5634 16725
rect 5715 16715 5915 16740
rect 5970 16731 6000 16919
rect 5944 16725 6000 16731
rect 5686 16665 5944 16685
rect 5996 16665 6000 16725
rect 5630 16655 6000 16665
rect 6030 16985 6400 16995
rect 6030 16925 6034 16985
rect 6086 16965 6344 16985
rect 6030 16919 6086 16925
rect 6030 16731 6060 16919
rect 6115 16910 6315 16935
rect 6396 16925 6400 16985
rect 6344 16919 6400 16925
rect 6115 16890 6185 16910
rect 6090 16850 6185 16890
rect 6245 16890 6315 16910
rect 6245 16850 6340 16890
rect 6090 16800 6340 16850
rect 6090 16760 6185 16800
rect 6115 16740 6185 16760
rect 6245 16760 6340 16800
rect 6245 16740 6315 16760
rect 6030 16725 6086 16731
rect 6030 16665 6034 16725
rect 6115 16715 6315 16740
rect 6370 16731 6400 16919
rect 6344 16725 6400 16731
rect 6086 16665 6344 16685
rect 6396 16665 6400 16725
rect 6030 16655 6400 16665
rect 6430 16985 6800 16995
rect 6430 16925 6434 16985
rect 6486 16965 6744 16985
rect 6430 16919 6486 16925
rect 6430 16731 6460 16919
rect 6515 16910 6715 16935
rect 6796 16925 6800 16985
rect 6744 16919 6800 16925
rect 6515 16890 6585 16910
rect 6490 16850 6585 16890
rect 6645 16890 6715 16910
rect 6645 16850 6740 16890
rect 6490 16800 6740 16850
rect 6490 16760 6585 16800
rect 6515 16740 6585 16760
rect 6645 16760 6740 16800
rect 6645 16740 6715 16760
rect 6430 16725 6486 16731
rect 6430 16665 6434 16725
rect 6515 16715 6715 16740
rect 6770 16731 6800 16919
rect 6744 16725 6800 16731
rect 6486 16665 6744 16685
rect 6796 16665 6800 16725
rect 6430 16655 6800 16665
rect 6830 16985 7200 16995
rect 6830 16925 6834 16985
rect 6886 16965 7144 16985
rect 6830 16919 6886 16925
rect 6830 16731 6860 16919
rect 6915 16910 7115 16935
rect 7196 16925 7200 16985
rect 7144 16919 7200 16925
rect 6915 16890 6985 16910
rect 6890 16850 6985 16890
rect 7045 16890 7115 16910
rect 7045 16850 7140 16890
rect 6890 16800 7140 16850
rect 6890 16760 6985 16800
rect 6915 16740 6985 16760
rect 7045 16760 7140 16800
rect 7045 16740 7115 16760
rect 6830 16725 6886 16731
rect 6830 16665 6834 16725
rect 6915 16715 7115 16740
rect 7170 16731 7200 16919
rect 7144 16725 7200 16731
rect 6886 16665 7144 16685
rect 7196 16665 7200 16725
rect 6830 16655 7200 16665
rect 7230 16985 7600 16995
rect 7230 16925 7234 16985
rect 7286 16965 7544 16985
rect 7230 16919 7286 16925
rect 7230 16731 7260 16919
rect 7315 16910 7515 16935
rect 7596 16925 7600 16985
rect 7544 16919 7600 16925
rect 7315 16890 7385 16910
rect 7290 16850 7385 16890
rect 7445 16890 7515 16910
rect 7445 16850 7540 16890
rect 7290 16800 7540 16850
rect 7290 16760 7385 16800
rect 7315 16740 7385 16760
rect 7445 16760 7540 16800
rect 7445 16740 7515 16760
rect 7230 16725 7286 16731
rect 7230 16665 7234 16725
rect 7315 16715 7515 16740
rect 7570 16731 7600 16919
rect 7544 16725 7600 16731
rect 7286 16665 7544 16685
rect 7596 16665 7600 16725
rect 7230 16655 7600 16665
rect 7630 16985 8000 16995
rect 7630 16925 7634 16985
rect 7686 16965 7944 16985
rect 7630 16919 7686 16925
rect 7630 16731 7660 16919
rect 7715 16910 7915 16935
rect 7996 16925 8000 16985
rect 7944 16919 8000 16925
rect 7715 16890 7785 16910
rect 7690 16850 7785 16890
rect 7845 16890 7915 16910
rect 7845 16850 7940 16890
rect 7690 16800 7940 16850
rect 7690 16760 7785 16800
rect 7715 16740 7785 16760
rect 7845 16760 7940 16800
rect 7845 16740 7915 16760
rect 7630 16725 7686 16731
rect 7630 16665 7634 16725
rect 7715 16715 7915 16740
rect 7970 16731 8000 16919
rect 7944 16725 8000 16731
rect 7686 16665 7944 16685
rect 7996 16665 8000 16725
rect 7630 16655 8000 16665
rect 8030 16985 8400 16995
rect 8030 16925 8034 16985
rect 8086 16965 8344 16985
rect 8030 16919 8086 16925
rect 8030 16731 8060 16919
rect 8115 16910 8315 16935
rect 8396 16925 8400 16985
rect 8344 16919 8400 16925
rect 8115 16890 8185 16910
rect 8090 16850 8185 16890
rect 8245 16890 8315 16910
rect 8245 16850 8340 16890
rect 8090 16800 8340 16850
rect 8090 16760 8185 16800
rect 8115 16740 8185 16760
rect 8245 16760 8340 16800
rect 8245 16740 8315 16760
rect 8030 16725 8086 16731
rect 8030 16665 8034 16725
rect 8115 16715 8315 16740
rect 8370 16731 8400 16919
rect 8344 16725 8400 16731
rect 8086 16665 8344 16685
rect 8396 16665 8400 16725
rect 8030 16655 8400 16665
rect 8430 16985 8800 16995
rect 8430 16925 8434 16985
rect 8486 16965 8744 16985
rect 8430 16919 8486 16925
rect 8430 16731 8460 16919
rect 8515 16910 8715 16935
rect 8796 16925 8800 16985
rect 8744 16919 8800 16925
rect 8515 16890 8585 16910
rect 8490 16850 8585 16890
rect 8645 16890 8715 16910
rect 8645 16850 8740 16890
rect 8490 16800 8740 16850
rect 8490 16760 8585 16800
rect 8515 16740 8585 16760
rect 8645 16760 8740 16800
rect 8645 16740 8715 16760
rect 8430 16725 8486 16731
rect 8430 16665 8434 16725
rect 8515 16715 8715 16740
rect 8770 16731 8800 16919
rect 8744 16725 8800 16731
rect 8486 16665 8744 16685
rect 8796 16665 8800 16725
rect 8430 16655 8800 16665
rect 8830 16985 9200 16995
rect 8830 16925 8834 16985
rect 8886 16965 9144 16985
rect 8830 16919 8886 16925
rect 8830 16731 8860 16919
rect 8915 16910 9115 16935
rect 9196 16925 9200 16985
rect 9144 16919 9200 16925
rect 8915 16890 8985 16910
rect 8890 16850 8985 16890
rect 9045 16890 9115 16910
rect 9045 16850 9140 16890
rect 8890 16800 9140 16850
rect 8890 16760 8985 16800
rect 8915 16740 8985 16760
rect 9045 16760 9140 16800
rect 9045 16740 9115 16760
rect 8830 16725 8886 16731
rect 8830 16665 8834 16725
rect 8915 16715 9115 16740
rect 9170 16731 9200 16919
rect 9144 16725 9200 16731
rect 8886 16665 9144 16685
rect 9196 16665 9200 16725
rect 8830 16655 9200 16665
rect 9230 16985 9600 16995
rect 9230 16925 9234 16985
rect 9286 16965 9544 16985
rect 9230 16919 9286 16925
rect 9230 16731 9260 16919
rect 9315 16910 9515 16935
rect 9596 16925 9600 16985
rect 9544 16919 9600 16925
rect 9315 16890 9385 16910
rect 9290 16850 9385 16890
rect 9445 16890 9515 16910
rect 9445 16850 9540 16890
rect 9290 16800 9540 16850
rect 9290 16760 9385 16800
rect 9315 16740 9385 16760
rect 9445 16760 9540 16800
rect 9445 16740 9515 16760
rect 9230 16725 9286 16731
rect 9230 16665 9234 16725
rect 9315 16715 9515 16740
rect 9570 16731 9600 16919
rect 9544 16725 9600 16731
rect 9286 16665 9544 16685
rect 9596 16665 9600 16725
rect 9230 16655 9600 16665
rect 9630 16985 10000 16995
rect 9630 16925 9634 16985
rect 9686 16965 9944 16985
rect 9630 16919 9686 16925
rect 9630 16731 9660 16919
rect 9715 16910 9915 16935
rect 9996 16925 10000 16985
rect 9944 16919 10000 16925
rect 9715 16890 9785 16910
rect 9690 16850 9785 16890
rect 9845 16890 9915 16910
rect 9845 16850 9940 16890
rect 9690 16800 9940 16850
rect 9690 16760 9785 16800
rect 9715 16740 9785 16760
rect 9845 16760 9940 16800
rect 9845 16740 9915 16760
rect 9630 16725 9686 16731
rect 9630 16665 9634 16725
rect 9715 16715 9915 16740
rect 9970 16731 10000 16919
rect 9944 16725 10000 16731
rect 9686 16665 9944 16685
rect 9996 16665 10000 16725
rect 9630 16655 10000 16665
rect 10030 16985 10400 16995
rect 10030 16925 10034 16985
rect 10086 16965 10344 16985
rect 10030 16919 10086 16925
rect 10030 16731 10060 16919
rect 10115 16910 10315 16935
rect 10396 16925 10400 16985
rect 10344 16919 10400 16925
rect 10115 16890 10185 16910
rect 10090 16850 10185 16890
rect 10245 16890 10315 16910
rect 10245 16850 10340 16890
rect 10090 16800 10340 16850
rect 10090 16760 10185 16800
rect 10115 16740 10185 16760
rect 10245 16760 10340 16800
rect 10245 16740 10315 16760
rect 10030 16725 10086 16731
rect 10030 16665 10034 16725
rect 10115 16715 10315 16740
rect 10370 16731 10400 16919
rect 10344 16725 10400 16731
rect 10086 16665 10344 16685
rect 10396 16665 10400 16725
rect 10030 16655 10400 16665
rect 10430 16985 10800 16995
rect 10430 16925 10434 16985
rect 10486 16965 10744 16985
rect 10430 16919 10486 16925
rect 10430 16731 10460 16919
rect 10515 16910 10715 16935
rect 10796 16925 10800 16985
rect 10744 16919 10800 16925
rect 10515 16890 10585 16910
rect 10490 16850 10585 16890
rect 10645 16890 10715 16910
rect 10645 16850 10740 16890
rect 10490 16800 10740 16850
rect 10490 16760 10585 16800
rect 10515 16740 10585 16760
rect 10645 16760 10740 16800
rect 10645 16740 10715 16760
rect 10430 16725 10486 16731
rect 10430 16665 10434 16725
rect 10515 16715 10715 16740
rect 10770 16731 10800 16919
rect 10744 16725 10800 16731
rect 10486 16665 10744 16685
rect 10796 16665 10800 16725
rect 10430 16655 10800 16665
rect 10830 16985 11200 16995
rect 10830 16925 10834 16985
rect 10886 16965 11144 16985
rect 10830 16919 10886 16925
rect 10830 16731 10860 16919
rect 10915 16910 11115 16935
rect 11196 16925 11200 16985
rect 11144 16919 11200 16925
rect 10915 16890 10985 16910
rect 10890 16850 10985 16890
rect 11045 16890 11115 16910
rect 11045 16850 11140 16890
rect 10890 16800 11140 16850
rect 10890 16760 10985 16800
rect 10915 16740 10985 16760
rect 11045 16760 11140 16800
rect 11045 16740 11115 16760
rect 10830 16725 10886 16731
rect 10830 16665 10834 16725
rect 10915 16715 11115 16740
rect 11170 16731 11200 16919
rect 11144 16725 11200 16731
rect 10886 16665 11144 16685
rect 11196 16665 11200 16725
rect 10830 16655 11200 16665
rect 11230 16985 11600 16995
rect 11230 16925 11234 16985
rect 11286 16965 11544 16985
rect 11230 16919 11286 16925
rect 11230 16731 11260 16919
rect 11315 16910 11515 16935
rect 11596 16925 11600 16985
rect 11544 16919 11600 16925
rect 11315 16890 11385 16910
rect 11290 16850 11385 16890
rect 11445 16890 11515 16910
rect 11445 16850 11540 16890
rect 11290 16800 11540 16850
rect 11290 16760 11385 16800
rect 11315 16740 11385 16760
rect 11445 16760 11540 16800
rect 11445 16740 11515 16760
rect 11230 16725 11286 16731
rect 11230 16665 11234 16725
rect 11315 16715 11515 16740
rect 11570 16731 11600 16919
rect 11544 16725 11600 16731
rect 11286 16665 11544 16685
rect 11596 16665 11600 16725
rect 11230 16655 11600 16665
rect 11630 16985 12000 16995
rect 11630 16925 11634 16985
rect 11686 16965 11944 16985
rect 11630 16919 11686 16925
rect 11630 16731 11660 16919
rect 11715 16910 11915 16935
rect 11996 16925 12000 16985
rect 11944 16919 12000 16925
rect 11715 16890 11785 16910
rect 11690 16850 11785 16890
rect 11845 16890 11915 16910
rect 11845 16850 11940 16890
rect 11690 16800 11940 16850
rect 11690 16760 11785 16800
rect 11715 16740 11785 16760
rect 11845 16760 11940 16800
rect 11845 16740 11915 16760
rect 11630 16725 11686 16731
rect 11630 16665 11634 16725
rect 11715 16715 11915 16740
rect 11970 16731 12000 16919
rect 11944 16725 12000 16731
rect 11686 16665 11944 16685
rect 11996 16665 12000 16725
rect 11630 16655 12000 16665
rect 12030 16985 12400 16995
rect 12030 16925 12034 16985
rect 12086 16965 12344 16985
rect 12030 16919 12086 16925
rect 12030 16731 12060 16919
rect 12115 16910 12315 16935
rect 12396 16925 12400 16985
rect 12344 16919 12400 16925
rect 12115 16890 12185 16910
rect 12090 16850 12185 16890
rect 12245 16890 12315 16910
rect 12245 16850 12340 16890
rect 12090 16800 12340 16850
rect 12090 16760 12185 16800
rect 12115 16740 12185 16760
rect 12245 16760 12340 16800
rect 12245 16740 12315 16760
rect 12030 16725 12086 16731
rect 12030 16665 12034 16725
rect 12115 16715 12315 16740
rect 12370 16731 12400 16919
rect 12344 16725 12400 16731
rect 12086 16665 12344 16685
rect 12396 16665 12400 16725
rect 12030 16655 12400 16665
rect 12430 16985 12800 16995
rect 12430 16925 12434 16985
rect 12486 16965 12744 16985
rect 12430 16919 12486 16925
rect 12430 16731 12460 16919
rect 12515 16910 12715 16935
rect 12796 16925 12800 16985
rect 12744 16919 12800 16925
rect 12515 16890 12585 16910
rect 12490 16850 12585 16890
rect 12645 16890 12715 16910
rect 12645 16850 12740 16890
rect 12490 16800 12740 16850
rect 12490 16760 12585 16800
rect 12515 16740 12585 16760
rect 12645 16760 12740 16800
rect 12645 16740 12715 16760
rect 12430 16725 12486 16731
rect 12430 16665 12434 16725
rect 12515 16715 12715 16740
rect 12770 16731 12800 16919
rect 12744 16725 12800 16731
rect 12486 16665 12744 16685
rect 12796 16665 12800 16725
rect 12430 16655 12800 16665
rect 12830 16985 13200 16995
rect 12830 16925 12834 16985
rect 12886 16965 13144 16985
rect 12830 16919 12886 16925
rect 12830 16731 12860 16919
rect 12915 16910 13115 16935
rect 13196 16925 13200 16985
rect 13144 16919 13200 16925
rect 12915 16890 12985 16910
rect 12890 16850 12985 16890
rect 13045 16890 13115 16910
rect 13045 16850 13140 16890
rect 12890 16800 13140 16850
rect 12890 16760 12985 16800
rect 12915 16740 12985 16760
rect 13045 16760 13140 16800
rect 13045 16740 13115 16760
rect 12830 16725 12886 16731
rect 12830 16665 12834 16725
rect 12915 16715 13115 16740
rect 13170 16731 13200 16919
rect 13144 16725 13200 16731
rect 12886 16665 13144 16685
rect 13196 16665 13200 16725
rect 12830 16655 13200 16665
rect -370 16615 0 16625
rect -370 16555 -366 16615
rect -314 16595 -56 16615
rect -370 16549 -314 16555
rect -370 16361 -340 16549
rect -285 16540 -85 16565
rect -4 16555 0 16615
rect -56 16549 0 16555
rect -285 16520 -215 16540
rect -310 16480 -215 16520
rect -155 16520 -85 16540
rect -155 16480 -60 16520
rect -310 16430 -60 16480
rect -310 16390 -215 16430
rect -285 16370 -215 16390
rect -155 16390 -60 16430
rect -155 16370 -85 16390
rect -370 16355 -314 16361
rect -370 16295 -366 16355
rect -285 16345 -85 16370
rect -30 16361 0 16549
rect -56 16355 0 16361
rect -314 16295 -56 16315
rect -4 16295 0 16355
rect -370 16285 0 16295
rect 30 16615 400 16625
rect 30 16555 34 16615
rect 86 16595 344 16615
rect 30 16549 86 16555
rect 30 16361 60 16549
rect 115 16540 315 16565
rect 396 16555 400 16615
rect 344 16549 400 16555
rect 115 16520 185 16540
rect 90 16480 185 16520
rect 245 16520 315 16540
rect 245 16480 340 16520
rect 90 16430 340 16480
rect 90 16390 185 16430
rect 115 16370 185 16390
rect 245 16390 340 16430
rect 245 16370 315 16390
rect 30 16355 86 16361
rect 30 16295 34 16355
rect 115 16345 315 16370
rect 370 16361 400 16549
rect 344 16355 400 16361
rect 86 16295 344 16315
rect 396 16295 400 16355
rect 30 16285 400 16295
rect 430 16615 800 16625
rect 430 16555 434 16615
rect 486 16595 744 16615
rect 430 16549 486 16555
rect 430 16361 460 16549
rect 515 16540 715 16565
rect 796 16555 800 16615
rect 744 16549 800 16555
rect 515 16520 585 16540
rect 490 16480 585 16520
rect 645 16520 715 16540
rect 645 16480 740 16520
rect 490 16430 740 16480
rect 490 16390 585 16430
rect 515 16370 585 16390
rect 645 16390 740 16430
rect 645 16370 715 16390
rect 430 16355 486 16361
rect 430 16295 434 16355
rect 515 16345 715 16370
rect 770 16361 800 16549
rect 744 16355 800 16361
rect 486 16295 744 16315
rect 796 16295 800 16355
rect 430 16285 800 16295
rect 830 16615 1200 16625
rect 830 16555 834 16615
rect 886 16595 1144 16615
rect 830 16549 886 16555
rect 830 16361 860 16549
rect 915 16540 1115 16565
rect 1196 16555 1200 16615
rect 1144 16549 1200 16555
rect 915 16520 985 16540
rect 890 16480 985 16520
rect 1045 16520 1115 16540
rect 1045 16480 1140 16520
rect 890 16430 1140 16480
rect 890 16390 985 16430
rect 915 16370 985 16390
rect 1045 16390 1140 16430
rect 1045 16370 1115 16390
rect 830 16355 886 16361
rect 830 16295 834 16355
rect 915 16345 1115 16370
rect 1170 16361 1200 16549
rect 1144 16355 1200 16361
rect 886 16295 1144 16315
rect 1196 16295 1200 16355
rect 830 16285 1200 16295
rect 1230 16615 1600 16625
rect 1230 16555 1234 16615
rect 1286 16595 1544 16615
rect 1230 16549 1286 16555
rect 1230 16361 1260 16549
rect 1315 16540 1515 16565
rect 1596 16555 1600 16615
rect 1544 16549 1600 16555
rect 1315 16520 1385 16540
rect 1290 16480 1385 16520
rect 1445 16520 1515 16540
rect 1445 16480 1540 16520
rect 1290 16430 1540 16480
rect 1290 16390 1385 16430
rect 1315 16370 1385 16390
rect 1445 16390 1540 16430
rect 1445 16370 1515 16390
rect 1230 16355 1286 16361
rect 1230 16295 1234 16355
rect 1315 16345 1515 16370
rect 1570 16361 1600 16549
rect 1544 16355 1600 16361
rect 1286 16295 1544 16315
rect 1596 16295 1600 16355
rect 1230 16285 1600 16295
rect 1630 16615 2000 16625
rect 1630 16555 1634 16615
rect 1686 16595 1944 16615
rect 1630 16549 1686 16555
rect 1630 16361 1660 16549
rect 1715 16540 1915 16565
rect 1996 16555 2000 16615
rect 1944 16549 2000 16555
rect 1715 16520 1785 16540
rect 1690 16480 1785 16520
rect 1845 16520 1915 16540
rect 1845 16480 1940 16520
rect 1690 16430 1940 16480
rect 1690 16390 1785 16430
rect 1715 16370 1785 16390
rect 1845 16390 1940 16430
rect 1845 16370 1915 16390
rect 1630 16355 1686 16361
rect 1630 16295 1634 16355
rect 1715 16345 1915 16370
rect 1970 16361 2000 16549
rect 1944 16355 2000 16361
rect 1686 16295 1944 16315
rect 1996 16295 2000 16355
rect 1630 16285 2000 16295
rect 2030 16615 2400 16625
rect 2030 16555 2034 16615
rect 2086 16595 2344 16615
rect 2030 16549 2086 16555
rect 2030 16361 2060 16549
rect 2115 16540 2315 16565
rect 2396 16555 2400 16615
rect 2344 16549 2400 16555
rect 2115 16520 2185 16540
rect 2090 16480 2185 16520
rect 2245 16520 2315 16540
rect 2245 16480 2340 16520
rect 2090 16430 2340 16480
rect 2090 16390 2185 16430
rect 2115 16370 2185 16390
rect 2245 16390 2340 16430
rect 2245 16370 2315 16390
rect 2030 16355 2086 16361
rect 2030 16295 2034 16355
rect 2115 16345 2315 16370
rect 2370 16361 2400 16549
rect 2344 16355 2400 16361
rect 2086 16295 2344 16315
rect 2396 16295 2400 16355
rect 2030 16285 2400 16295
rect 2430 16615 2800 16625
rect 2430 16555 2434 16615
rect 2486 16595 2744 16615
rect 2430 16549 2486 16555
rect 2430 16361 2460 16549
rect 2515 16540 2715 16565
rect 2796 16555 2800 16615
rect 2744 16549 2800 16555
rect 2515 16520 2585 16540
rect 2490 16480 2585 16520
rect 2645 16520 2715 16540
rect 2645 16480 2740 16520
rect 2490 16430 2740 16480
rect 2490 16390 2585 16430
rect 2515 16370 2585 16390
rect 2645 16390 2740 16430
rect 2645 16370 2715 16390
rect 2430 16355 2486 16361
rect 2430 16295 2434 16355
rect 2515 16345 2715 16370
rect 2770 16361 2800 16549
rect 2744 16355 2800 16361
rect 2486 16295 2744 16315
rect 2796 16295 2800 16355
rect 2430 16285 2800 16295
rect 2830 16615 3200 16625
rect 2830 16555 2834 16615
rect 2886 16595 3144 16615
rect 2830 16549 2886 16555
rect 2830 16361 2860 16549
rect 2915 16540 3115 16565
rect 3196 16555 3200 16615
rect 3144 16549 3200 16555
rect 2915 16520 2985 16540
rect 2890 16480 2985 16520
rect 3045 16520 3115 16540
rect 3045 16480 3140 16520
rect 2890 16430 3140 16480
rect 2890 16390 2985 16430
rect 2915 16370 2985 16390
rect 3045 16390 3140 16430
rect 3045 16370 3115 16390
rect 2830 16355 2886 16361
rect 2830 16295 2834 16355
rect 2915 16345 3115 16370
rect 3170 16361 3200 16549
rect 3144 16355 3200 16361
rect 2886 16295 3144 16315
rect 3196 16295 3200 16355
rect 2830 16285 3200 16295
rect 3230 16615 3600 16625
rect 3230 16555 3234 16615
rect 3286 16595 3544 16615
rect 3230 16549 3286 16555
rect 3230 16361 3260 16549
rect 3315 16540 3515 16565
rect 3596 16555 3600 16615
rect 3544 16549 3600 16555
rect 3315 16520 3385 16540
rect 3290 16480 3385 16520
rect 3445 16520 3515 16540
rect 3445 16480 3540 16520
rect 3290 16430 3540 16480
rect 3290 16390 3385 16430
rect 3315 16370 3385 16390
rect 3445 16390 3540 16430
rect 3445 16370 3515 16390
rect 3230 16355 3286 16361
rect 3230 16295 3234 16355
rect 3315 16345 3515 16370
rect 3570 16361 3600 16549
rect 3544 16355 3600 16361
rect 3286 16295 3544 16315
rect 3596 16295 3600 16355
rect 3230 16285 3600 16295
rect 3630 16615 4000 16625
rect 3630 16555 3634 16615
rect 3686 16595 3944 16615
rect 3630 16549 3686 16555
rect 3630 16361 3660 16549
rect 3715 16540 3915 16565
rect 3996 16555 4000 16615
rect 3944 16549 4000 16555
rect 3715 16520 3785 16540
rect 3690 16480 3785 16520
rect 3845 16520 3915 16540
rect 3845 16480 3940 16520
rect 3690 16430 3940 16480
rect 3690 16390 3785 16430
rect 3715 16370 3785 16390
rect 3845 16390 3940 16430
rect 3845 16370 3915 16390
rect 3630 16355 3686 16361
rect 3630 16295 3634 16355
rect 3715 16345 3915 16370
rect 3970 16361 4000 16549
rect 3944 16355 4000 16361
rect 3686 16295 3944 16315
rect 3996 16295 4000 16355
rect 3630 16285 4000 16295
rect 4030 16615 4400 16625
rect 4030 16555 4034 16615
rect 4086 16595 4344 16615
rect 4030 16549 4086 16555
rect 4030 16361 4060 16549
rect 4115 16540 4315 16565
rect 4396 16555 4400 16615
rect 4344 16549 4400 16555
rect 4115 16520 4185 16540
rect 4090 16480 4185 16520
rect 4245 16520 4315 16540
rect 4245 16480 4340 16520
rect 4090 16430 4340 16480
rect 4090 16390 4185 16430
rect 4115 16370 4185 16390
rect 4245 16390 4340 16430
rect 4245 16370 4315 16390
rect 4030 16355 4086 16361
rect 4030 16295 4034 16355
rect 4115 16345 4315 16370
rect 4370 16361 4400 16549
rect 4344 16355 4400 16361
rect 4086 16295 4344 16315
rect 4396 16295 4400 16355
rect 4030 16285 4400 16295
rect 4430 16615 4800 16625
rect 4430 16555 4434 16615
rect 4486 16595 4744 16615
rect 4430 16549 4486 16555
rect 4430 16361 4460 16549
rect 4515 16540 4715 16565
rect 4796 16555 4800 16615
rect 4744 16549 4800 16555
rect 4515 16520 4585 16540
rect 4490 16480 4585 16520
rect 4645 16520 4715 16540
rect 4645 16480 4740 16520
rect 4490 16430 4740 16480
rect 4490 16390 4585 16430
rect 4515 16370 4585 16390
rect 4645 16390 4740 16430
rect 4645 16370 4715 16390
rect 4430 16355 4486 16361
rect 4430 16295 4434 16355
rect 4515 16345 4715 16370
rect 4770 16361 4800 16549
rect 4744 16355 4800 16361
rect 4486 16295 4744 16315
rect 4796 16295 4800 16355
rect 4430 16285 4800 16295
rect 4830 16615 5200 16625
rect 4830 16555 4834 16615
rect 4886 16595 5144 16615
rect 4830 16549 4886 16555
rect 4830 16361 4860 16549
rect 4915 16540 5115 16565
rect 5196 16555 5200 16615
rect 5144 16549 5200 16555
rect 4915 16520 4985 16540
rect 4890 16480 4985 16520
rect 5045 16520 5115 16540
rect 5045 16480 5140 16520
rect 4890 16430 5140 16480
rect 4890 16390 4985 16430
rect 4915 16370 4985 16390
rect 5045 16390 5140 16430
rect 5045 16370 5115 16390
rect 4830 16355 4886 16361
rect 4830 16295 4834 16355
rect 4915 16345 5115 16370
rect 5170 16361 5200 16549
rect 5144 16355 5200 16361
rect 4886 16295 5144 16315
rect 5196 16295 5200 16355
rect 4830 16285 5200 16295
rect 5230 16615 5600 16625
rect 5230 16555 5234 16615
rect 5286 16595 5544 16615
rect 5230 16549 5286 16555
rect 5230 16361 5260 16549
rect 5315 16540 5515 16565
rect 5596 16555 5600 16615
rect 5544 16549 5600 16555
rect 5315 16520 5385 16540
rect 5290 16480 5385 16520
rect 5445 16520 5515 16540
rect 5445 16480 5540 16520
rect 5290 16430 5540 16480
rect 5290 16390 5385 16430
rect 5315 16370 5385 16390
rect 5445 16390 5540 16430
rect 5445 16370 5515 16390
rect 5230 16355 5286 16361
rect 5230 16295 5234 16355
rect 5315 16345 5515 16370
rect 5570 16361 5600 16549
rect 5544 16355 5600 16361
rect 5286 16295 5544 16315
rect 5596 16295 5600 16355
rect 5230 16285 5600 16295
rect 5630 16615 6000 16625
rect 5630 16555 5634 16615
rect 5686 16595 5944 16615
rect 5630 16549 5686 16555
rect 5630 16361 5660 16549
rect 5715 16540 5915 16565
rect 5996 16555 6000 16615
rect 5944 16549 6000 16555
rect 5715 16520 5785 16540
rect 5690 16480 5785 16520
rect 5845 16520 5915 16540
rect 5845 16480 5940 16520
rect 5690 16430 5940 16480
rect 5690 16390 5785 16430
rect 5715 16370 5785 16390
rect 5845 16390 5940 16430
rect 5845 16370 5915 16390
rect 5630 16355 5686 16361
rect 5630 16295 5634 16355
rect 5715 16345 5915 16370
rect 5970 16361 6000 16549
rect 5944 16355 6000 16361
rect 5686 16295 5944 16315
rect 5996 16295 6000 16355
rect 5630 16285 6000 16295
rect 6030 16615 6400 16625
rect 6030 16555 6034 16615
rect 6086 16595 6344 16615
rect 6030 16549 6086 16555
rect 6030 16361 6060 16549
rect 6115 16540 6315 16565
rect 6396 16555 6400 16615
rect 6344 16549 6400 16555
rect 6115 16520 6185 16540
rect 6090 16480 6185 16520
rect 6245 16520 6315 16540
rect 6245 16480 6340 16520
rect 6090 16430 6340 16480
rect 6090 16390 6185 16430
rect 6115 16370 6185 16390
rect 6245 16390 6340 16430
rect 6245 16370 6315 16390
rect 6030 16355 6086 16361
rect 6030 16295 6034 16355
rect 6115 16345 6315 16370
rect 6370 16361 6400 16549
rect 6344 16355 6400 16361
rect 6086 16295 6344 16315
rect 6396 16295 6400 16355
rect 6030 16285 6400 16295
rect 6430 16615 6800 16625
rect 6430 16555 6434 16615
rect 6486 16595 6744 16615
rect 6430 16549 6486 16555
rect 6430 16361 6460 16549
rect 6515 16540 6715 16565
rect 6796 16555 6800 16615
rect 6744 16549 6800 16555
rect 6515 16520 6585 16540
rect 6490 16480 6585 16520
rect 6645 16520 6715 16540
rect 6645 16480 6740 16520
rect 6490 16430 6740 16480
rect 6490 16390 6585 16430
rect 6515 16370 6585 16390
rect 6645 16390 6740 16430
rect 6645 16370 6715 16390
rect 6430 16355 6486 16361
rect 6430 16295 6434 16355
rect 6515 16345 6715 16370
rect 6770 16361 6800 16549
rect 6744 16355 6800 16361
rect 6486 16295 6744 16315
rect 6796 16295 6800 16355
rect 6430 16285 6800 16295
rect 6830 16615 7200 16625
rect 6830 16555 6834 16615
rect 6886 16595 7144 16615
rect 6830 16549 6886 16555
rect 6830 16361 6860 16549
rect 6915 16540 7115 16565
rect 7196 16555 7200 16615
rect 7144 16549 7200 16555
rect 6915 16520 6985 16540
rect 6890 16480 6985 16520
rect 7045 16520 7115 16540
rect 7045 16480 7140 16520
rect 6890 16430 7140 16480
rect 6890 16390 6985 16430
rect 6915 16370 6985 16390
rect 7045 16390 7140 16430
rect 7045 16370 7115 16390
rect 6830 16355 6886 16361
rect 6830 16295 6834 16355
rect 6915 16345 7115 16370
rect 7170 16361 7200 16549
rect 7144 16355 7200 16361
rect 6886 16295 7144 16315
rect 7196 16295 7200 16355
rect 6830 16285 7200 16295
rect 7230 16615 7600 16625
rect 7230 16555 7234 16615
rect 7286 16595 7544 16615
rect 7230 16549 7286 16555
rect 7230 16361 7260 16549
rect 7315 16540 7515 16565
rect 7596 16555 7600 16615
rect 7544 16549 7600 16555
rect 7315 16520 7385 16540
rect 7290 16480 7385 16520
rect 7445 16520 7515 16540
rect 7445 16480 7540 16520
rect 7290 16430 7540 16480
rect 7290 16390 7385 16430
rect 7315 16370 7385 16390
rect 7445 16390 7540 16430
rect 7445 16370 7515 16390
rect 7230 16355 7286 16361
rect 7230 16295 7234 16355
rect 7315 16345 7515 16370
rect 7570 16361 7600 16549
rect 7544 16355 7600 16361
rect 7286 16295 7544 16315
rect 7596 16295 7600 16355
rect 7230 16285 7600 16295
rect 7630 16615 8000 16625
rect 7630 16555 7634 16615
rect 7686 16595 7944 16615
rect 7630 16549 7686 16555
rect 7630 16361 7660 16549
rect 7715 16540 7915 16565
rect 7996 16555 8000 16615
rect 7944 16549 8000 16555
rect 7715 16520 7785 16540
rect 7690 16480 7785 16520
rect 7845 16520 7915 16540
rect 7845 16480 7940 16520
rect 7690 16430 7940 16480
rect 7690 16390 7785 16430
rect 7715 16370 7785 16390
rect 7845 16390 7940 16430
rect 7845 16370 7915 16390
rect 7630 16355 7686 16361
rect 7630 16295 7634 16355
rect 7715 16345 7915 16370
rect 7970 16361 8000 16549
rect 7944 16355 8000 16361
rect 7686 16295 7944 16315
rect 7996 16295 8000 16355
rect 7630 16285 8000 16295
rect 8030 16615 8400 16625
rect 8030 16555 8034 16615
rect 8086 16595 8344 16615
rect 8030 16549 8086 16555
rect 8030 16361 8060 16549
rect 8115 16540 8315 16565
rect 8396 16555 8400 16615
rect 8344 16549 8400 16555
rect 8115 16520 8185 16540
rect 8090 16480 8185 16520
rect 8245 16520 8315 16540
rect 8245 16480 8340 16520
rect 8090 16430 8340 16480
rect 8090 16390 8185 16430
rect 8115 16370 8185 16390
rect 8245 16390 8340 16430
rect 8245 16370 8315 16390
rect 8030 16355 8086 16361
rect 8030 16295 8034 16355
rect 8115 16345 8315 16370
rect 8370 16361 8400 16549
rect 8344 16355 8400 16361
rect 8086 16295 8344 16315
rect 8396 16295 8400 16355
rect 8030 16285 8400 16295
rect 8430 16615 8800 16625
rect 8430 16555 8434 16615
rect 8486 16595 8744 16615
rect 8430 16549 8486 16555
rect 8430 16361 8460 16549
rect 8515 16540 8715 16565
rect 8796 16555 8800 16615
rect 8744 16549 8800 16555
rect 8515 16520 8585 16540
rect 8490 16480 8585 16520
rect 8645 16520 8715 16540
rect 8645 16480 8740 16520
rect 8490 16430 8740 16480
rect 8490 16390 8585 16430
rect 8515 16370 8585 16390
rect 8645 16390 8740 16430
rect 8645 16370 8715 16390
rect 8430 16355 8486 16361
rect 8430 16295 8434 16355
rect 8515 16345 8715 16370
rect 8770 16361 8800 16549
rect 8744 16355 8800 16361
rect 8486 16295 8744 16315
rect 8796 16295 8800 16355
rect 8430 16285 8800 16295
rect 8830 16615 9200 16625
rect 8830 16555 8834 16615
rect 8886 16595 9144 16615
rect 8830 16549 8886 16555
rect 8830 16361 8860 16549
rect 8915 16540 9115 16565
rect 9196 16555 9200 16615
rect 9144 16549 9200 16555
rect 8915 16520 8985 16540
rect 8890 16480 8985 16520
rect 9045 16520 9115 16540
rect 9045 16480 9140 16520
rect 8890 16430 9140 16480
rect 8890 16390 8985 16430
rect 8915 16370 8985 16390
rect 9045 16390 9140 16430
rect 9045 16370 9115 16390
rect 8830 16355 8886 16361
rect 8830 16295 8834 16355
rect 8915 16345 9115 16370
rect 9170 16361 9200 16549
rect 9144 16355 9200 16361
rect 8886 16295 9144 16315
rect 9196 16295 9200 16355
rect 8830 16285 9200 16295
rect 9230 16615 9600 16625
rect 9230 16555 9234 16615
rect 9286 16595 9544 16615
rect 9230 16549 9286 16555
rect 9230 16361 9260 16549
rect 9315 16540 9515 16565
rect 9596 16555 9600 16615
rect 9544 16549 9600 16555
rect 9315 16520 9385 16540
rect 9290 16480 9385 16520
rect 9445 16520 9515 16540
rect 9445 16480 9540 16520
rect 9290 16430 9540 16480
rect 9290 16390 9385 16430
rect 9315 16370 9385 16390
rect 9445 16390 9540 16430
rect 9445 16370 9515 16390
rect 9230 16355 9286 16361
rect 9230 16295 9234 16355
rect 9315 16345 9515 16370
rect 9570 16361 9600 16549
rect 9544 16355 9600 16361
rect 9286 16295 9544 16315
rect 9596 16295 9600 16355
rect 9230 16285 9600 16295
rect 9630 16615 10000 16625
rect 9630 16555 9634 16615
rect 9686 16595 9944 16615
rect 9630 16549 9686 16555
rect 9630 16361 9660 16549
rect 9715 16540 9915 16565
rect 9996 16555 10000 16615
rect 9944 16549 10000 16555
rect 9715 16520 9785 16540
rect 9690 16480 9785 16520
rect 9845 16520 9915 16540
rect 9845 16480 9940 16520
rect 9690 16430 9940 16480
rect 9690 16390 9785 16430
rect 9715 16370 9785 16390
rect 9845 16390 9940 16430
rect 9845 16370 9915 16390
rect 9630 16355 9686 16361
rect 9630 16295 9634 16355
rect 9715 16345 9915 16370
rect 9970 16361 10000 16549
rect 9944 16355 10000 16361
rect 9686 16295 9944 16315
rect 9996 16295 10000 16355
rect 9630 16285 10000 16295
rect 10030 16615 10400 16625
rect 10030 16555 10034 16615
rect 10086 16595 10344 16615
rect 10030 16549 10086 16555
rect 10030 16361 10060 16549
rect 10115 16540 10315 16565
rect 10396 16555 10400 16615
rect 10344 16549 10400 16555
rect 10115 16520 10185 16540
rect 10090 16480 10185 16520
rect 10245 16520 10315 16540
rect 10245 16480 10340 16520
rect 10090 16430 10340 16480
rect 10090 16390 10185 16430
rect 10115 16370 10185 16390
rect 10245 16390 10340 16430
rect 10245 16370 10315 16390
rect 10030 16355 10086 16361
rect 10030 16295 10034 16355
rect 10115 16345 10315 16370
rect 10370 16361 10400 16549
rect 10344 16355 10400 16361
rect 10086 16295 10344 16315
rect 10396 16295 10400 16355
rect 10030 16285 10400 16295
rect 10430 16615 10800 16625
rect 10430 16555 10434 16615
rect 10486 16595 10744 16615
rect 10430 16549 10486 16555
rect 10430 16361 10460 16549
rect 10515 16540 10715 16565
rect 10796 16555 10800 16615
rect 10744 16549 10800 16555
rect 10515 16520 10585 16540
rect 10490 16480 10585 16520
rect 10645 16520 10715 16540
rect 10645 16480 10740 16520
rect 10490 16430 10740 16480
rect 10490 16390 10585 16430
rect 10515 16370 10585 16390
rect 10645 16390 10740 16430
rect 10645 16370 10715 16390
rect 10430 16355 10486 16361
rect 10430 16295 10434 16355
rect 10515 16345 10715 16370
rect 10770 16361 10800 16549
rect 10744 16355 10800 16361
rect 10486 16295 10744 16315
rect 10796 16295 10800 16355
rect 10430 16285 10800 16295
rect 10830 16615 11200 16625
rect 10830 16555 10834 16615
rect 10886 16595 11144 16615
rect 10830 16549 10886 16555
rect 10830 16361 10860 16549
rect 10915 16540 11115 16565
rect 11196 16555 11200 16615
rect 11144 16549 11200 16555
rect 10915 16520 10985 16540
rect 10890 16480 10985 16520
rect 11045 16520 11115 16540
rect 11045 16480 11140 16520
rect 10890 16430 11140 16480
rect 10890 16390 10985 16430
rect 10915 16370 10985 16390
rect 11045 16390 11140 16430
rect 11045 16370 11115 16390
rect 10830 16355 10886 16361
rect 10830 16295 10834 16355
rect 10915 16345 11115 16370
rect 11170 16361 11200 16549
rect 11144 16355 11200 16361
rect 10886 16295 11144 16315
rect 11196 16295 11200 16355
rect 10830 16285 11200 16295
rect 11230 16615 11600 16625
rect 11230 16555 11234 16615
rect 11286 16595 11544 16615
rect 11230 16549 11286 16555
rect 11230 16361 11260 16549
rect 11315 16540 11515 16565
rect 11596 16555 11600 16615
rect 11544 16549 11600 16555
rect 11315 16520 11385 16540
rect 11290 16480 11385 16520
rect 11445 16520 11515 16540
rect 11445 16480 11540 16520
rect 11290 16430 11540 16480
rect 11290 16390 11385 16430
rect 11315 16370 11385 16390
rect 11445 16390 11540 16430
rect 11445 16370 11515 16390
rect 11230 16355 11286 16361
rect 11230 16295 11234 16355
rect 11315 16345 11515 16370
rect 11570 16361 11600 16549
rect 11544 16355 11600 16361
rect 11286 16295 11544 16315
rect 11596 16295 11600 16355
rect 11230 16285 11600 16295
rect 11630 16615 12000 16625
rect 11630 16555 11634 16615
rect 11686 16595 11944 16615
rect 11630 16549 11686 16555
rect 11630 16361 11660 16549
rect 11715 16540 11915 16565
rect 11996 16555 12000 16615
rect 11944 16549 12000 16555
rect 11715 16520 11785 16540
rect 11690 16480 11785 16520
rect 11845 16520 11915 16540
rect 11845 16480 11940 16520
rect 11690 16430 11940 16480
rect 11690 16390 11785 16430
rect 11715 16370 11785 16390
rect 11845 16390 11940 16430
rect 11845 16370 11915 16390
rect 11630 16355 11686 16361
rect 11630 16295 11634 16355
rect 11715 16345 11915 16370
rect 11970 16361 12000 16549
rect 11944 16355 12000 16361
rect 11686 16295 11944 16315
rect 11996 16295 12000 16355
rect 11630 16285 12000 16295
rect 12030 16615 12400 16625
rect 12030 16555 12034 16615
rect 12086 16595 12344 16615
rect 12030 16549 12086 16555
rect 12030 16361 12060 16549
rect 12115 16540 12315 16565
rect 12396 16555 12400 16615
rect 12344 16549 12400 16555
rect 12115 16520 12185 16540
rect 12090 16480 12185 16520
rect 12245 16520 12315 16540
rect 12245 16480 12340 16520
rect 12090 16430 12340 16480
rect 12090 16390 12185 16430
rect 12115 16370 12185 16390
rect 12245 16390 12340 16430
rect 12245 16370 12315 16390
rect 12030 16355 12086 16361
rect 12030 16295 12034 16355
rect 12115 16345 12315 16370
rect 12370 16361 12400 16549
rect 12344 16355 12400 16361
rect 12086 16295 12344 16315
rect 12396 16295 12400 16355
rect 12030 16285 12400 16295
rect 12430 16615 12800 16625
rect 12430 16555 12434 16615
rect 12486 16595 12744 16615
rect 12430 16549 12486 16555
rect 12430 16361 12460 16549
rect 12515 16540 12715 16565
rect 12796 16555 12800 16615
rect 12744 16549 12800 16555
rect 12515 16520 12585 16540
rect 12490 16480 12585 16520
rect 12645 16520 12715 16540
rect 12645 16480 12740 16520
rect 12490 16430 12740 16480
rect 12490 16390 12585 16430
rect 12515 16370 12585 16390
rect 12645 16390 12740 16430
rect 12645 16370 12715 16390
rect 12430 16355 12486 16361
rect 12430 16295 12434 16355
rect 12515 16345 12715 16370
rect 12770 16361 12800 16549
rect 12744 16355 12800 16361
rect 12486 16295 12744 16315
rect 12796 16295 12800 16355
rect 12430 16285 12800 16295
rect 12830 16615 13200 16625
rect 12830 16555 12834 16615
rect 12886 16595 13144 16615
rect 12830 16549 12886 16555
rect 12830 16361 12860 16549
rect 12915 16540 13115 16565
rect 13196 16555 13200 16615
rect 13144 16549 13200 16555
rect 12915 16520 12985 16540
rect 12890 16480 12985 16520
rect 13045 16520 13115 16540
rect 13045 16480 13140 16520
rect 12890 16430 13140 16480
rect 12890 16390 12985 16430
rect 12915 16370 12985 16390
rect 13045 16390 13140 16430
rect 13045 16370 13115 16390
rect 12830 16355 12886 16361
rect 12830 16295 12834 16355
rect 12915 16345 13115 16370
rect 13170 16361 13200 16549
rect 13144 16355 13200 16361
rect 12886 16295 13144 16315
rect 13196 16295 13200 16355
rect 12830 16285 13200 16295
rect -370 16245 0 16255
rect -370 16185 -366 16245
rect -314 16225 -56 16245
rect -370 16179 -314 16185
rect -370 15991 -340 16179
rect -285 16170 -85 16195
rect -4 16185 0 16245
rect -56 16179 0 16185
rect -285 16150 -215 16170
rect -310 16110 -215 16150
rect -155 16150 -85 16170
rect -155 16110 -60 16150
rect -310 16060 -60 16110
rect -310 16020 -215 16060
rect -285 16000 -215 16020
rect -155 16020 -60 16060
rect -155 16000 -85 16020
rect -370 15985 -314 15991
rect -370 15925 -366 15985
rect -285 15975 -85 16000
rect -30 15991 0 16179
rect -56 15985 0 15991
rect -314 15925 -56 15945
rect -4 15925 0 15985
rect -370 15915 0 15925
rect 30 16245 400 16255
rect 30 16185 34 16245
rect 86 16225 344 16245
rect 30 16179 86 16185
rect 30 15991 60 16179
rect 115 16170 315 16195
rect 396 16185 400 16245
rect 344 16179 400 16185
rect 115 16150 185 16170
rect 90 16110 185 16150
rect 245 16150 315 16170
rect 245 16110 340 16150
rect 90 16060 340 16110
rect 90 16020 185 16060
rect 115 16000 185 16020
rect 245 16020 340 16060
rect 245 16000 315 16020
rect 30 15985 86 15991
rect 30 15925 34 15985
rect 115 15975 315 16000
rect 370 15991 400 16179
rect 344 15985 400 15991
rect 86 15925 344 15945
rect 396 15925 400 15985
rect 30 15915 400 15925
rect 430 16245 800 16255
rect 430 16185 434 16245
rect 486 16225 744 16245
rect 430 16179 486 16185
rect 430 15991 460 16179
rect 515 16170 715 16195
rect 796 16185 800 16245
rect 744 16179 800 16185
rect 515 16150 585 16170
rect 490 16110 585 16150
rect 645 16150 715 16170
rect 645 16110 740 16150
rect 490 16060 740 16110
rect 490 16020 585 16060
rect 515 16000 585 16020
rect 645 16020 740 16060
rect 645 16000 715 16020
rect 430 15985 486 15991
rect 430 15925 434 15985
rect 515 15975 715 16000
rect 770 15991 800 16179
rect 744 15985 800 15991
rect 486 15925 744 15945
rect 796 15925 800 15985
rect 430 15915 800 15925
rect 830 16245 1200 16255
rect 830 16185 834 16245
rect 886 16225 1144 16245
rect 830 16179 886 16185
rect 830 15991 860 16179
rect 915 16170 1115 16195
rect 1196 16185 1200 16245
rect 1144 16179 1200 16185
rect 915 16150 985 16170
rect 890 16110 985 16150
rect 1045 16150 1115 16170
rect 1045 16110 1140 16150
rect 890 16060 1140 16110
rect 890 16020 985 16060
rect 915 16000 985 16020
rect 1045 16020 1140 16060
rect 1045 16000 1115 16020
rect 830 15985 886 15991
rect 830 15925 834 15985
rect 915 15975 1115 16000
rect 1170 15991 1200 16179
rect 1144 15985 1200 15991
rect 886 15925 1144 15945
rect 1196 15925 1200 15985
rect 830 15915 1200 15925
rect 1230 16245 1600 16255
rect 1230 16185 1234 16245
rect 1286 16225 1544 16245
rect 1230 16179 1286 16185
rect 1230 15991 1260 16179
rect 1315 16170 1515 16195
rect 1596 16185 1600 16245
rect 1544 16179 1600 16185
rect 1315 16150 1385 16170
rect 1290 16110 1385 16150
rect 1445 16150 1515 16170
rect 1445 16110 1540 16150
rect 1290 16060 1540 16110
rect 1290 16020 1385 16060
rect 1315 16000 1385 16020
rect 1445 16020 1540 16060
rect 1445 16000 1515 16020
rect 1230 15985 1286 15991
rect 1230 15925 1234 15985
rect 1315 15975 1515 16000
rect 1570 15991 1600 16179
rect 1544 15985 1600 15991
rect 1286 15925 1544 15945
rect 1596 15925 1600 15985
rect 1230 15915 1600 15925
rect 1630 16245 2000 16255
rect 1630 16185 1634 16245
rect 1686 16225 1944 16245
rect 1630 16179 1686 16185
rect 1630 15991 1660 16179
rect 1715 16170 1915 16195
rect 1996 16185 2000 16245
rect 1944 16179 2000 16185
rect 1715 16150 1785 16170
rect 1690 16110 1785 16150
rect 1845 16150 1915 16170
rect 1845 16110 1940 16150
rect 1690 16060 1940 16110
rect 1690 16020 1785 16060
rect 1715 16000 1785 16020
rect 1845 16020 1940 16060
rect 1845 16000 1915 16020
rect 1630 15985 1686 15991
rect 1630 15925 1634 15985
rect 1715 15975 1915 16000
rect 1970 15991 2000 16179
rect 1944 15985 2000 15991
rect 1686 15925 1944 15945
rect 1996 15925 2000 15985
rect 1630 15915 2000 15925
rect 2030 16245 2400 16255
rect 2030 16185 2034 16245
rect 2086 16225 2344 16245
rect 2030 16179 2086 16185
rect 2030 15991 2060 16179
rect 2115 16170 2315 16195
rect 2396 16185 2400 16245
rect 2344 16179 2400 16185
rect 2115 16150 2185 16170
rect 2090 16110 2185 16150
rect 2245 16150 2315 16170
rect 2245 16110 2340 16150
rect 2090 16060 2340 16110
rect 2090 16020 2185 16060
rect 2115 16000 2185 16020
rect 2245 16020 2340 16060
rect 2245 16000 2315 16020
rect 2030 15985 2086 15991
rect 2030 15925 2034 15985
rect 2115 15975 2315 16000
rect 2370 15991 2400 16179
rect 2344 15985 2400 15991
rect 2086 15925 2344 15945
rect 2396 15925 2400 15985
rect 2030 15915 2400 15925
rect 2430 16245 2800 16255
rect 2430 16185 2434 16245
rect 2486 16225 2744 16245
rect 2430 16179 2486 16185
rect 2430 15991 2460 16179
rect 2515 16170 2715 16195
rect 2796 16185 2800 16245
rect 2744 16179 2800 16185
rect 2515 16150 2585 16170
rect 2490 16110 2585 16150
rect 2645 16150 2715 16170
rect 2645 16110 2740 16150
rect 2490 16060 2740 16110
rect 2490 16020 2585 16060
rect 2515 16000 2585 16020
rect 2645 16020 2740 16060
rect 2645 16000 2715 16020
rect 2430 15985 2486 15991
rect 2430 15925 2434 15985
rect 2515 15975 2715 16000
rect 2770 15991 2800 16179
rect 2744 15985 2800 15991
rect 2486 15925 2744 15945
rect 2796 15925 2800 15985
rect 2430 15915 2800 15925
rect 2830 16245 3200 16255
rect 2830 16185 2834 16245
rect 2886 16225 3144 16245
rect 2830 16179 2886 16185
rect 2830 15991 2860 16179
rect 2915 16170 3115 16195
rect 3196 16185 3200 16245
rect 3144 16179 3200 16185
rect 2915 16150 2985 16170
rect 2890 16110 2985 16150
rect 3045 16150 3115 16170
rect 3045 16110 3140 16150
rect 2890 16060 3140 16110
rect 2890 16020 2985 16060
rect 2915 16000 2985 16020
rect 3045 16020 3140 16060
rect 3045 16000 3115 16020
rect 2830 15985 2886 15991
rect 2830 15925 2834 15985
rect 2915 15975 3115 16000
rect 3170 15991 3200 16179
rect 3144 15985 3200 15991
rect 2886 15925 3144 15945
rect 3196 15925 3200 15985
rect 2830 15915 3200 15925
rect 3230 16245 3600 16255
rect 3230 16185 3234 16245
rect 3286 16225 3544 16245
rect 3230 16179 3286 16185
rect 3230 15991 3260 16179
rect 3315 16170 3515 16195
rect 3596 16185 3600 16245
rect 3544 16179 3600 16185
rect 3315 16150 3385 16170
rect 3290 16110 3385 16150
rect 3445 16150 3515 16170
rect 3445 16110 3540 16150
rect 3290 16060 3540 16110
rect 3290 16020 3385 16060
rect 3315 16000 3385 16020
rect 3445 16020 3540 16060
rect 3445 16000 3515 16020
rect 3230 15985 3286 15991
rect 3230 15925 3234 15985
rect 3315 15975 3515 16000
rect 3570 15991 3600 16179
rect 3544 15985 3600 15991
rect 3286 15925 3544 15945
rect 3596 15925 3600 15985
rect 3230 15915 3600 15925
rect 3630 16245 4000 16255
rect 3630 16185 3634 16245
rect 3686 16225 3944 16245
rect 3630 16179 3686 16185
rect 3630 15991 3660 16179
rect 3715 16170 3915 16195
rect 3996 16185 4000 16245
rect 3944 16179 4000 16185
rect 3715 16150 3785 16170
rect 3690 16110 3785 16150
rect 3845 16150 3915 16170
rect 3845 16110 3940 16150
rect 3690 16060 3940 16110
rect 3690 16020 3785 16060
rect 3715 16000 3785 16020
rect 3845 16020 3940 16060
rect 3845 16000 3915 16020
rect 3630 15985 3686 15991
rect 3630 15925 3634 15985
rect 3715 15975 3915 16000
rect 3970 15991 4000 16179
rect 3944 15985 4000 15991
rect 3686 15925 3944 15945
rect 3996 15925 4000 15985
rect 3630 15915 4000 15925
rect 4030 16245 4400 16255
rect 4030 16185 4034 16245
rect 4086 16225 4344 16245
rect 4030 16179 4086 16185
rect 4030 15991 4060 16179
rect 4115 16170 4315 16195
rect 4396 16185 4400 16245
rect 4344 16179 4400 16185
rect 4115 16150 4185 16170
rect 4090 16110 4185 16150
rect 4245 16150 4315 16170
rect 4245 16110 4340 16150
rect 4090 16060 4340 16110
rect 4090 16020 4185 16060
rect 4115 16000 4185 16020
rect 4245 16020 4340 16060
rect 4245 16000 4315 16020
rect 4030 15985 4086 15991
rect 4030 15925 4034 15985
rect 4115 15975 4315 16000
rect 4370 15991 4400 16179
rect 4344 15985 4400 15991
rect 4086 15925 4344 15945
rect 4396 15925 4400 15985
rect 4030 15915 4400 15925
rect 4430 16245 4800 16255
rect 4430 16185 4434 16245
rect 4486 16225 4744 16245
rect 4430 16179 4486 16185
rect 4430 15991 4460 16179
rect 4515 16170 4715 16195
rect 4796 16185 4800 16245
rect 4744 16179 4800 16185
rect 4515 16150 4585 16170
rect 4490 16110 4585 16150
rect 4645 16150 4715 16170
rect 4645 16110 4740 16150
rect 4490 16060 4740 16110
rect 4490 16020 4585 16060
rect 4515 16000 4585 16020
rect 4645 16020 4740 16060
rect 4645 16000 4715 16020
rect 4430 15985 4486 15991
rect 4430 15925 4434 15985
rect 4515 15975 4715 16000
rect 4770 15991 4800 16179
rect 4744 15985 4800 15991
rect 4486 15925 4744 15945
rect 4796 15925 4800 15985
rect 4430 15915 4800 15925
rect 4830 16245 5200 16255
rect 4830 16185 4834 16245
rect 4886 16225 5144 16245
rect 4830 16179 4886 16185
rect 4830 15991 4860 16179
rect 4915 16170 5115 16195
rect 5196 16185 5200 16245
rect 5144 16179 5200 16185
rect 4915 16150 4985 16170
rect 4890 16110 4985 16150
rect 5045 16150 5115 16170
rect 5045 16110 5140 16150
rect 4890 16060 5140 16110
rect 4890 16020 4985 16060
rect 4915 16000 4985 16020
rect 5045 16020 5140 16060
rect 5045 16000 5115 16020
rect 4830 15985 4886 15991
rect 4830 15925 4834 15985
rect 4915 15975 5115 16000
rect 5170 15991 5200 16179
rect 5144 15985 5200 15991
rect 4886 15925 5144 15945
rect 5196 15925 5200 15985
rect 4830 15915 5200 15925
rect 5230 16245 5600 16255
rect 5230 16185 5234 16245
rect 5286 16225 5544 16245
rect 5230 16179 5286 16185
rect 5230 15991 5260 16179
rect 5315 16170 5515 16195
rect 5596 16185 5600 16245
rect 5544 16179 5600 16185
rect 5315 16150 5385 16170
rect 5290 16110 5385 16150
rect 5445 16150 5515 16170
rect 5445 16110 5540 16150
rect 5290 16060 5540 16110
rect 5290 16020 5385 16060
rect 5315 16000 5385 16020
rect 5445 16020 5540 16060
rect 5445 16000 5515 16020
rect 5230 15985 5286 15991
rect 5230 15925 5234 15985
rect 5315 15975 5515 16000
rect 5570 15991 5600 16179
rect 5544 15985 5600 15991
rect 5286 15925 5544 15945
rect 5596 15925 5600 15985
rect 5230 15915 5600 15925
rect 5630 16245 6000 16255
rect 5630 16185 5634 16245
rect 5686 16225 5944 16245
rect 5630 16179 5686 16185
rect 5630 15991 5660 16179
rect 5715 16170 5915 16195
rect 5996 16185 6000 16245
rect 5944 16179 6000 16185
rect 5715 16150 5785 16170
rect 5690 16110 5785 16150
rect 5845 16150 5915 16170
rect 5845 16110 5940 16150
rect 5690 16060 5940 16110
rect 5690 16020 5785 16060
rect 5715 16000 5785 16020
rect 5845 16020 5940 16060
rect 5845 16000 5915 16020
rect 5630 15985 5686 15991
rect 5630 15925 5634 15985
rect 5715 15975 5915 16000
rect 5970 15991 6000 16179
rect 5944 15985 6000 15991
rect 5686 15925 5944 15945
rect 5996 15925 6000 15985
rect 5630 15915 6000 15925
rect 6030 16245 6400 16255
rect 6030 16185 6034 16245
rect 6086 16225 6344 16245
rect 6030 16179 6086 16185
rect 6030 15991 6060 16179
rect 6115 16170 6315 16195
rect 6396 16185 6400 16245
rect 6344 16179 6400 16185
rect 6115 16150 6185 16170
rect 6090 16110 6185 16150
rect 6245 16150 6315 16170
rect 6245 16110 6340 16150
rect 6090 16060 6340 16110
rect 6090 16020 6185 16060
rect 6115 16000 6185 16020
rect 6245 16020 6340 16060
rect 6245 16000 6315 16020
rect 6030 15985 6086 15991
rect 6030 15925 6034 15985
rect 6115 15975 6315 16000
rect 6370 15991 6400 16179
rect 6344 15985 6400 15991
rect 6086 15925 6344 15945
rect 6396 15925 6400 15985
rect 6030 15915 6400 15925
rect 6430 16245 6800 16255
rect 6430 16185 6434 16245
rect 6486 16225 6744 16245
rect 6430 16179 6486 16185
rect 6430 15991 6460 16179
rect 6515 16170 6715 16195
rect 6796 16185 6800 16245
rect 6744 16179 6800 16185
rect 6515 16150 6585 16170
rect 6490 16110 6585 16150
rect 6645 16150 6715 16170
rect 6645 16110 6740 16150
rect 6490 16060 6740 16110
rect 6490 16020 6585 16060
rect 6515 16000 6585 16020
rect 6645 16020 6740 16060
rect 6645 16000 6715 16020
rect 6430 15985 6486 15991
rect 6430 15925 6434 15985
rect 6515 15975 6715 16000
rect 6770 15991 6800 16179
rect 6744 15985 6800 15991
rect 6486 15925 6744 15945
rect 6796 15925 6800 15985
rect 6430 15915 6800 15925
rect 6830 16245 7200 16255
rect 6830 16185 6834 16245
rect 6886 16225 7144 16245
rect 6830 16179 6886 16185
rect 6830 15991 6860 16179
rect 6915 16170 7115 16195
rect 7196 16185 7200 16245
rect 7144 16179 7200 16185
rect 6915 16150 6985 16170
rect 6890 16110 6985 16150
rect 7045 16150 7115 16170
rect 7045 16110 7140 16150
rect 6890 16060 7140 16110
rect 6890 16020 6985 16060
rect 6915 16000 6985 16020
rect 7045 16020 7140 16060
rect 7045 16000 7115 16020
rect 6830 15985 6886 15991
rect 6830 15925 6834 15985
rect 6915 15975 7115 16000
rect 7170 15991 7200 16179
rect 7144 15985 7200 15991
rect 6886 15925 7144 15945
rect 7196 15925 7200 15985
rect 6830 15915 7200 15925
rect 7230 16245 7600 16255
rect 7230 16185 7234 16245
rect 7286 16225 7544 16245
rect 7230 16179 7286 16185
rect 7230 15991 7260 16179
rect 7315 16170 7515 16195
rect 7596 16185 7600 16245
rect 7544 16179 7600 16185
rect 7315 16150 7385 16170
rect 7290 16110 7385 16150
rect 7445 16150 7515 16170
rect 7445 16110 7540 16150
rect 7290 16060 7540 16110
rect 7290 16020 7385 16060
rect 7315 16000 7385 16020
rect 7445 16020 7540 16060
rect 7445 16000 7515 16020
rect 7230 15985 7286 15991
rect 7230 15925 7234 15985
rect 7315 15975 7515 16000
rect 7570 15991 7600 16179
rect 7544 15985 7600 15991
rect 7286 15925 7544 15945
rect 7596 15925 7600 15985
rect 7230 15915 7600 15925
rect 7630 16245 8000 16255
rect 7630 16185 7634 16245
rect 7686 16225 7944 16245
rect 7630 16179 7686 16185
rect 7630 15991 7660 16179
rect 7715 16170 7915 16195
rect 7996 16185 8000 16245
rect 7944 16179 8000 16185
rect 7715 16150 7785 16170
rect 7690 16110 7785 16150
rect 7845 16150 7915 16170
rect 7845 16110 7940 16150
rect 7690 16060 7940 16110
rect 7690 16020 7785 16060
rect 7715 16000 7785 16020
rect 7845 16020 7940 16060
rect 7845 16000 7915 16020
rect 7630 15985 7686 15991
rect 7630 15925 7634 15985
rect 7715 15975 7915 16000
rect 7970 15991 8000 16179
rect 7944 15985 8000 15991
rect 7686 15925 7944 15945
rect 7996 15925 8000 15985
rect 7630 15915 8000 15925
rect 8030 16245 8400 16255
rect 8030 16185 8034 16245
rect 8086 16225 8344 16245
rect 8030 16179 8086 16185
rect 8030 15991 8060 16179
rect 8115 16170 8315 16195
rect 8396 16185 8400 16245
rect 8344 16179 8400 16185
rect 8115 16150 8185 16170
rect 8090 16110 8185 16150
rect 8245 16150 8315 16170
rect 8245 16110 8340 16150
rect 8090 16060 8340 16110
rect 8090 16020 8185 16060
rect 8115 16000 8185 16020
rect 8245 16020 8340 16060
rect 8245 16000 8315 16020
rect 8030 15985 8086 15991
rect 8030 15925 8034 15985
rect 8115 15975 8315 16000
rect 8370 15991 8400 16179
rect 8344 15985 8400 15991
rect 8086 15925 8344 15945
rect 8396 15925 8400 15985
rect 8030 15915 8400 15925
rect 8430 16245 8800 16255
rect 8430 16185 8434 16245
rect 8486 16225 8744 16245
rect 8430 16179 8486 16185
rect 8430 15991 8460 16179
rect 8515 16170 8715 16195
rect 8796 16185 8800 16245
rect 8744 16179 8800 16185
rect 8515 16150 8585 16170
rect 8490 16110 8585 16150
rect 8645 16150 8715 16170
rect 8645 16110 8740 16150
rect 8490 16060 8740 16110
rect 8490 16020 8585 16060
rect 8515 16000 8585 16020
rect 8645 16020 8740 16060
rect 8645 16000 8715 16020
rect 8430 15985 8486 15991
rect 8430 15925 8434 15985
rect 8515 15975 8715 16000
rect 8770 15991 8800 16179
rect 8744 15985 8800 15991
rect 8486 15925 8744 15945
rect 8796 15925 8800 15985
rect 8430 15915 8800 15925
rect 8830 16245 9200 16255
rect 8830 16185 8834 16245
rect 8886 16225 9144 16245
rect 8830 16179 8886 16185
rect 8830 15991 8860 16179
rect 8915 16170 9115 16195
rect 9196 16185 9200 16245
rect 9144 16179 9200 16185
rect 8915 16150 8985 16170
rect 8890 16110 8985 16150
rect 9045 16150 9115 16170
rect 9045 16110 9140 16150
rect 8890 16060 9140 16110
rect 8890 16020 8985 16060
rect 8915 16000 8985 16020
rect 9045 16020 9140 16060
rect 9045 16000 9115 16020
rect 8830 15985 8886 15991
rect 8830 15925 8834 15985
rect 8915 15975 9115 16000
rect 9170 15991 9200 16179
rect 9144 15985 9200 15991
rect 8886 15925 9144 15945
rect 9196 15925 9200 15985
rect 8830 15915 9200 15925
rect 9230 16245 9600 16255
rect 9230 16185 9234 16245
rect 9286 16225 9544 16245
rect 9230 16179 9286 16185
rect 9230 15991 9260 16179
rect 9315 16170 9515 16195
rect 9596 16185 9600 16245
rect 9544 16179 9600 16185
rect 9315 16150 9385 16170
rect 9290 16110 9385 16150
rect 9445 16150 9515 16170
rect 9445 16110 9540 16150
rect 9290 16060 9540 16110
rect 9290 16020 9385 16060
rect 9315 16000 9385 16020
rect 9445 16020 9540 16060
rect 9445 16000 9515 16020
rect 9230 15985 9286 15991
rect 9230 15925 9234 15985
rect 9315 15975 9515 16000
rect 9570 15991 9600 16179
rect 9544 15985 9600 15991
rect 9286 15925 9544 15945
rect 9596 15925 9600 15985
rect 9230 15915 9600 15925
rect 9630 16245 10000 16255
rect 9630 16185 9634 16245
rect 9686 16225 9944 16245
rect 9630 16179 9686 16185
rect 9630 15991 9660 16179
rect 9715 16170 9915 16195
rect 9996 16185 10000 16245
rect 9944 16179 10000 16185
rect 9715 16150 9785 16170
rect 9690 16110 9785 16150
rect 9845 16150 9915 16170
rect 9845 16110 9940 16150
rect 9690 16060 9940 16110
rect 9690 16020 9785 16060
rect 9715 16000 9785 16020
rect 9845 16020 9940 16060
rect 9845 16000 9915 16020
rect 9630 15985 9686 15991
rect 9630 15925 9634 15985
rect 9715 15975 9915 16000
rect 9970 15991 10000 16179
rect 9944 15985 10000 15991
rect 9686 15925 9944 15945
rect 9996 15925 10000 15985
rect 9630 15915 10000 15925
rect 10030 16245 10400 16255
rect 10030 16185 10034 16245
rect 10086 16225 10344 16245
rect 10030 16179 10086 16185
rect 10030 15991 10060 16179
rect 10115 16170 10315 16195
rect 10396 16185 10400 16245
rect 10344 16179 10400 16185
rect 10115 16150 10185 16170
rect 10090 16110 10185 16150
rect 10245 16150 10315 16170
rect 10245 16110 10340 16150
rect 10090 16060 10340 16110
rect 10090 16020 10185 16060
rect 10115 16000 10185 16020
rect 10245 16020 10340 16060
rect 10245 16000 10315 16020
rect 10030 15985 10086 15991
rect 10030 15925 10034 15985
rect 10115 15975 10315 16000
rect 10370 15991 10400 16179
rect 10344 15985 10400 15991
rect 10086 15925 10344 15945
rect 10396 15925 10400 15985
rect 10030 15915 10400 15925
rect 10430 16245 10800 16255
rect 10430 16185 10434 16245
rect 10486 16225 10744 16245
rect 10430 16179 10486 16185
rect 10430 15991 10460 16179
rect 10515 16170 10715 16195
rect 10796 16185 10800 16245
rect 10744 16179 10800 16185
rect 10515 16150 10585 16170
rect 10490 16110 10585 16150
rect 10645 16150 10715 16170
rect 10645 16110 10740 16150
rect 10490 16060 10740 16110
rect 10490 16020 10585 16060
rect 10515 16000 10585 16020
rect 10645 16020 10740 16060
rect 10645 16000 10715 16020
rect 10430 15985 10486 15991
rect 10430 15925 10434 15985
rect 10515 15975 10715 16000
rect 10770 15991 10800 16179
rect 10744 15985 10800 15991
rect 10486 15925 10744 15945
rect 10796 15925 10800 15985
rect 10430 15915 10800 15925
rect 10830 16245 11200 16255
rect 10830 16185 10834 16245
rect 10886 16225 11144 16245
rect 10830 16179 10886 16185
rect 10830 15991 10860 16179
rect 10915 16170 11115 16195
rect 11196 16185 11200 16245
rect 11144 16179 11200 16185
rect 10915 16150 10985 16170
rect 10890 16110 10985 16150
rect 11045 16150 11115 16170
rect 11045 16110 11140 16150
rect 10890 16060 11140 16110
rect 10890 16020 10985 16060
rect 10915 16000 10985 16020
rect 11045 16020 11140 16060
rect 11045 16000 11115 16020
rect 10830 15985 10886 15991
rect 10830 15925 10834 15985
rect 10915 15975 11115 16000
rect 11170 15991 11200 16179
rect 11144 15985 11200 15991
rect 10886 15925 11144 15945
rect 11196 15925 11200 15985
rect 10830 15915 11200 15925
rect 11230 16245 11600 16255
rect 11230 16185 11234 16245
rect 11286 16225 11544 16245
rect 11230 16179 11286 16185
rect 11230 15991 11260 16179
rect 11315 16170 11515 16195
rect 11596 16185 11600 16245
rect 11544 16179 11600 16185
rect 11315 16150 11385 16170
rect 11290 16110 11385 16150
rect 11445 16150 11515 16170
rect 11445 16110 11540 16150
rect 11290 16060 11540 16110
rect 11290 16020 11385 16060
rect 11315 16000 11385 16020
rect 11445 16020 11540 16060
rect 11445 16000 11515 16020
rect 11230 15985 11286 15991
rect 11230 15925 11234 15985
rect 11315 15975 11515 16000
rect 11570 15991 11600 16179
rect 11544 15985 11600 15991
rect 11286 15925 11544 15945
rect 11596 15925 11600 15985
rect 11230 15915 11600 15925
rect 11630 16245 12000 16255
rect 11630 16185 11634 16245
rect 11686 16225 11944 16245
rect 11630 16179 11686 16185
rect 11630 15991 11660 16179
rect 11715 16170 11915 16195
rect 11996 16185 12000 16245
rect 11944 16179 12000 16185
rect 11715 16150 11785 16170
rect 11690 16110 11785 16150
rect 11845 16150 11915 16170
rect 11845 16110 11940 16150
rect 11690 16060 11940 16110
rect 11690 16020 11785 16060
rect 11715 16000 11785 16020
rect 11845 16020 11940 16060
rect 11845 16000 11915 16020
rect 11630 15985 11686 15991
rect 11630 15925 11634 15985
rect 11715 15975 11915 16000
rect 11970 15991 12000 16179
rect 11944 15985 12000 15991
rect 11686 15925 11944 15945
rect 11996 15925 12000 15985
rect 11630 15915 12000 15925
rect 12030 16245 12400 16255
rect 12030 16185 12034 16245
rect 12086 16225 12344 16245
rect 12030 16179 12086 16185
rect 12030 15991 12060 16179
rect 12115 16170 12315 16195
rect 12396 16185 12400 16245
rect 12344 16179 12400 16185
rect 12115 16150 12185 16170
rect 12090 16110 12185 16150
rect 12245 16150 12315 16170
rect 12245 16110 12340 16150
rect 12090 16060 12340 16110
rect 12090 16020 12185 16060
rect 12115 16000 12185 16020
rect 12245 16020 12340 16060
rect 12245 16000 12315 16020
rect 12030 15985 12086 15991
rect 12030 15925 12034 15985
rect 12115 15975 12315 16000
rect 12370 15991 12400 16179
rect 12344 15985 12400 15991
rect 12086 15925 12344 15945
rect 12396 15925 12400 15985
rect 12030 15915 12400 15925
rect 12430 16245 12800 16255
rect 12430 16185 12434 16245
rect 12486 16225 12744 16245
rect 12430 16179 12486 16185
rect 12430 15991 12460 16179
rect 12515 16170 12715 16195
rect 12796 16185 12800 16245
rect 12744 16179 12800 16185
rect 12515 16150 12585 16170
rect 12490 16110 12585 16150
rect 12645 16150 12715 16170
rect 12645 16110 12740 16150
rect 12490 16060 12740 16110
rect 12490 16020 12585 16060
rect 12515 16000 12585 16020
rect 12645 16020 12740 16060
rect 12645 16000 12715 16020
rect 12430 15985 12486 15991
rect 12430 15925 12434 15985
rect 12515 15975 12715 16000
rect 12770 15991 12800 16179
rect 12744 15985 12800 15991
rect 12486 15925 12744 15945
rect 12796 15925 12800 15985
rect 12430 15915 12800 15925
rect 12830 16245 13200 16255
rect 12830 16185 12834 16245
rect 12886 16225 13144 16245
rect 12830 16179 12886 16185
rect 12830 15991 12860 16179
rect 12915 16170 13115 16195
rect 13196 16185 13200 16245
rect 13144 16179 13200 16185
rect 12915 16150 12985 16170
rect 12890 16110 12985 16150
rect 13045 16150 13115 16170
rect 13045 16110 13140 16150
rect 12890 16060 13140 16110
rect 12890 16020 12985 16060
rect 12915 16000 12985 16020
rect 13045 16020 13140 16060
rect 13045 16000 13115 16020
rect 12830 15985 12886 15991
rect 12830 15925 12834 15985
rect 12915 15975 13115 16000
rect 13170 15991 13200 16179
rect 13144 15985 13200 15991
rect 12886 15925 13144 15945
rect 13196 15925 13200 15985
rect 12830 15915 13200 15925
rect -370 15875 0 15885
rect -370 15815 -366 15875
rect -314 15855 -56 15875
rect -370 15809 -314 15815
rect -370 15621 -340 15809
rect -285 15800 -85 15825
rect -4 15815 0 15875
rect -56 15809 0 15815
rect -285 15780 -215 15800
rect -310 15740 -215 15780
rect -155 15780 -85 15800
rect -155 15740 -60 15780
rect -310 15690 -60 15740
rect -310 15650 -215 15690
rect -285 15630 -215 15650
rect -155 15650 -60 15690
rect -155 15630 -85 15650
rect -370 15615 -314 15621
rect -370 15555 -366 15615
rect -285 15605 -85 15630
rect -30 15621 0 15809
rect -56 15615 0 15621
rect -314 15555 -56 15575
rect -4 15555 0 15615
rect -370 15545 0 15555
rect 30 15875 400 15885
rect 30 15815 34 15875
rect 86 15855 344 15875
rect 30 15809 86 15815
rect 30 15621 60 15809
rect 115 15800 315 15825
rect 396 15815 400 15875
rect 344 15809 400 15815
rect 115 15780 185 15800
rect 90 15740 185 15780
rect 245 15780 315 15800
rect 245 15740 340 15780
rect 90 15690 340 15740
rect 90 15650 185 15690
rect 115 15630 185 15650
rect 245 15650 340 15690
rect 245 15630 315 15650
rect 30 15615 86 15621
rect 30 15555 34 15615
rect 115 15605 315 15630
rect 370 15621 400 15809
rect 344 15615 400 15621
rect 86 15555 344 15575
rect 396 15555 400 15615
rect 30 15545 400 15555
rect 430 15875 800 15885
rect 430 15815 434 15875
rect 486 15855 744 15875
rect 430 15809 486 15815
rect 430 15621 460 15809
rect 515 15800 715 15825
rect 796 15815 800 15875
rect 744 15809 800 15815
rect 515 15780 585 15800
rect 490 15740 585 15780
rect 645 15780 715 15800
rect 645 15740 740 15780
rect 490 15690 740 15740
rect 490 15650 585 15690
rect 515 15630 585 15650
rect 645 15650 740 15690
rect 645 15630 715 15650
rect 430 15615 486 15621
rect 430 15555 434 15615
rect 515 15605 715 15630
rect 770 15621 800 15809
rect 744 15615 800 15621
rect 486 15555 744 15575
rect 796 15555 800 15615
rect 430 15545 800 15555
rect 830 15875 1200 15885
rect 830 15815 834 15875
rect 886 15855 1144 15875
rect 830 15809 886 15815
rect 830 15621 860 15809
rect 915 15800 1115 15825
rect 1196 15815 1200 15875
rect 1144 15809 1200 15815
rect 915 15780 985 15800
rect 890 15740 985 15780
rect 1045 15780 1115 15800
rect 1045 15740 1140 15780
rect 890 15690 1140 15740
rect 890 15650 985 15690
rect 915 15630 985 15650
rect 1045 15650 1140 15690
rect 1045 15630 1115 15650
rect 830 15615 886 15621
rect 830 15555 834 15615
rect 915 15605 1115 15630
rect 1170 15621 1200 15809
rect 1144 15615 1200 15621
rect 886 15555 1144 15575
rect 1196 15555 1200 15615
rect 830 15545 1200 15555
rect 1230 15875 1600 15885
rect 1230 15815 1234 15875
rect 1286 15855 1544 15875
rect 1230 15809 1286 15815
rect 1230 15621 1260 15809
rect 1315 15800 1515 15825
rect 1596 15815 1600 15875
rect 1544 15809 1600 15815
rect 1315 15780 1385 15800
rect 1290 15740 1385 15780
rect 1445 15780 1515 15800
rect 1445 15740 1540 15780
rect 1290 15690 1540 15740
rect 1290 15650 1385 15690
rect 1315 15630 1385 15650
rect 1445 15650 1540 15690
rect 1445 15630 1515 15650
rect 1230 15615 1286 15621
rect 1230 15555 1234 15615
rect 1315 15605 1515 15630
rect 1570 15621 1600 15809
rect 1544 15615 1600 15621
rect 1286 15555 1544 15575
rect 1596 15555 1600 15615
rect 1230 15545 1600 15555
rect 1630 15875 2000 15885
rect 1630 15815 1634 15875
rect 1686 15855 1944 15875
rect 1630 15809 1686 15815
rect 1630 15621 1660 15809
rect 1715 15800 1915 15825
rect 1996 15815 2000 15875
rect 1944 15809 2000 15815
rect 1715 15780 1785 15800
rect 1690 15740 1785 15780
rect 1845 15780 1915 15800
rect 1845 15740 1940 15780
rect 1690 15690 1940 15740
rect 1690 15650 1785 15690
rect 1715 15630 1785 15650
rect 1845 15650 1940 15690
rect 1845 15630 1915 15650
rect 1630 15615 1686 15621
rect 1630 15555 1634 15615
rect 1715 15605 1915 15630
rect 1970 15621 2000 15809
rect 1944 15615 2000 15621
rect 1686 15555 1944 15575
rect 1996 15555 2000 15615
rect 1630 15545 2000 15555
rect 2030 15875 2400 15885
rect 2030 15815 2034 15875
rect 2086 15855 2344 15875
rect 2030 15809 2086 15815
rect 2030 15621 2060 15809
rect 2115 15800 2315 15825
rect 2396 15815 2400 15875
rect 2344 15809 2400 15815
rect 2115 15780 2185 15800
rect 2090 15740 2185 15780
rect 2245 15780 2315 15800
rect 2245 15740 2340 15780
rect 2090 15690 2340 15740
rect 2090 15650 2185 15690
rect 2115 15630 2185 15650
rect 2245 15650 2340 15690
rect 2245 15630 2315 15650
rect 2030 15615 2086 15621
rect 2030 15555 2034 15615
rect 2115 15605 2315 15630
rect 2370 15621 2400 15809
rect 2344 15615 2400 15621
rect 2086 15555 2344 15575
rect 2396 15555 2400 15615
rect 2030 15545 2400 15555
rect 2430 15875 2800 15885
rect 2430 15815 2434 15875
rect 2486 15855 2744 15875
rect 2430 15809 2486 15815
rect 2430 15621 2460 15809
rect 2515 15800 2715 15825
rect 2796 15815 2800 15875
rect 2744 15809 2800 15815
rect 2515 15780 2585 15800
rect 2490 15740 2585 15780
rect 2645 15780 2715 15800
rect 2645 15740 2740 15780
rect 2490 15690 2740 15740
rect 2490 15650 2585 15690
rect 2515 15630 2585 15650
rect 2645 15650 2740 15690
rect 2645 15630 2715 15650
rect 2430 15615 2486 15621
rect 2430 15555 2434 15615
rect 2515 15605 2715 15630
rect 2770 15621 2800 15809
rect 2744 15615 2800 15621
rect 2486 15555 2744 15575
rect 2796 15555 2800 15615
rect 2430 15545 2800 15555
rect 2830 15875 3200 15885
rect 2830 15815 2834 15875
rect 2886 15855 3144 15875
rect 2830 15809 2886 15815
rect 2830 15621 2860 15809
rect 2915 15800 3115 15825
rect 3196 15815 3200 15875
rect 3144 15809 3200 15815
rect 2915 15780 2985 15800
rect 2890 15740 2985 15780
rect 3045 15780 3115 15800
rect 3045 15740 3140 15780
rect 2890 15690 3140 15740
rect 2890 15650 2985 15690
rect 2915 15630 2985 15650
rect 3045 15650 3140 15690
rect 3045 15630 3115 15650
rect 2830 15615 2886 15621
rect 2830 15555 2834 15615
rect 2915 15605 3115 15630
rect 3170 15621 3200 15809
rect 3144 15615 3200 15621
rect 2886 15555 3144 15575
rect 3196 15555 3200 15615
rect 2830 15545 3200 15555
rect 3230 15875 3600 15885
rect 3230 15815 3234 15875
rect 3286 15855 3544 15875
rect 3230 15809 3286 15815
rect 3230 15621 3260 15809
rect 3315 15800 3515 15825
rect 3596 15815 3600 15875
rect 3544 15809 3600 15815
rect 3315 15780 3385 15800
rect 3290 15740 3385 15780
rect 3445 15780 3515 15800
rect 3445 15740 3540 15780
rect 3290 15690 3540 15740
rect 3290 15650 3385 15690
rect 3315 15630 3385 15650
rect 3445 15650 3540 15690
rect 3445 15630 3515 15650
rect 3230 15615 3286 15621
rect 3230 15555 3234 15615
rect 3315 15605 3515 15630
rect 3570 15621 3600 15809
rect 3544 15615 3600 15621
rect 3286 15555 3544 15575
rect 3596 15555 3600 15615
rect 3230 15545 3600 15555
rect 3630 15875 4000 15885
rect 3630 15815 3634 15875
rect 3686 15855 3944 15875
rect 3630 15809 3686 15815
rect 3630 15621 3660 15809
rect 3715 15800 3915 15825
rect 3996 15815 4000 15875
rect 3944 15809 4000 15815
rect 3715 15780 3785 15800
rect 3690 15740 3785 15780
rect 3845 15780 3915 15800
rect 3845 15740 3940 15780
rect 3690 15690 3940 15740
rect 3690 15650 3785 15690
rect 3715 15630 3785 15650
rect 3845 15650 3940 15690
rect 3845 15630 3915 15650
rect 3630 15615 3686 15621
rect 3630 15555 3634 15615
rect 3715 15605 3915 15630
rect 3970 15621 4000 15809
rect 3944 15615 4000 15621
rect 3686 15555 3944 15575
rect 3996 15555 4000 15615
rect 3630 15545 4000 15555
rect 4030 15875 4400 15885
rect 4030 15815 4034 15875
rect 4086 15855 4344 15875
rect 4030 15809 4086 15815
rect 4030 15621 4060 15809
rect 4115 15800 4315 15825
rect 4396 15815 4400 15875
rect 4344 15809 4400 15815
rect 4115 15780 4185 15800
rect 4090 15740 4185 15780
rect 4245 15780 4315 15800
rect 4245 15740 4340 15780
rect 4090 15690 4340 15740
rect 4090 15650 4185 15690
rect 4115 15630 4185 15650
rect 4245 15650 4340 15690
rect 4245 15630 4315 15650
rect 4030 15615 4086 15621
rect 4030 15555 4034 15615
rect 4115 15605 4315 15630
rect 4370 15621 4400 15809
rect 4344 15615 4400 15621
rect 4086 15555 4344 15575
rect 4396 15555 4400 15615
rect 4030 15545 4400 15555
rect 4430 15875 4800 15885
rect 4430 15815 4434 15875
rect 4486 15855 4744 15875
rect 4430 15809 4486 15815
rect 4430 15621 4460 15809
rect 4515 15800 4715 15825
rect 4796 15815 4800 15875
rect 4744 15809 4800 15815
rect 4515 15780 4585 15800
rect 4490 15740 4585 15780
rect 4645 15780 4715 15800
rect 4645 15740 4740 15780
rect 4490 15690 4740 15740
rect 4490 15650 4585 15690
rect 4515 15630 4585 15650
rect 4645 15650 4740 15690
rect 4645 15630 4715 15650
rect 4430 15615 4486 15621
rect 4430 15555 4434 15615
rect 4515 15605 4715 15630
rect 4770 15621 4800 15809
rect 4744 15615 4800 15621
rect 4486 15555 4744 15575
rect 4796 15555 4800 15615
rect 4430 15545 4800 15555
rect 4830 15875 5200 15885
rect 4830 15815 4834 15875
rect 4886 15855 5144 15875
rect 4830 15809 4886 15815
rect 4830 15621 4860 15809
rect 4915 15800 5115 15825
rect 5196 15815 5200 15875
rect 5144 15809 5200 15815
rect 4915 15780 4985 15800
rect 4890 15740 4985 15780
rect 5045 15780 5115 15800
rect 5045 15740 5140 15780
rect 4890 15690 5140 15740
rect 4890 15650 4985 15690
rect 4915 15630 4985 15650
rect 5045 15650 5140 15690
rect 5045 15630 5115 15650
rect 4830 15615 4886 15621
rect 4830 15555 4834 15615
rect 4915 15605 5115 15630
rect 5170 15621 5200 15809
rect 5144 15615 5200 15621
rect 4886 15555 5144 15575
rect 5196 15555 5200 15615
rect 4830 15545 5200 15555
rect 5230 15875 5600 15885
rect 5230 15815 5234 15875
rect 5286 15855 5544 15875
rect 5230 15809 5286 15815
rect 5230 15621 5260 15809
rect 5315 15800 5515 15825
rect 5596 15815 5600 15875
rect 5544 15809 5600 15815
rect 5315 15780 5385 15800
rect 5290 15740 5385 15780
rect 5445 15780 5515 15800
rect 5445 15740 5540 15780
rect 5290 15690 5540 15740
rect 5290 15650 5385 15690
rect 5315 15630 5385 15650
rect 5445 15650 5540 15690
rect 5445 15630 5515 15650
rect 5230 15615 5286 15621
rect 5230 15555 5234 15615
rect 5315 15605 5515 15630
rect 5570 15621 5600 15809
rect 5544 15615 5600 15621
rect 5286 15555 5544 15575
rect 5596 15555 5600 15615
rect 5230 15545 5600 15555
rect 5630 15875 6000 15885
rect 5630 15815 5634 15875
rect 5686 15855 5944 15875
rect 5630 15809 5686 15815
rect 5630 15621 5660 15809
rect 5715 15800 5915 15825
rect 5996 15815 6000 15875
rect 5944 15809 6000 15815
rect 5715 15780 5785 15800
rect 5690 15740 5785 15780
rect 5845 15780 5915 15800
rect 5845 15740 5940 15780
rect 5690 15690 5940 15740
rect 5690 15650 5785 15690
rect 5715 15630 5785 15650
rect 5845 15650 5940 15690
rect 5845 15630 5915 15650
rect 5630 15615 5686 15621
rect 5630 15555 5634 15615
rect 5715 15605 5915 15630
rect 5970 15621 6000 15809
rect 5944 15615 6000 15621
rect 5686 15555 5944 15575
rect 5996 15555 6000 15615
rect 5630 15545 6000 15555
rect 6030 15875 6400 15885
rect 6030 15815 6034 15875
rect 6086 15855 6344 15875
rect 6030 15809 6086 15815
rect 6030 15621 6060 15809
rect 6115 15800 6315 15825
rect 6396 15815 6400 15875
rect 6344 15809 6400 15815
rect 6115 15780 6185 15800
rect 6090 15740 6185 15780
rect 6245 15780 6315 15800
rect 6245 15740 6340 15780
rect 6090 15690 6340 15740
rect 6090 15650 6185 15690
rect 6115 15630 6185 15650
rect 6245 15650 6340 15690
rect 6245 15630 6315 15650
rect 6030 15615 6086 15621
rect 6030 15555 6034 15615
rect 6115 15605 6315 15630
rect 6370 15621 6400 15809
rect 6344 15615 6400 15621
rect 6086 15555 6344 15575
rect 6396 15555 6400 15615
rect 6030 15545 6400 15555
rect 6430 15875 6800 15885
rect 6430 15815 6434 15875
rect 6486 15855 6744 15875
rect 6430 15809 6486 15815
rect 6430 15621 6460 15809
rect 6515 15800 6715 15825
rect 6796 15815 6800 15875
rect 6744 15809 6800 15815
rect 6515 15780 6585 15800
rect 6490 15740 6585 15780
rect 6645 15780 6715 15800
rect 6645 15740 6740 15780
rect 6490 15690 6740 15740
rect 6490 15650 6585 15690
rect 6515 15630 6585 15650
rect 6645 15650 6740 15690
rect 6645 15630 6715 15650
rect 6430 15615 6486 15621
rect 6430 15555 6434 15615
rect 6515 15605 6715 15630
rect 6770 15621 6800 15809
rect 6744 15615 6800 15621
rect 6486 15555 6744 15575
rect 6796 15555 6800 15615
rect 6430 15545 6800 15555
rect 6830 15875 7200 15885
rect 6830 15815 6834 15875
rect 6886 15855 7144 15875
rect 6830 15809 6886 15815
rect 6830 15621 6860 15809
rect 6915 15800 7115 15825
rect 7196 15815 7200 15875
rect 7144 15809 7200 15815
rect 6915 15780 6985 15800
rect 6890 15740 6985 15780
rect 7045 15780 7115 15800
rect 7045 15740 7140 15780
rect 6890 15690 7140 15740
rect 6890 15650 6985 15690
rect 6915 15630 6985 15650
rect 7045 15650 7140 15690
rect 7045 15630 7115 15650
rect 6830 15615 6886 15621
rect 6830 15555 6834 15615
rect 6915 15605 7115 15630
rect 7170 15621 7200 15809
rect 7144 15615 7200 15621
rect 6886 15555 7144 15575
rect 7196 15555 7200 15615
rect 6830 15545 7200 15555
rect 7230 15875 7600 15885
rect 7230 15815 7234 15875
rect 7286 15855 7544 15875
rect 7230 15809 7286 15815
rect 7230 15621 7260 15809
rect 7315 15800 7515 15825
rect 7596 15815 7600 15875
rect 7544 15809 7600 15815
rect 7315 15780 7385 15800
rect 7290 15740 7385 15780
rect 7445 15780 7515 15800
rect 7445 15740 7540 15780
rect 7290 15690 7540 15740
rect 7290 15650 7385 15690
rect 7315 15630 7385 15650
rect 7445 15650 7540 15690
rect 7445 15630 7515 15650
rect 7230 15615 7286 15621
rect 7230 15555 7234 15615
rect 7315 15605 7515 15630
rect 7570 15621 7600 15809
rect 7544 15615 7600 15621
rect 7286 15555 7544 15575
rect 7596 15555 7600 15615
rect 7230 15545 7600 15555
rect 7630 15875 8000 15885
rect 7630 15815 7634 15875
rect 7686 15855 7944 15875
rect 7630 15809 7686 15815
rect 7630 15621 7660 15809
rect 7715 15800 7915 15825
rect 7996 15815 8000 15875
rect 7944 15809 8000 15815
rect 7715 15780 7785 15800
rect 7690 15740 7785 15780
rect 7845 15780 7915 15800
rect 7845 15740 7940 15780
rect 7690 15690 7940 15740
rect 7690 15650 7785 15690
rect 7715 15630 7785 15650
rect 7845 15650 7940 15690
rect 7845 15630 7915 15650
rect 7630 15615 7686 15621
rect 7630 15555 7634 15615
rect 7715 15605 7915 15630
rect 7970 15621 8000 15809
rect 7944 15615 8000 15621
rect 7686 15555 7944 15575
rect 7996 15555 8000 15615
rect 7630 15545 8000 15555
rect 8030 15875 8400 15885
rect 8030 15815 8034 15875
rect 8086 15855 8344 15875
rect 8030 15809 8086 15815
rect 8030 15621 8060 15809
rect 8115 15800 8315 15825
rect 8396 15815 8400 15875
rect 8344 15809 8400 15815
rect 8115 15780 8185 15800
rect 8090 15740 8185 15780
rect 8245 15780 8315 15800
rect 8245 15740 8340 15780
rect 8090 15690 8340 15740
rect 8090 15650 8185 15690
rect 8115 15630 8185 15650
rect 8245 15650 8340 15690
rect 8245 15630 8315 15650
rect 8030 15615 8086 15621
rect 8030 15555 8034 15615
rect 8115 15605 8315 15630
rect 8370 15621 8400 15809
rect 8344 15615 8400 15621
rect 8086 15555 8344 15575
rect 8396 15555 8400 15615
rect 8030 15545 8400 15555
rect 8430 15875 8800 15885
rect 8430 15815 8434 15875
rect 8486 15855 8744 15875
rect 8430 15809 8486 15815
rect 8430 15621 8460 15809
rect 8515 15800 8715 15825
rect 8796 15815 8800 15875
rect 8744 15809 8800 15815
rect 8515 15780 8585 15800
rect 8490 15740 8585 15780
rect 8645 15780 8715 15800
rect 8645 15740 8740 15780
rect 8490 15690 8740 15740
rect 8490 15650 8585 15690
rect 8515 15630 8585 15650
rect 8645 15650 8740 15690
rect 8645 15630 8715 15650
rect 8430 15615 8486 15621
rect 8430 15555 8434 15615
rect 8515 15605 8715 15630
rect 8770 15621 8800 15809
rect 8744 15615 8800 15621
rect 8486 15555 8744 15575
rect 8796 15555 8800 15615
rect 8430 15545 8800 15555
rect 8830 15875 9200 15885
rect 8830 15815 8834 15875
rect 8886 15855 9144 15875
rect 8830 15809 8886 15815
rect 8830 15621 8860 15809
rect 8915 15800 9115 15825
rect 9196 15815 9200 15875
rect 9144 15809 9200 15815
rect 8915 15780 8985 15800
rect 8890 15740 8985 15780
rect 9045 15780 9115 15800
rect 9045 15740 9140 15780
rect 8890 15690 9140 15740
rect 8890 15650 8985 15690
rect 8915 15630 8985 15650
rect 9045 15650 9140 15690
rect 9045 15630 9115 15650
rect 8830 15615 8886 15621
rect 8830 15555 8834 15615
rect 8915 15605 9115 15630
rect 9170 15621 9200 15809
rect 9144 15615 9200 15621
rect 8886 15555 9144 15575
rect 9196 15555 9200 15615
rect 8830 15545 9200 15555
rect 9230 15875 9600 15885
rect 9230 15815 9234 15875
rect 9286 15855 9544 15875
rect 9230 15809 9286 15815
rect 9230 15621 9260 15809
rect 9315 15800 9515 15825
rect 9596 15815 9600 15875
rect 9544 15809 9600 15815
rect 9315 15780 9385 15800
rect 9290 15740 9385 15780
rect 9445 15780 9515 15800
rect 9445 15740 9540 15780
rect 9290 15690 9540 15740
rect 9290 15650 9385 15690
rect 9315 15630 9385 15650
rect 9445 15650 9540 15690
rect 9445 15630 9515 15650
rect 9230 15615 9286 15621
rect 9230 15555 9234 15615
rect 9315 15605 9515 15630
rect 9570 15621 9600 15809
rect 9544 15615 9600 15621
rect 9286 15555 9544 15575
rect 9596 15555 9600 15615
rect 9230 15545 9600 15555
rect 9630 15875 10000 15885
rect 9630 15815 9634 15875
rect 9686 15855 9944 15875
rect 9630 15809 9686 15815
rect 9630 15621 9660 15809
rect 9715 15800 9915 15825
rect 9996 15815 10000 15875
rect 9944 15809 10000 15815
rect 9715 15780 9785 15800
rect 9690 15740 9785 15780
rect 9845 15780 9915 15800
rect 9845 15740 9940 15780
rect 9690 15690 9940 15740
rect 9690 15650 9785 15690
rect 9715 15630 9785 15650
rect 9845 15650 9940 15690
rect 9845 15630 9915 15650
rect 9630 15615 9686 15621
rect 9630 15555 9634 15615
rect 9715 15605 9915 15630
rect 9970 15621 10000 15809
rect 9944 15615 10000 15621
rect 9686 15555 9944 15575
rect 9996 15555 10000 15615
rect 9630 15545 10000 15555
rect 10030 15875 10400 15885
rect 10030 15815 10034 15875
rect 10086 15855 10344 15875
rect 10030 15809 10086 15815
rect 10030 15621 10060 15809
rect 10115 15800 10315 15825
rect 10396 15815 10400 15875
rect 10344 15809 10400 15815
rect 10115 15780 10185 15800
rect 10090 15740 10185 15780
rect 10245 15780 10315 15800
rect 10245 15740 10340 15780
rect 10090 15690 10340 15740
rect 10090 15650 10185 15690
rect 10115 15630 10185 15650
rect 10245 15650 10340 15690
rect 10245 15630 10315 15650
rect 10030 15615 10086 15621
rect 10030 15555 10034 15615
rect 10115 15605 10315 15630
rect 10370 15621 10400 15809
rect 10344 15615 10400 15621
rect 10086 15555 10344 15575
rect 10396 15555 10400 15615
rect 10030 15545 10400 15555
rect 10430 15875 10800 15885
rect 10430 15815 10434 15875
rect 10486 15855 10744 15875
rect 10430 15809 10486 15815
rect 10430 15621 10460 15809
rect 10515 15800 10715 15825
rect 10796 15815 10800 15875
rect 10744 15809 10800 15815
rect 10515 15780 10585 15800
rect 10490 15740 10585 15780
rect 10645 15780 10715 15800
rect 10645 15740 10740 15780
rect 10490 15690 10740 15740
rect 10490 15650 10585 15690
rect 10515 15630 10585 15650
rect 10645 15650 10740 15690
rect 10645 15630 10715 15650
rect 10430 15615 10486 15621
rect 10430 15555 10434 15615
rect 10515 15605 10715 15630
rect 10770 15621 10800 15809
rect 10744 15615 10800 15621
rect 10486 15555 10744 15575
rect 10796 15555 10800 15615
rect 10430 15545 10800 15555
rect 10830 15875 11200 15885
rect 10830 15815 10834 15875
rect 10886 15855 11144 15875
rect 10830 15809 10886 15815
rect 10830 15621 10860 15809
rect 10915 15800 11115 15825
rect 11196 15815 11200 15875
rect 11144 15809 11200 15815
rect 10915 15780 10985 15800
rect 10890 15740 10985 15780
rect 11045 15780 11115 15800
rect 11045 15740 11140 15780
rect 10890 15690 11140 15740
rect 10890 15650 10985 15690
rect 10915 15630 10985 15650
rect 11045 15650 11140 15690
rect 11045 15630 11115 15650
rect 10830 15615 10886 15621
rect 10830 15555 10834 15615
rect 10915 15605 11115 15630
rect 11170 15621 11200 15809
rect 11144 15615 11200 15621
rect 10886 15555 11144 15575
rect 11196 15555 11200 15615
rect 10830 15545 11200 15555
rect 11230 15875 11600 15885
rect 11230 15815 11234 15875
rect 11286 15855 11544 15875
rect 11230 15809 11286 15815
rect 11230 15621 11260 15809
rect 11315 15800 11515 15825
rect 11596 15815 11600 15875
rect 11544 15809 11600 15815
rect 11315 15780 11385 15800
rect 11290 15740 11385 15780
rect 11445 15780 11515 15800
rect 11445 15740 11540 15780
rect 11290 15690 11540 15740
rect 11290 15650 11385 15690
rect 11315 15630 11385 15650
rect 11445 15650 11540 15690
rect 11445 15630 11515 15650
rect 11230 15615 11286 15621
rect 11230 15555 11234 15615
rect 11315 15605 11515 15630
rect 11570 15621 11600 15809
rect 11544 15615 11600 15621
rect 11286 15555 11544 15575
rect 11596 15555 11600 15615
rect 11230 15545 11600 15555
rect 11630 15875 12000 15885
rect 11630 15815 11634 15875
rect 11686 15855 11944 15875
rect 11630 15809 11686 15815
rect 11630 15621 11660 15809
rect 11715 15800 11915 15825
rect 11996 15815 12000 15875
rect 11944 15809 12000 15815
rect 11715 15780 11785 15800
rect 11690 15740 11785 15780
rect 11845 15780 11915 15800
rect 11845 15740 11940 15780
rect 11690 15690 11940 15740
rect 11690 15650 11785 15690
rect 11715 15630 11785 15650
rect 11845 15650 11940 15690
rect 11845 15630 11915 15650
rect 11630 15615 11686 15621
rect 11630 15555 11634 15615
rect 11715 15605 11915 15630
rect 11970 15621 12000 15809
rect 11944 15615 12000 15621
rect 11686 15555 11944 15575
rect 11996 15555 12000 15615
rect 11630 15545 12000 15555
rect 12030 15875 12400 15885
rect 12030 15815 12034 15875
rect 12086 15855 12344 15875
rect 12030 15809 12086 15815
rect 12030 15621 12060 15809
rect 12115 15800 12315 15825
rect 12396 15815 12400 15875
rect 12344 15809 12400 15815
rect 12115 15780 12185 15800
rect 12090 15740 12185 15780
rect 12245 15780 12315 15800
rect 12245 15740 12340 15780
rect 12090 15690 12340 15740
rect 12090 15650 12185 15690
rect 12115 15630 12185 15650
rect 12245 15650 12340 15690
rect 12245 15630 12315 15650
rect 12030 15615 12086 15621
rect 12030 15555 12034 15615
rect 12115 15605 12315 15630
rect 12370 15621 12400 15809
rect 12344 15615 12400 15621
rect 12086 15555 12344 15575
rect 12396 15555 12400 15615
rect 12030 15545 12400 15555
rect 12430 15875 12800 15885
rect 12430 15815 12434 15875
rect 12486 15855 12744 15875
rect 12430 15809 12486 15815
rect 12430 15621 12460 15809
rect 12515 15800 12715 15825
rect 12796 15815 12800 15875
rect 12744 15809 12800 15815
rect 12515 15780 12585 15800
rect 12490 15740 12585 15780
rect 12645 15780 12715 15800
rect 12645 15740 12740 15780
rect 12490 15690 12740 15740
rect 12490 15650 12585 15690
rect 12515 15630 12585 15650
rect 12645 15650 12740 15690
rect 12645 15630 12715 15650
rect 12430 15615 12486 15621
rect 12430 15555 12434 15615
rect 12515 15605 12715 15630
rect 12770 15621 12800 15809
rect 12744 15615 12800 15621
rect 12486 15555 12744 15575
rect 12796 15555 12800 15615
rect 12430 15545 12800 15555
rect 12830 15875 13200 15885
rect 12830 15815 12834 15875
rect 12886 15855 13144 15875
rect 12830 15809 12886 15815
rect 12830 15621 12860 15809
rect 12915 15800 13115 15825
rect 13196 15815 13200 15875
rect 13144 15809 13200 15815
rect 12915 15780 12985 15800
rect 12890 15740 12985 15780
rect 13045 15780 13115 15800
rect 13045 15740 13140 15780
rect 12890 15690 13140 15740
rect 12890 15650 12985 15690
rect 12915 15630 12985 15650
rect 13045 15650 13140 15690
rect 13045 15630 13115 15650
rect 12830 15615 12886 15621
rect 12830 15555 12834 15615
rect 12915 15605 13115 15630
rect 13170 15621 13200 15809
rect 13144 15615 13200 15621
rect 12886 15555 13144 15575
rect 13196 15555 13200 15615
rect 12830 15545 13200 15555
rect -370 15505 0 15515
rect -370 15445 -366 15505
rect -314 15485 -56 15505
rect -370 15439 -314 15445
rect -370 15251 -340 15439
rect -285 15430 -85 15455
rect -4 15445 0 15505
rect -56 15439 0 15445
rect -285 15410 -215 15430
rect -310 15370 -215 15410
rect -155 15410 -85 15430
rect -155 15370 -60 15410
rect -310 15320 -60 15370
rect -310 15280 -215 15320
rect -285 15260 -215 15280
rect -155 15280 -60 15320
rect -155 15260 -85 15280
rect -370 15245 -314 15251
rect -370 15185 -366 15245
rect -285 15235 -85 15260
rect -30 15251 0 15439
rect -56 15245 0 15251
rect -314 15185 -56 15205
rect -4 15185 0 15245
rect -370 15175 0 15185
rect 30 15505 400 15515
rect 30 15445 34 15505
rect 86 15485 344 15505
rect 30 15439 86 15445
rect 30 15251 60 15439
rect 115 15430 315 15455
rect 396 15445 400 15505
rect 344 15439 400 15445
rect 115 15410 185 15430
rect 90 15370 185 15410
rect 245 15410 315 15430
rect 245 15370 340 15410
rect 90 15320 340 15370
rect 90 15280 185 15320
rect 115 15260 185 15280
rect 245 15280 340 15320
rect 245 15260 315 15280
rect 30 15245 86 15251
rect 30 15185 34 15245
rect 115 15235 315 15260
rect 370 15251 400 15439
rect 344 15245 400 15251
rect 86 15185 344 15205
rect 396 15185 400 15245
rect 30 15175 400 15185
rect 430 15505 800 15515
rect 430 15445 434 15505
rect 486 15485 744 15505
rect 430 15439 486 15445
rect 430 15251 460 15439
rect 515 15430 715 15455
rect 796 15445 800 15505
rect 744 15439 800 15445
rect 515 15410 585 15430
rect 490 15370 585 15410
rect 645 15410 715 15430
rect 645 15370 740 15410
rect 490 15320 740 15370
rect 490 15280 585 15320
rect 515 15260 585 15280
rect 645 15280 740 15320
rect 645 15260 715 15280
rect 430 15245 486 15251
rect 430 15185 434 15245
rect 515 15235 715 15260
rect 770 15251 800 15439
rect 744 15245 800 15251
rect 486 15185 744 15205
rect 796 15185 800 15245
rect 430 15175 800 15185
rect 830 15505 1200 15515
rect 830 15445 834 15505
rect 886 15485 1144 15505
rect 830 15439 886 15445
rect 830 15251 860 15439
rect 915 15430 1115 15455
rect 1196 15445 1200 15505
rect 1144 15439 1200 15445
rect 915 15410 985 15430
rect 890 15370 985 15410
rect 1045 15410 1115 15430
rect 1045 15370 1140 15410
rect 890 15320 1140 15370
rect 890 15280 985 15320
rect 915 15260 985 15280
rect 1045 15280 1140 15320
rect 1045 15260 1115 15280
rect 830 15245 886 15251
rect 830 15185 834 15245
rect 915 15235 1115 15260
rect 1170 15251 1200 15439
rect 1144 15245 1200 15251
rect 886 15185 1144 15205
rect 1196 15185 1200 15245
rect 830 15175 1200 15185
rect 1230 15505 1600 15515
rect 1230 15445 1234 15505
rect 1286 15485 1544 15505
rect 1230 15439 1286 15445
rect 1230 15251 1260 15439
rect 1315 15430 1515 15455
rect 1596 15445 1600 15505
rect 1544 15439 1600 15445
rect 1315 15410 1385 15430
rect 1290 15370 1385 15410
rect 1445 15410 1515 15430
rect 1445 15370 1540 15410
rect 1290 15320 1540 15370
rect 1290 15280 1385 15320
rect 1315 15260 1385 15280
rect 1445 15280 1540 15320
rect 1445 15260 1515 15280
rect 1230 15245 1286 15251
rect 1230 15185 1234 15245
rect 1315 15235 1515 15260
rect 1570 15251 1600 15439
rect 1544 15245 1600 15251
rect 1286 15185 1544 15205
rect 1596 15185 1600 15245
rect 1230 15175 1600 15185
rect 1630 15505 2000 15515
rect 1630 15445 1634 15505
rect 1686 15485 1944 15505
rect 1630 15439 1686 15445
rect 1630 15251 1660 15439
rect 1715 15430 1915 15455
rect 1996 15445 2000 15505
rect 1944 15439 2000 15445
rect 1715 15410 1785 15430
rect 1690 15370 1785 15410
rect 1845 15410 1915 15430
rect 1845 15370 1940 15410
rect 1690 15320 1940 15370
rect 1690 15280 1785 15320
rect 1715 15260 1785 15280
rect 1845 15280 1940 15320
rect 1845 15260 1915 15280
rect 1630 15245 1686 15251
rect 1630 15185 1634 15245
rect 1715 15235 1915 15260
rect 1970 15251 2000 15439
rect 1944 15245 2000 15251
rect 1686 15185 1944 15205
rect 1996 15185 2000 15245
rect 1630 15175 2000 15185
rect 2030 15505 2400 15515
rect 2030 15445 2034 15505
rect 2086 15485 2344 15505
rect 2030 15439 2086 15445
rect 2030 15251 2060 15439
rect 2115 15430 2315 15455
rect 2396 15445 2400 15505
rect 2344 15439 2400 15445
rect 2115 15410 2185 15430
rect 2090 15370 2185 15410
rect 2245 15410 2315 15430
rect 2245 15370 2340 15410
rect 2090 15320 2340 15370
rect 2090 15280 2185 15320
rect 2115 15260 2185 15280
rect 2245 15280 2340 15320
rect 2245 15260 2315 15280
rect 2030 15245 2086 15251
rect 2030 15185 2034 15245
rect 2115 15235 2315 15260
rect 2370 15251 2400 15439
rect 2344 15245 2400 15251
rect 2086 15185 2344 15205
rect 2396 15185 2400 15245
rect 2030 15175 2400 15185
rect 2430 15505 2800 15515
rect 2430 15445 2434 15505
rect 2486 15485 2744 15505
rect 2430 15439 2486 15445
rect 2430 15251 2460 15439
rect 2515 15430 2715 15455
rect 2796 15445 2800 15505
rect 2744 15439 2800 15445
rect 2515 15410 2585 15430
rect 2490 15370 2585 15410
rect 2645 15410 2715 15430
rect 2645 15370 2740 15410
rect 2490 15320 2740 15370
rect 2490 15280 2585 15320
rect 2515 15260 2585 15280
rect 2645 15280 2740 15320
rect 2645 15260 2715 15280
rect 2430 15245 2486 15251
rect 2430 15185 2434 15245
rect 2515 15235 2715 15260
rect 2770 15251 2800 15439
rect 2744 15245 2800 15251
rect 2486 15185 2744 15205
rect 2796 15185 2800 15245
rect 2430 15175 2800 15185
rect 2830 15505 3200 15515
rect 2830 15445 2834 15505
rect 2886 15485 3144 15505
rect 2830 15439 2886 15445
rect 2830 15251 2860 15439
rect 2915 15430 3115 15455
rect 3196 15445 3200 15505
rect 3144 15439 3200 15445
rect 2915 15410 2985 15430
rect 2890 15370 2985 15410
rect 3045 15410 3115 15430
rect 3045 15370 3140 15410
rect 2890 15320 3140 15370
rect 2890 15280 2985 15320
rect 2915 15260 2985 15280
rect 3045 15280 3140 15320
rect 3045 15260 3115 15280
rect 2830 15245 2886 15251
rect 2830 15185 2834 15245
rect 2915 15235 3115 15260
rect 3170 15251 3200 15439
rect 3144 15245 3200 15251
rect 2886 15185 3144 15205
rect 3196 15185 3200 15245
rect 2830 15175 3200 15185
rect 3230 15505 3600 15515
rect 3230 15445 3234 15505
rect 3286 15485 3544 15505
rect 3230 15439 3286 15445
rect 3230 15251 3260 15439
rect 3315 15430 3515 15455
rect 3596 15445 3600 15505
rect 3544 15439 3600 15445
rect 3315 15410 3385 15430
rect 3290 15370 3385 15410
rect 3445 15410 3515 15430
rect 3445 15370 3540 15410
rect 3290 15320 3540 15370
rect 3290 15280 3385 15320
rect 3315 15260 3385 15280
rect 3445 15280 3540 15320
rect 3445 15260 3515 15280
rect 3230 15245 3286 15251
rect 3230 15185 3234 15245
rect 3315 15235 3515 15260
rect 3570 15251 3600 15439
rect 3544 15245 3600 15251
rect 3286 15185 3544 15205
rect 3596 15185 3600 15245
rect 3230 15175 3600 15185
rect 3630 15505 4000 15515
rect 3630 15445 3634 15505
rect 3686 15485 3944 15505
rect 3630 15439 3686 15445
rect 3630 15251 3660 15439
rect 3715 15430 3915 15455
rect 3996 15445 4000 15505
rect 3944 15439 4000 15445
rect 3715 15410 3785 15430
rect 3690 15370 3785 15410
rect 3845 15410 3915 15430
rect 3845 15370 3940 15410
rect 3690 15320 3940 15370
rect 3690 15280 3785 15320
rect 3715 15260 3785 15280
rect 3845 15280 3940 15320
rect 3845 15260 3915 15280
rect 3630 15245 3686 15251
rect 3630 15185 3634 15245
rect 3715 15235 3915 15260
rect 3970 15251 4000 15439
rect 3944 15245 4000 15251
rect 3686 15185 3944 15205
rect 3996 15185 4000 15245
rect 3630 15175 4000 15185
rect 4030 15505 4400 15515
rect 4030 15445 4034 15505
rect 4086 15485 4344 15505
rect 4030 15439 4086 15445
rect 4030 15251 4060 15439
rect 4115 15430 4315 15455
rect 4396 15445 4400 15505
rect 4344 15439 4400 15445
rect 4115 15410 4185 15430
rect 4090 15370 4185 15410
rect 4245 15410 4315 15430
rect 4245 15370 4340 15410
rect 4090 15320 4340 15370
rect 4090 15280 4185 15320
rect 4115 15260 4185 15280
rect 4245 15280 4340 15320
rect 4245 15260 4315 15280
rect 4030 15245 4086 15251
rect 4030 15185 4034 15245
rect 4115 15235 4315 15260
rect 4370 15251 4400 15439
rect 4344 15245 4400 15251
rect 4086 15185 4344 15205
rect 4396 15185 4400 15245
rect 4030 15175 4400 15185
rect 4430 15505 4800 15515
rect 4430 15445 4434 15505
rect 4486 15485 4744 15505
rect 4430 15439 4486 15445
rect 4430 15251 4460 15439
rect 4515 15430 4715 15455
rect 4796 15445 4800 15505
rect 4744 15439 4800 15445
rect 4515 15410 4585 15430
rect 4490 15370 4585 15410
rect 4645 15410 4715 15430
rect 4645 15370 4740 15410
rect 4490 15320 4740 15370
rect 4490 15280 4585 15320
rect 4515 15260 4585 15280
rect 4645 15280 4740 15320
rect 4645 15260 4715 15280
rect 4430 15245 4486 15251
rect 4430 15185 4434 15245
rect 4515 15235 4715 15260
rect 4770 15251 4800 15439
rect 4744 15245 4800 15251
rect 4486 15185 4744 15205
rect 4796 15185 4800 15245
rect 4430 15175 4800 15185
rect 4830 15505 5200 15515
rect 4830 15445 4834 15505
rect 4886 15485 5144 15505
rect 4830 15439 4886 15445
rect 4830 15251 4860 15439
rect 4915 15430 5115 15455
rect 5196 15445 5200 15505
rect 5144 15439 5200 15445
rect 4915 15410 4985 15430
rect 4890 15370 4985 15410
rect 5045 15410 5115 15430
rect 5045 15370 5140 15410
rect 4890 15320 5140 15370
rect 4890 15280 4985 15320
rect 4915 15260 4985 15280
rect 5045 15280 5140 15320
rect 5045 15260 5115 15280
rect 4830 15245 4886 15251
rect 4830 15185 4834 15245
rect 4915 15235 5115 15260
rect 5170 15251 5200 15439
rect 5144 15245 5200 15251
rect 4886 15185 5144 15205
rect 5196 15185 5200 15245
rect 4830 15175 5200 15185
rect 5230 15505 5600 15515
rect 5230 15445 5234 15505
rect 5286 15485 5544 15505
rect 5230 15439 5286 15445
rect 5230 15251 5260 15439
rect 5315 15430 5515 15455
rect 5596 15445 5600 15505
rect 5544 15439 5600 15445
rect 5315 15410 5385 15430
rect 5290 15370 5385 15410
rect 5445 15410 5515 15430
rect 5445 15370 5540 15410
rect 5290 15320 5540 15370
rect 5290 15280 5385 15320
rect 5315 15260 5385 15280
rect 5445 15280 5540 15320
rect 5445 15260 5515 15280
rect 5230 15245 5286 15251
rect 5230 15185 5234 15245
rect 5315 15235 5515 15260
rect 5570 15251 5600 15439
rect 5544 15245 5600 15251
rect 5286 15185 5544 15205
rect 5596 15185 5600 15245
rect 5230 15175 5600 15185
rect 5630 15505 6000 15515
rect 5630 15445 5634 15505
rect 5686 15485 5944 15505
rect 5630 15439 5686 15445
rect 5630 15251 5660 15439
rect 5715 15430 5915 15455
rect 5996 15445 6000 15505
rect 5944 15439 6000 15445
rect 5715 15410 5785 15430
rect 5690 15370 5785 15410
rect 5845 15410 5915 15430
rect 5845 15370 5940 15410
rect 5690 15320 5940 15370
rect 5690 15280 5785 15320
rect 5715 15260 5785 15280
rect 5845 15280 5940 15320
rect 5845 15260 5915 15280
rect 5630 15245 5686 15251
rect 5630 15185 5634 15245
rect 5715 15235 5915 15260
rect 5970 15251 6000 15439
rect 5944 15245 6000 15251
rect 5686 15185 5944 15205
rect 5996 15185 6000 15245
rect 5630 15175 6000 15185
rect 6030 15505 6400 15515
rect 6030 15445 6034 15505
rect 6086 15485 6344 15505
rect 6030 15439 6086 15445
rect 6030 15251 6060 15439
rect 6115 15430 6315 15455
rect 6396 15445 6400 15505
rect 6344 15439 6400 15445
rect 6115 15410 6185 15430
rect 6090 15370 6185 15410
rect 6245 15410 6315 15430
rect 6245 15370 6340 15410
rect 6090 15320 6340 15370
rect 6090 15280 6185 15320
rect 6115 15260 6185 15280
rect 6245 15280 6340 15320
rect 6245 15260 6315 15280
rect 6030 15245 6086 15251
rect 6030 15185 6034 15245
rect 6115 15235 6315 15260
rect 6370 15251 6400 15439
rect 6344 15245 6400 15251
rect 6086 15185 6344 15205
rect 6396 15185 6400 15245
rect 6030 15175 6400 15185
rect 6430 15505 6800 15515
rect 6430 15445 6434 15505
rect 6486 15485 6744 15505
rect 6430 15439 6486 15445
rect 6430 15251 6460 15439
rect 6515 15430 6715 15455
rect 6796 15445 6800 15505
rect 6744 15439 6800 15445
rect 6515 15410 6585 15430
rect 6490 15370 6585 15410
rect 6645 15410 6715 15430
rect 6645 15370 6740 15410
rect 6490 15320 6740 15370
rect 6490 15280 6585 15320
rect 6515 15260 6585 15280
rect 6645 15280 6740 15320
rect 6645 15260 6715 15280
rect 6430 15245 6486 15251
rect 6430 15185 6434 15245
rect 6515 15235 6715 15260
rect 6770 15251 6800 15439
rect 6744 15245 6800 15251
rect 6486 15185 6744 15205
rect 6796 15185 6800 15245
rect 6430 15175 6800 15185
rect 6830 15505 7200 15515
rect 6830 15445 6834 15505
rect 6886 15485 7144 15505
rect 6830 15439 6886 15445
rect 6830 15251 6860 15439
rect 6915 15430 7115 15455
rect 7196 15445 7200 15505
rect 7144 15439 7200 15445
rect 6915 15410 6985 15430
rect 6890 15370 6985 15410
rect 7045 15410 7115 15430
rect 7045 15370 7140 15410
rect 6890 15320 7140 15370
rect 6890 15280 6985 15320
rect 6915 15260 6985 15280
rect 7045 15280 7140 15320
rect 7045 15260 7115 15280
rect 6830 15245 6886 15251
rect 6830 15185 6834 15245
rect 6915 15235 7115 15260
rect 7170 15251 7200 15439
rect 7144 15245 7200 15251
rect 6886 15185 7144 15205
rect 7196 15185 7200 15245
rect 6830 15175 7200 15185
rect 7230 15505 7600 15515
rect 7230 15445 7234 15505
rect 7286 15485 7544 15505
rect 7230 15439 7286 15445
rect 7230 15251 7260 15439
rect 7315 15430 7515 15455
rect 7596 15445 7600 15505
rect 7544 15439 7600 15445
rect 7315 15410 7385 15430
rect 7290 15370 7385 15410
rect 7445 15410 7515 15430
rect 7445 15370 7540 15410
rect 7290 15320 7540 15370
rect 7290 15280 7385 15320
rect 7315 15260 7385 15280
rect 7445 15280 7540 15320
rect 7445 15260 7515 15280
rect 7230 15245 7286 15251
rect 7230 15185 7234 15245
rect 7315 15235 7515 15260
rect 7570 15251 7600 15439
rect 7544 15245 7600 15251
rect 7286 15185 7544 15205
rect 7596 15185 7600 15245
rect 7230 15175 7600 15185
rect 7630 15505 8000 15515
rect 7630 15445 7634 15505
rect 7686 15485 7944 15505
rect 7630 15439 7686 15445
rect 7630 15251 7660 15439
rect 7715 15430 7915 15455
rect 7996 15445 8000 15505
rect 7944 15439 8000 15445
rect 7715 15410 7785 15430
rect 7690 15370 7785 15410
rect 7845 15410 7915 15430
rect 7845 15370 7940 15410
rect 7690 15320 7940 15370
rect 7690 15280 7785 15320
rect 7715 15260 7785 15280
rect 7845 15280 7940 15320
rect 7845 15260 7915 15280
rect 7630 15245 7686 15251
rect 7630 15185 7634 15245
rect 7715 15235 7915 15260
rect 7970 15251 8000 15439
rect 7944 15245 8000 15251
rect 7686 15185 7944 15205
rect 7996 15185 8000 15245
rect 7630 15175 8000 15185
rect 8030 15505 8400 15515
rect 8030 15445 8034 15505
rect 8086 15485 8344 15505
rect 8030 15439 8086 15445
rect 8030 15251 8060 15439
rect 8115 15430 8315 15455
rect 8396 15445 8400 15505
rect 8344 15439 8400 15445
rect 8115 15410 8185 15430
rect 8090 15370 8185 15410
rect 8245 15410 8315 15430
rect 8245 15370 8340 15410
rect 8090 15320 8340 15370
rect 8090 15280 8185 15320
rect 8115 15260 8185 15280
rect 8245 15280 8340 15320
rect 8245 15260 8315 15280
rect 8030 15245 8086 15251
rect 8030 15185 8034 15245
rect 8115 15235 8315 15260
rect 8370 15251 8400 15439
rect 8344 15245 8400 15251
rect 8086 15185 8344 15205
rect 8396 15185 8400 15245
rect 8030 15175 8400 15185
rect 8430 15505 8800 15515
rect 8430 15445 8434 15505
rect 8486 15485 8744 15505
rect 8430 15439 8486 15445
rect 8430 15251 8460 15439
rect 8515 15430 8715 15455
rect 8796 15445 8800 15505
rect 8744 15439 8800 15445
rect 8515 15410 8585 15430
rect 8490 15370 8585 15410
rect 8645 15410 8715 15430
rect 8645 15370 8740 15410
rect 8490 15320 8740 15370
rect 8490 15280 8585 15320
rect 8515 15260 8585 15280
rect 8645 15280 8740 15320
rect 8645 15260 8715 15280
rect 8430 15245 8486 15251
rect 8430 15185 8434 15245
rect 8515 15235 8715 15260
rect 8770 15251 8800 15439
rect 8744 15245 8800 15251
rect 8486 15185 8744 15205
rect 8796 15185 8800 15245
rect 8430 15175 8800 15185
rect 8830 15505 9200 15515
rect 8830 15445 8834 15505
rect 8886 15485 9144 15505
rect 8830 15439 8886 15445
rect 8830 15251 8860 15439
rect 8915 15430 9115 15455
rect 9196 15445 9200 15505
rect 9144 15439 9200 15445
rect 8915 15410 8985 15430
rect 8890 15370 8985 15410
rect 9045 15410 9115 15430
rect 9045 15370 9140 15410
rect 8890 15320 9140 15370
rect 8890 15280 8985 15320
rect 8915 15260 8985 15280
rect 9045 15280 9140 15320
rect 9045 15260 9115 15280
rect 8830 15245 8886 15251
rect 8830 15185 8834 15245
rect 8915 15235 9115 15260
rect 9170 15251 9200 15439
rect 9144 15245 9200 15251
rect 8886 15185 9144 15205
rect 9196 15185 9200 15245
rect 8830 15175 9200 15185
rect 9230 15505 9600 15515
rect 9230 15445 9234 15505
rect 9286 15485 9544 15505
rect 9230 15439 9286 15445
rect 9230 15251 9260 15439
rect 9315 15430 9515 15455
rect 9596 15445 9600 15505
rect 9544 15439 9600 15445
rect 9315 15410 9385 15430
rect 9290 15370 9385 15410
rect 9445 15410 9515 15430
rect 9445 15370 9540 15410
rect 9290 15320 9540 15370
rect 9290 15280 9385 15320
rect 9315 15260 9385 15280
rect 9445 15280 9540 15320
rect 9445 15260 9515 15280
rect 9230 15245 9286 15251
rect 9230 15185 9234 15245
rect 9315 15235 9515 15260
rect 9570 15251 9600 15439
rect 9544 15245 9600 15251
rect 9286 15185 9544 15205
rect 9596 15185 9600 15245
rect 9230 15175 9600 15185
rect 9630 15505 10000 15515
rect 9630 15445 9634 15505
rect 9686 15485 9944 15505
rect 9630 15439 9686 15445
rect 9630 15251 9660 15439
rect 9715 15430 9915 15455
rect 9996 15445 10000 15505
rect 9944 15439 10000 15445
rect 9715 15410 9785 15430
rect 9690 15370 9785 15410
rect 9845 15410 9915 15430
rect 9845 15370 9940 15410
rect 9690 15320 9940 15370
rect 9690 15280 9785 15320
rect 9715 15260 9785 15280
rect 9845 15280 9940 15320
rect 9845 15260 9915 15280
rect 9630 15245 9686 15251
rect 9630 15185 9634 15245
rect 9715 15235 9915 15260
rect 9970 15251 10000 15439
rect 9944 15245 10000 15251
rect 9686 15185 9944 15205
rect 9996 15185 10000 15245
rect 9630 15175 10000 15185
rect 10030 15505 10400 15515
rect 10030 15445 10034 15505
rect 10086 15485 10344 15505
rect 10030 15439 10086 15445
rect 10030 15251 10060 15439
rect 10115 15430 10315 15455
rect 10396 15445 10400 15505
rect 10344 15439 10400 15445
rect 10115 15410 10185 15430
rect 10090 15370 10185 15410
rect 10245 15410 10315 15430
rect 10245 15370 10340 15410
rect 10090 15320 10340 15370
rect 10090 15280 10185 15320
rect 10115 15260 10185 15280
rect 10245 15280 10340 15320
rect 10245 15260 10315 15280
rect 10030 15245 10086 15251
rect 10030 15185 10034 15245
rect 10115 15235 10315 15260
rect 10370 15251 10400 15439
rect 10344 15245 10400 15251
rect 10086 15185 10344 15205
rect 10396 15185 10400 15245
rect 10030 15175 10400 15185
rect 10430 15505 10800 15515
rect 10430 15445 10434 15505
rect 10486 15485 10744 15505
rect 10430 15439 10486 15445
rect 10430 15251 10460 15439
rect 10515 15430 10715 15455
rect 10796 15445 10800 15505
rect 10744 15439 10800 15445
rect 10515 15410 10585 15430
rect 10490 15370 10585 15410
rect 10645 15410 10715 15430
rect 10645 15370 10740 15410
rect 10490 15320 10740 15370
rect 10490 15280 10585 15320
rect 10515 15260 10585 15280
rect 10645 15280 10740 15320
rect 10645 15260 10715 15280
rect 10430 15245 10486 15251
rect 10430 15185 10434 15245
rect 10515 15235 10715 15260
rect 10770 15251 10800 15439
rect 10744 15245 10800 15251
rect 10486 15185 10744 15205
rect 10796 15185 10800 15245
rect 10430 15175 10800 15185
rect 10830 15505 11200 15515
rect 10830 15445 10834 15505
rect 10886 15485 11144 15505
rect 10830 15439 10886 15445
rect 10830 15251 10860 15439
rect 10915 15430 11115 15455
rect 11196 15445 11200 15505
rect 11144 15439 11200 15445
rect 10915 15410 10985 15430
rect 10890 15370 10985 15410
rect 11045 15410 11115 15430
rect 11045 15370 11140 15410
rect 10890 15320 11140 15370
rect 10890 15280 10985 15320
rect 10915 15260 10985 15280
rect 11045 15280 11140 15320
rect 11045 15260 11115 15280
rect 10830 15245 10886 15251
rect 10830 15185 10834 15245
rect 10915 15235 11115 15260
rect 11170 15251 11200 15439
rect 11144 15245 11200 15251
rect 10886 15185 11144 15205
rect 11196 15185 11200 15245
rect 10830 15175 11200 15185
rect 11230 15505 11600 15515
rect 11230 15445 11234 15505
rect 11286 15485 11544 15505
rect 11230 15439 11286 15445
rect 11230 15251 11260 15439
rect 11315 15430 11515 15455
rect 11596 15445 11600 15505
rect 11544 15439 11600 15445
rect 11315 15410 11385 15430
rect 11290 15370 11385 15410
rect 11445 15410 11515 15430
rect 11445 15370 11540 15410
rect 11290 15320 11540 15370
rect 11290 15280 11385 15320
rect 11315 15260 11385 15280
rect 11445 15280 11540 15320
rect 11445 15260 11515 15280
rect 11230 15245 11286 15251
rect 11230 15185 11234 15245
rect 11315 15235 11515 15260
rect 11570 15251 11600 15439
rect 11544 15245 11600 15251
rect 11286 15185 11544 15205
rect 11596 15185 11600 15245
rect 11230 15175 11600 15185
rect 11630 15505 12000 15515
rect 11630 15445 11634 15505
rect 11686 15485 11944 15505
rect 11630 15439 11686 15445
rect 11630 15251 11660 15439
rect 11715 15430 11915 15455
rect 11996 15445 12000 15505
rect 11944 15439 12000 15445
rect 11715 15410 11785 15430
rect 11690 15370 11785 15410
rect 11845 15410 11915 15430
rect 11845 15370 11940 15410
rect 11690 15320 11940 15370
rect 11690 15280 11785 15320
rect 11715 15260 11785 15280
rect 11845 15280 11940 15320
rect 11845 15260 11915 15280
rect 11630 15245 11686 15251
rect 11630 15185 11634 15245
rect 11715 15235 11915 15260
rect 11970 15251 12000 15439
rect 11944 15245 12000 15251
rect 11686 15185 11944 15205
rect 11996 15185 12000 15245
rect 11630 15175 12000 15185
rect 12030 15505 12400 15515
rect 12030 15445 12034 15505
rect 12086 15485 12344 15505
rect 12030 15439 12086 15445
rect 12030 15251 12060 15439
rect 12115 15430 12315 15455
rect 12396 15445 12400 15505
rect 12344 15439 12400 15445
rect 12115 15410 12185 15430
rect 12090 15370 12185 15410
rect 12245 15410 12315 15430
rect 12245 15370 12340 15410
rect 12090 15320 12340 15370
rect 12090 15280 12185 15320
rect 12115 15260 12185 15280
rect 12245 15280 12340 15320
rect 12245 15260 12315 15280
rect 12030 15245 12086 15251
rect 12030 15185 12034 15245
rect 12115 15235 12315 15260
rect 12370 15251 12400 15439
rect 12344 15245 12400 15251
rect 12086 15185 12344 15205
rect 12396 15185 12400 15245
rect 12030 15175 12400 15185
rect 12430 15505 12800 15515
rect 12430 15445 12434 15505
rect 12486 15485 12744 15505
rect 12430 15439 12486 15445
rect 12430 15251 12460 15439
rect 12515 15430 12715 15455
rect 12796 15445 12800 15505
rect 12744 15439 12800 15445
rect 12515 15410 12585 15430
rect 12490 15370 12585 15410
rect 12645 15410 12715 15430
rect 12645 15370 12740 15410
rect 12490 15320 12740 15370
rect 12490 15280 12585 15320
rect 12515 15260 12585 15280
rect 12645 15280 12740 15320
rect 12645 15260 12715 15280
rect 12430 15245 12486 15251
rect 12430 15185 12434 15245
rect 12515 15235 12715 15260
rect 12770 15251 12800 15439
rect 12744 15245 12800 15251
rect 12486 15185 12744 15205
rect 12796 15185 12800 15245
rect 12430 15175 12800 15185
rect 12830 15505 13200 15515
rect 12830 15445 12834 15505
rect 12886 15485 13144 15505
rect 12830 15439 12886 15445
rect 12830 15251 12860 15439
rect 12915 15430 13115 15455
rect 13196 15445 13200 15505
rect 13144 15439 13200 15445
rect 12915 15410 12985 15430
rect 12890 15370 12985 15410
rect 13045 15410 13115 15430
rect 13045 15370 13140 15410
rect 12890 15320 13140 15370
rect 12890 15280 12985 15320
rect 12915 15260 12985 15280
rect 13045 15280 13140 15320
rect 13045 15260 13115 15280
rect 12830 15245 12886 15251
rect 12830 15185 12834 15245
rect 12915 15235 13115 15260
rect 13170 15251 13200 15439
rect 13144 15245 13200 15251
rect 12886 15185 13144 15205
rect 13196 15185 13200 15245
rect 12830 15175 13200 15185
rect -370 15135 0 15145
rect -370 15075 -366 15135
rect -314 15115 -56 15135
rect -370 15069 -314 15075
rect -370 14881 -340 15069
rect -285 15060 -85 15085
rect -4 15075 0 15135
rect -56 15069 0 15075
rect -285 15040 -215 15060
rect -310 15000 -215 15040
rect -155 15040 -85 15060
rect -155 15000 -60 15040
rect -310 14950 -60 15000
rect -310 14910 -215 14950
rect -285 14890 -215 14910
rect -155 14910 -60 14950
rect -155 14890 -85 14910
rect -370 14875 -314 14881
rect -370 14815 -366 14875
rect -285 14865 -85 14890
rect -30 14881 0 15069
rect -56 14875 0 14881
rect -314 14815 -56 14835
rect -4 14815 0 14875
rect -370 14805 0 14815
rect 30 15135 400 15145
rect 30 15075 34 15135
rect 86 15115 344 15135
rect 30 15069 86 15075
rect 30 14881 60 15069
rect 115 15060 315 15085
rect 396 15075 400 15135
rect 344 15069 400 15075
rect 115 15040 185 15060
rect 90 15000 185 15040
rect 245 15040 315 15060
rect 245 15000 340 15040
rect 90 14950 340 15000
rect 90 14910 185 14950
rect 115 14890 185 14910
rect 245 14910 340 14950
rect 245 14890 315 14910
rect 30 14875 86 14881
rect 30 14815 34 14875
rect 115 14865 315 14890
rect 370 14881 400 15069
rect 344 14875 400 14881
rect 86 14815 344 14835
rect 396 14815 400 14875
rect 30 14805 400 14815
rect 430 15135 800 15145
rect 430 15075 434 15135
rect 486 15115 744 15135
rect 430 15069 486 15075
rect 430 14881 460 15069
rect 515 15060 715 15085
rect 796 15075 800 15135
rect 744 15069 800 15075
rect 515 15040 585 15060
rect 490 15000 585 15040
rect 645 15040 715 15060
rect 645 15000 740 15040
rect 490 14950 740 15000
rect 490 14910 585 14950
rect 515 14890 585 14910
rect 645 14910 740 14950
rect 645 14890 715 14910
rect 430 14875 486 14881
rect 430 14815 434 14875
rect 515 14865 715 14890
rect 770 14881 800 15069
rect 744 14875 800 14881
rect 486 14815 744 14835
rect 796 14815 800 14875
rect 430 14805 800 14815
rect 830 15135 1200 15145
rect 830 15075 834 15135
rect 886 15115 1144 15135
rect 830 15069 886 15075
rect 830 14881 860 15069
rect 915 15060 1115 15085
rect 1196 15075 1200 15135
rect 1144 15069 1200 15075
rect 915 15040 985 15060
rect 890 15000 985 15040
rect 1045 15040 1115 15060
rect 1045 15000 1140 15040
rect 890 14950 1140 15000
rect 890 14910 985 14950
rect 915 14890 985 14910
rect 1045 14910 1140 14950
rect 1045 14890 1115 14910
rect 830 14875 886 14881
rect 830 14815 834 14875
rect 915 14865 1115 14890
rect 1170 14881 1200 15069
rect 1144 14875 1200 14881
rect 886 14815 1144 14835
rect 1196 14815 1200 14875
rect 830 14805 1200 14815
rect 1230 15135 1600 15145
rect 1230 15075 1234 15135
rect 1286 15115 1544 15135
rect 1230 15069 1286 15075
rect 1230 14881 1260 15069
rect 1315 15060 1515 15085
rect 1596 15075 1600 15135
rect 1544 15069 1600 15075
rect 1315 15040 1385 15060
rect 1290 15000 1385 15040
rect 1445 15040 1515 15060
rect 1445 15000 1540 15040
rect 1290 14950 1540 15000
rect 1290 14910 1385 14950
rect 1315 14890 1385 14910
rect 1445 14910 1540 14950
rect 1445 14890 1515 14910
rect 1230 14875 1286 14881
rect 1230 14815 1234 14875
rect 1315 14865 1515 14890
rect 1570 14881 1600 15069
rect 1544 14875 1600 14881
rect 1286 14815 1544 14835
rect 1596 14815 1600 14875
rect 1230 14805 1600 14815
rect 1630 15135 2000 15145
rect 1630 15075 1634 15135
rect 1686 15115 1944 15135
rect 1630 15069 1686 15075
rect 1630 14881 1660 15069
rect 1715 15060 1915 15085
rect 1996 15075 2000 15135
rect 1944 15069 2000 15075
rect 1715 15040 1785 15060
rect 1690 15000 1785 15040
rect 1845 15040 1915 15060
rect 1845 15000 1940 15040
rect 1690 14950 1940 15000
rect 1690 14910 1785 14950
rect 1715 14890 1785 14910
rect 1845 14910 1940 14950
rect 1845 14890 1915 14910
rect 1630 14875 1686 14881
rect 1630 14815 1634 14875
rect 1715 14865 1915 14890
rect 1970 14881 2000 15069
rect 1944 14875 2000 14881
rect 1686 14815 1944 14835
rect 1996 14815 2000 14875
rect 1630 14805 2000 14815
rect 2030 15135 2400 15145
rect 2030 15075 2034 15135
rect 2086 15115 2344 15135
rect 2030 15069 2086 15075
rect 2030 14881 2060 15069
rect 2115 15060 2315 15085
rect 2396 15075 2400 15135
rect 2344 15069 2400 15075
rect 2115 15040 2185 15060
rect 2090 15000 2185 15040
rect 2245 15040 2315 15060
rect 2245 15000 2340 15040
rect 2090 14950 2340 15000
rect 2090 14910 2185 14950
rect 2115 14890 2185 14910
rect 2245 14910 2340 14950
rect 2245 14890 2315 14910
rect 2030 14875 2086 14881
rect 2030 14815 2034 14875
rect 2115 14865 2315 14890
rect 2370 14881 2400 15069
rect 2344 14875 2400 14881
rect 2086 14815 2344 14835
rect 2396 14815 2400 14875
rect 2030 14805 2400 14815
rect 2430 15135 2800 15145
rect 2430 15075 2434 15135
rect 2486 15115 2744 15135
rect 2430 15069 2486 15075
rect 2430 14881 2460 15069
rect 2515 15060 2715 15085
rect 2796 15075 2800 15135
rect 2744 15069 2800 15075
rect 2515 15040 2585 15060
rect 2490 15000 2585 15040
rect 2645 15040 2715 15060
rect 2645 15000 2740 15040
rect 2490 14950 2740 15000
rect 2490 14910 2585 14950
rect 2515 14890 2585 14910
rect 2645 14910 2740 14950
rect 2645 14890 2715 14910
rect 2430 14875 2486 14881
rect 2430 14815 2434 14875
rect 2515 14865 2715 14890
rect 2770 14881 2800 15069
rect 2744 14875 2800 14881
rect 2486 14815 2744 14835
rect 2796 14815 2800 14875
rect 2430 14805 2800 14815
rect 2830 15135 3200 15145
rect 2830 15075 2834 15135
rect 2886 15115 3144 15135
rect 2830 15069 2886 15075
rect 2830 14881 2860 15069
rect 2915 15060 3115 15085
rect 3196 15075 3200 15135
rect 3144 15069 3200 15075
rect 2915 15040 2985 15060
rect 2890 15000 2985 15040
rect 3045 15040 3115 15060
rect 3045 15000 3140 15040
rect 2890 14950 3140 15000
rect 2890 14910 2985 14950
rect 2915 14890 2985 14910
rect 3045 14910 3140 14950
rect 3045 14890 3115 14910
rect 2830 14875 2886 14881
rect 2830 14815 2834 14875
rect 2915 14865 3115 14890
rect 3170 14881 3200 15069
rect 3144 14875 3200 14881
rect 2886 14815 3144 14835
rect 3196 14815 3200 14875
rect 2830 14805 3200 14815
rect 3230 15135 3600 15145
rect 3230 15075 3234 15135
rect 3286 15115 3544 15135
rect 3230 15069 3286 15075
rect 3230 14881 3260 15069
rect 3315 15060 3515 15085
rect 3596 15075 3600 15135
rect 3544 15069 3600 15075
rect 3315 15040 3385 15060
rect 3290 15000 3385 15040
rect 3445 15040 3515 15060
rect 3445 15000 3540 15040
rect 3290 14950 3540 15000
rect 3290 14910 3385 14950
rect 3315 14890 3385 14910
rect 3445 14910 3540 14950
rect 3445 14890 3515 14910
rect 3230 14875 3286 14881
rect 3230 14815 3234 14875
rect 3315 14865 3515 14890
rect 3570 14881 3600 15069
rect 3544 14875 3600 14881
rect 3286 14815 3544 14835
rect 3596 14815 3600 14875
rect 3230 14805 3600 14815
rect 3630 15135 4000 15145
rect 3630 15075 3634 15135
rect 3686 15115 3944 15135
rect 3630 15069 3686 15075
rect 3630 14881 3660 15069
rect 3715 15060 3915 15085
rect 3996 15075 4000 15135
rect 3944 15069 4000 15075
rect 3715 15040 3785 15060
rect 3690 15000 3785 15040
rect 3845 15040 3915 15060
rect 3845 15000 3940 15040
rect 3690 14950 3940 15000
rect 3690 14910 3785 14950
rect 3715 14890 3785 14910
rect 3845 14910 3940 14950
rect 3845 14890 3915 14910
rect 3630 14875 3686 14881
rect 3630 14815 3634 14875
rect 3715 14865 3915 14890
rect 3970 14881 4000 15069
rect 3944 14875 4000 14881
rect 3686 14815 3944 14835
rect 3996 14815 4000 14875
rect 3630 14805 4000 14815
rect 4030 15135 4400 15145
rect 4030 15075 4034 15135
rect 4086 15115 4344 15135
rect 4030 15069 4086 15075
rect 4030 14881 4060 15069
rect 4115 15060 4315 15085
rect 4396 15075 4400 15135
rect 4344 15069 4400 15075
rect 4115 15040 4185 15060
rect 4090 15000 4185 15040
rect 4245 15040 4315 15060
rect 4245 15000 4340 15040
rect 4090 14950 4340 15000
rect 4090 14910 4185 14950
rect 4115 14890 4185 14910
rect 4245 14910 4340 14950
rect 4245 14890 4315 14910
rect 4030 14875 4086 14881
rect 4030 14815 4034 14875
rect 4115 14865 4315 14890
rect 4370 14881 4400 15069
rect 4344 14875 4400 14881
rect 4086 14815 4344 14835
rect 4396 14815 4400 14875
rect 4030 14805 4400 14815
rect 4430 15135 4800 15145
rect 4430 15075 4434 15135
rect 4486 15115 4744 15135
rect 4430 15069 4486 15075
rect 4430 14881 4460 15069
rect 4515 15060 4715 15085
rect 4796 15075 4800 15135
rect 4744 15069 4800 15075
rect 4515 15040 4585 15060
rect 4490 15000 4585 15040
rect 4645 15040 4715 15060
rect 4645 15000 4740 15040
rect 4490 14950 4740 15000
rect 4490 14910 4585 14950
rect 4515 14890 4585 14910
rect 4645 14910 4740 14950
rect 4645 14890 4715 14910
rect 4430 14875 4486 14881
rect 4430 14815 4434 14875
rect 4515 14865 4715 14890
rect 4770 14881 4800 15069
rect 4744 14875 4800 14881
rect 4486 14815 4744 14835
rect 4796 14815 4800 14875
rect 4430 14805 4800 14815
rect 4830 15135 5200 15145
rect 4830 15075 4834 15135
rect 4886 15115 5144 15135
rect 4830 15069 4886 15075
rect 4830 14881 4860 15069
rect 4915 15060 5115 15085
rect 5196 15075 5200 15135
rect 5144 15069 5200 15075
rect 4915 15040 4985 15060
rect 4890 15000 4985 15040
rect 5045 15040 5115 15060
rect 5045 15000 5140 15040
rect 4890 14950 5140 15000
rect 4890 14910 4985 14950
rect 4915 14890 4985 14910
rect 5045 14910 5140 14950
rect 5045 14890 5115 14910
rect 4830 14875 4886 14881
rect 4830 14815 4834 14875
rect 4915 14865 5115 14890
rect 5170 14881 5200 15069
rect 5144 14875 5200 14881
rect 4886 14815 5144 14835
rect 5196 14815 5200 14875
rect 4830 14805 5200 14815
rect 5230 15135 5600 15145
rect 5230 15075 5234 15135
rect 5286 15115 5544 15135
rect 5230 15069 5286 15075
rect 5230 14881 5260 15069
rect 5315 15060 5515 15085
rect 5596 15075 5600 15135
rect 5544 15069 5600 15075
rect 5315 15040 5385 15060
rect 5290 15000 5385 15040
rect 5445 15040 5515 15060
rect 5445 15000 5540 15040
rect 5290 14950 5540 15000
rect 5290 14910 5385 14950
rect 5315 14890 5385 14910
rect 5445 14910 5540 14950
rect 5445 14890 5515 14910
rect 5230 14875 5286 14881
rect 5230 14815 5234 14875
rect 5315 14865 5515 14890
rect 5570 14881 5600 15069
rect 5544 14875 5600 14881
rect 5286 14815 5544 14835
rect 5596 14815 5600 14875
rect 5230 14805 5600 14815
rect 5630 15135 6000 15145
rect 5630 15075 5634 15135
rect 5686 15115 5944 15135
rect 5630 15069 5686 15075
rect 5630 14881 5660 15069
rect 5715 15060 5915 15085
rect 5996 15075 6000 15135
rect 5944 15069 6000 15075
rect 5715 15040 5785 15060
rect 5690 15000 5785 15040
rect 5845 15040 5915 15060
rect 5845 15000 5940 15040
rect 5690 14950 5940 15000
rect 5690 14910 5785 14950
rect 5715 14890 5785 14910
rect 5845 14910 5940 14950
rect 5845 14890 5915 14910
rect 5630 14875 5686 14881
rect 5630 14815 5634 14875
rect 5715 14865 5915 14890
rect 5970 14881 6000 15069
rect 5944 14875 6000 14881
rect 5686 14815 5944 14835
rect 5996 14815 6000 14875
rect 5630 14805 6000 14815
rect 6030 15135 6400 15145
rect 6030 15075 6034 15135
rect 6086 15115 6344 15135
rect 6030 15069 6086 15075
rect 6030 14881 6060 15069
rect 6115 15060 6315 15085
rect 6396 15075 6400 15135
rect 6344 15069 6400 15075
rect 6115 15040 6185 15060
rect 6090 15000 6185 15040
rect 6245 15040 6315 15060
rect 6245 15000 6340 15040
rect 6090 14950 6340 15000
rect 6090 14910 6185 14950
rect 6115 14890 6185 14910
rect 6245 14910 6340 14950
rect 6245 14890 6315 14910
rect 6030 14875 6086 14881
rect 6030 14815 6034 14875
rect 6115 14865 6315 14890
rect 6370 14881 6400 15069
rect 6344 14875 6400 14881
rect 6086 14815 6344 14835
rect 6396 14815 6400 14875
rect 6030 14805 6400 14815
rect 6430 15135 6800 15145
rect 6430 15075 6434 15135
rect 6486 15115 6744 15135
rect 6430 15069 6486 15075
rect 6430 14881 6460 15069
rect 6515 15060 6715 15085
rect 6796 15075 6800 15135
rect 6744 15069 6800 15075
rect 6515 15040 6585 15060
rect 6490 15000 6585 15040
rect 6645 15040 6715 15060
rect 6645 15000 6740 15040
rect 6490 14950 6740 15000
rect 6490 14910 6585 14950
rect 6515 14890 6585 14910
rect 6645 14910 6740 14950
rect 6645 14890 6715 14910
rect 6430 14875 6486 14881
rect 6430 14815 6434 14875
rect 6515 14865 6715 14890
rect 6770 14881 6800 15069
rect 6744 14875 6800 14881
rect 6486 14815 6744 14835
rect 6796 14815 6800 14875
rect 6430 14805 6800 14815
rect 6830 15135 7200 15145
rect 6830 15075 6834 15135
rect 6886 15115 7144 15135
rect 6830 15069 6886 15075
rect 6830 14881 6860 15069
rect 6915 15060 7115 15085
rect 7196 15075 7200 15135
rect 7144 15069 7200 15075
rect 6915 15040 6985 15060
rect 6890 15000 6985 15040
rect 7045 15040 7115 15060
rect 7045 15000 7140 15040
rect 6890 14950 7140 15000
rect 6890 14910 6985 14950
rect 6915 14890 6985 14910
rect 7045 14910 7140 14950
rect 7045 14890 7115 14910
rect 6830 14875 6886 14881
rect 6830 14815 6834 14875
rect 6915 14865 7115 14890
rect 7170 14881 7200 15069
rect 7144 14875 7200 14881
rect 6886 14815 7144 14835
rect 7196 14815 7200 14875
rect 6830 14805 7200 14815
rect 7230 15135 7600 15145
rect 7230 15075 7234 15135
rect 7286 15115 7544 15135
rect 7230 15069 7286 15075
rect 7230 14881 7260 15069
rect 7315 15060 7515 15085
rect 7596 15075 7600 15135
rect 7544 15069 7600 15075
rect 7315 15040 7385 15060
rect 7290 15000 7385 15040
rect 7445 15040 7515 15060
rect 7445 15000 7540 15040
rect 7290 14950 7540 15000
rect 7290 14910 7385 14950
rect 7315 14890 7385 14910
rect 7445 14910 7540 14950
rect 7445 14890 7515 14910
rect 7230 14875 7286 14881
rect 7230 14815 7234 14875
rect 7315 14865 7515 14890
rect 7570 14881 7600 15069
rect 7544 14875 7600 14881
rect 7286 14815 7544 14835
rect 7596 14815 7600 14875
rect 7230 14805 7600 14815
rect 7630 15135 8000 15145
rect 7630 15075 7634 15135
rect 7686 15115 7944 15135
rect 7630 15069 7686 15075
rect 7630 14881 7660 15069
rect 7715 15060 7915 15085
rect 7996 15075 8000 15135
rect 7944 15069 8000 15075
rect 7715 15040 7785 15060
rect 7690 15000 7785 15040
rect 7845 15040 7915 15060
rect 7845 15000 7940 15040
rect 7690 14950 7940 15000
rect 7690 14910 7785 14950
rect 7715 14890 7785 14910
rect 7845 14910 7940 14950
rect 7845 14890 7915 14910
rect 7630 14875 7686 14881
rect 7630 14815 7634 14875
rect 7715 14865 7915 14890
rect 7970 14881 8000 15069
rect 7944 14875 8000 14881
rect 7686 14815 7944 14835
rect 7996 14815 8000 14875
rect 7630 14805 8000 14815
rect 8030 15135 8400 15145
rect 8030 15075 8034 15135
rect 8086 15115 8344 15135
rect 8030 15069 8086 15075
rect 8030 14881 8060 15069
rect 8115 15060 8315 15085
rect 8396 15075 8400 15135
rect 8344 15069 8400 15075
rect 8115 15040 8185 15060
rect 8090 15000 8185 15040
rect 8245 15040 8315 15060
rect 8245 15000 8340 15040
rect 8090 14950 8340 15000
rect 8090 14910 8185 14950
rect 8115 14890 8185 14910
rect 8245 14910 8340 14950
rect 8245 14890 8315 14910
rect 8030 14875 8086 14881
rect 8030 14815 8034 14875
rect 8115 14865 8315 14890
rect 8370 14881 8400 15069
rect 8344 14875 8400 14881
rect 8086 14815 8344 14835
rect 8396 14815 8400 14875
rect 8030 14805 8400 14815
rect 8430 15135 8800 15145
rect 8430 15075 8434 15135
rect 8486 15115 8744 15135
rect 8430 15069 8486 15075
rect 8430 14881 8460 15069
rect 8515 15060 8715 15085
rect 8796 15075 8800 15135
rect 8744 15069 8800 15075
rect 8515 15040 8585 15060
rect 8490 15000 8585 15040
rect 8645 15040 8715 15060
rect 8645 15000 8740 15040
rect 8490 14950 8740 15000
rect 8490 14910 8585 14950
rect 8515 14890 8585 14910
rect 8645 14910 8740 14950
rect 8645 14890 8715 14910
rect 8430 14875 8486 14881
rect 8430 14815 8434 14875
rect 8515 14865 8715 14890
rect 8770 14881 8800 15069
rect 8744 14875 8800 14881
rect 8486 14815 8744 14835
rect 8796 14815 8800 14875
rect 8430 14805 8800 14815
rect 8830 15135 9200 15145
rect 8830 15075 8834 15135
rect 8886 15115 9144 15135
rect 8830 15069 8886 15075
rect 8830 14881 8860 15069
rect 8915 15060 9115 15085
rect 9196 15075 9200 15135
rect 9144 15069 9200 15075
rect 8915 15040 8985 15060
rect 8890 15000 8985 15040
rect 9045 15040 9115 15060
rect 9045 15000 9140 15040
rect 8890 14950 9140 15000
rect 8890 14910 8985 14950
rect 8915 14890 8985 14910
rect 9045 14910 9140 14950
rect 9045 14890 9115 14910
rect 8830 14875 8886 14881
rect 8830 14815 8834 14875
rect 8915 14865 9115 14890
rect 9170 14881 9200 15069
rect 9144 14875 9200 14881
rect 8886 14815 9144 14835
rect 9196 14815 9200 14875
rect 8830 14805 9200 14815
rect 9230 15135 9600 15145
rect 9230 15075 9234 15135
rect 9286 15115 9544 15135
rect 9230 15069 9286 15075
rect 9230 14881 9260 15069
rect 9315 15060 9515 15085
rect 9596 15075 9600 15135
rect 9544 15069 9600 15075
rect 9315 15040 9385 15060
rect 9290 15000 9385 15040
rect 9445 15040 9515 15060
rect 9445 15000 9540 15040
rect 9290 14950 9540 15000
rect 9290 14910 9385 14950
rect 9315 14890 9385 14910
rect 9445 14910 9540 14950
rect 9445 14890 9515 14910
rect 9230 14875 9286 14881
rect 9230 14815 9234 14875
rect 9315 14865 9515 14890
rect 9570 14881 9600 15069
rect 9544 14875 9600 14881
rect 9286 14815 9544 14835
rect 9596 14815 9600 14875
rect 9230 14805 9600 14815
rect 9630 15135 10000 15145
rect 9630 15075 9634 15135
rect 9686 15115 9944 15135
rect 9630 15069 9686 15075
rect 9630 14881 9660 15069
rect 9715 15060 9915 15085
rect 9996 15075 10000 15135
rect 9944 15069 10000 15075
rect 9715 15040 9785 15060
rect 9690 15000 9785 15040
rect 9845 15040 9915 15060
rect 9845 15000 9940 15040
rect 9690 14950 9940 15000
rect 9690 14910 9785 14950
rect 9715 14890 9785 14910
rect 9845 14910 9940 14950
rect 9845 14890 9915 14910
rect 9630 14875 9686 14881
rect 9630 14815 9634 14875
rect 9715 14865 9915 14890
rect 9970 14881 10000 15069
rect 9944 14875 10000 14881
rect 9686 14815 9944 14835
rect 9996 14815 10000 14875
rect 9630 14805 10000 14815
rect 10030 15135 10400 15145
rect 10030 15075 10034 15135
rect 10086 15115 10344 15135
rect 10030 15069 10086 15075
rect 10030 14881 10060 15069
rect 10115 15060 10315 15085
rect 10396 15075 10400 15135
rect 10344 15069 10400 15075
rect 10115 15040 10185 15060
rect 10090 15000 10185 15040
rect 10245 15040 10315 15060
rect 10245 15000 10340 15040
rect 10090 14950 10340 15000
rect 10090 14910 10185 14950
rect 10115 14890 10185 14910
rect 10245 14910 10340 14950
rect 10245 14890 10315 14910
rect 10030 14875 10086 14881
rect 10030 14815 10034 14875
rect 10115 14865 10315 14890
rect 10370 14881 10400 15069
rect 10344 14875 10400 14881
rect 10086 14815 10344 14835
rect 10396 14815 10400 14875
rect 10030 14805 10400 14815
rect 10430 15135 10800 15145
rect 10430 15075 10434 15135
rect 10486 15115 10744 15135
rect 10430 15069 10486 15075
rect 10430 14881 10460 15069
rect 10515 15060 10715 15085
rect 10796 15075 10800 15135
rect 10744 15069 10800 15075
rect 10515 15040 10585 15060
rect 10490 15000 10585 15040
rect 10645 15040 10715 15060
rect 10645 15000 10740 15040
rect 10490 14950 10740 15000
rect 10490 14910 10585 14950
rect 10515 14890 10585 14910
rect 10645 14910 10740 14950
rect 10645 14890 10715 14910
rect 10430 14875 10486 14881
rect 10430 14815 10434 14875
rect 10515 14865 10715 14890
rect 10770 14881 10800 15069
rect 10744 14875 10800 14881
rect 10486 14815 10744 14835
rect 10796 14815 10800 14875
rect 10430 14805 10800 14815
rect 10830 15135 11200 15145
rect 10830 15075 10834 15135
rect 10886 15115 11144 15135
rect 10830 15069 10886 15075
rect 10830 14881 10860 15069
rect 10915 15060 11115 15085
rect 11196 15075 11200 15135
rect 11144 15069 11200 15075
rect 10915 15040 10985 15060
rect 10890 15000 10985 15040
rect 11045 15040 11115 15060
rect 11045 15000 11140 15040
rect 10890 14950 11140 15000
rect 10890 14910 10985 14950
rect 10915 14890 10985 14910
rect 11045 14910 11140 14950
rect 11045 14890 11115 14910
rect 10830 14875 10886 14881
rect 10830 14815 10834 14875
rect 10915 14865 11115 14890
rect 11170 14881 11200 15069
rect 11144 14875 11200 14881
rect 10886 14815 11144 14835
rect 11196 14815 11200 14875
rect 10830 14805 11200 14815
rect 11230 15135 11600 15145
rect 11230 15075 11234 15135
rect 11286 15115 11544 15135
rect 11230 15069 11286 15075
rect 11230 14881 11260 15069
rect 11315 15060 11515 15085
rect 11596 15075 11600 15135
rect 11544 15069 11600 15075
rect 11315 15040 11385 15060
rect 11290 15000 11385 15040
rect 11445 15040 11515 15060
rect 11445 15000 11540 15040
rect 11290 14950 11540 15000
rect 11290 14910 11385 14950
rect 11315 14890 11385 14910
rect 11445 14910 11540 14950
rect 11445 14890 11515 14910
rect 11230 14875 11286 14881
rect 11230 14815 11234 14875
rect 11315 14865 11515 14890
rect 11570 14881 11600 15069
rect 11544 14875 11600 14881
rect 11286 14815 11544 14835
rect 11596 14815 11600 14875
rect 11230 14805 11600 14815
rect 11630 15135 12000 15145
rect 11630 15075 11634 15135
rect 11686 15115 11944 15135
rect 11630 15069 11686 15075
rect 11630 14881 11660 15069
rect 11715 15060 11915 15085
rect 11996 15075 12000 15135
rect 11944 15069 12000 15075
rect 11715 15040 11785 15060
rect 11690 15000 11785 15040
rect 11845 15040 11915 15060
rect 11845 15000 11940 15040
rect 11690 14950 11940 15000
rect 11690 14910 11785 14950
rect 11715 14890 11785 14910
rect 11845 14910 11940 14950
rect 11845 14890 11915 14910
rect 11630 14875 11686 14881
rect 11630 14815 11634 14875
rect 11715 14865 11915 14890
rect 11970 14881 12000 15069
rect 11944 14875 12000 14881
rect 11686 14815 11944 14835
rect 11996 14815 12000 14875
rect 11630 14805 12000 14815
rect 12030 15135 12400 15145
rect 12030 15075 12034 15135
rect 12086 15115 12344 15135
rect 12030 15069 12086 15075
rect 12030 14881 12060 15069
rect 12115 15060 12315 15085
rect 12396 15075 12400 15135
rect 12344 15069 12400 15075
rect 12115 15040 12185 15060
rect 12090 15000 12185 15040
rect 12245 15040 12315 15060
rect 12245 15000 12340 15040
rect 12090 14950 12340 15000
rect 12090 14910 12185 14950
rect 12115 14890 12185 14910
rect 12245 14910 12340 14950
rect 12245 14890 12315 14910
rect 12030 14875 12086 14881
rect 12030 14815 12034 14875
rect 12115 14865 12315 14890
rect 12370 14881 12400 15069
rect 12344 14875 12400 14881
rect 12086 14815 12344 14835
rect 12396 14815 12400 14875
rect 12030 14805 12400 14815
rect 12430 15135 12800 15145
rect 12430 15075 12434 15135
rect 12486 15115 12744 15135
rect 12430 15069 12486 15075
rect 12430 14881 12460 15069
rect 12515 15060 12715 15085
rect 12796 15075 12800 15135
rect 12744 15069 12800 15075
rect 12515 15040 12585 15060
rect 12490 15000 12585 15040
rect 12645 15040 12715 15060
rect 12645 15000 12740 15040
rect 12490 14950 12740 15000
rect 12490 14910 12585 14950
rect 12515 14890 12585 14910
rect 12645 14910 12740 14950
rect 12645 14890 12715 14910
rect 12430 14875 12486 14881
rect 12430 14815 12434 14875
rect 12515 14865 12715 14890
rect 12770 14881 12800 15069
rect 12744 14875 12800 14881
rect 12486 14815 12744 14835
rect 12796 14815 12800 14875
rect 12430 14805 12800 14815
rect 12830 15135 13200 15145
rect 12830 15075 12834 15135
rect 12886 15115 13144 15135
rect 12830 15069 12886 15075
rect 12830 14881 12860 15069
rect 12915 15060 13115 15085
rect 13196 15075 13200 15135
rect 13144 15069 13200 15075
rect 12915 15040 12985 15060
rect 12890 15000 12985 15040
rect 13045 15040 13115 15060
rect 13045 15000 13140 15040
rect 12890 14950 13140 15000
rect 12890 14910 12985 14950
rect 12915 14890 12985 14910
rect 13045 14910 13140 14950
rect 13045 14890 13115 14910
rect 12830 14875 12886 14881
rect 12830 14815 12834 14875
rect 12915 14865 13115 14890
rect 13170 14881 13200 15069
rect 13144 14875 13200 14881
rect 12886 14815 13144 14835
rect 13196 14815 13200 14875
rect 12830 14805 13200 14815
rect -370 14765 0 14775
rect -370 14705 -366 14765
rect -314 14745 -56 14765
rect -370 14699 -314 14705
rect -370 14511 -340 14699
rect -285 14690 -85 14715
rect -4 14705 0 14765
rect -56 14699 0 14705
rect -285 14670 -215 14690
rect -310 14630 -215 14670
rect -155 14670 -85 14690
rect -155 14630 -60 14670
rect -310 14580 -60 14630
rect -310 14540 -215 14580
rect -285 14520 -215 14540
rect -155 14540 -60 14580
rect -155 14520 -85 14540
rect -370 14505 -314 14511
rect -370 14445 -366 14505
rect -285 14495 -85 14520
rect -30 14511 0 14699
rect -56 14505 0 14511
rect -314 14445 -56 14465
rect -4 14445 0 14505
rect -370 14435 0 14445
rect 30 14765 400 14775
rect 30 14705 34 14765
rect 86 14745 344 14765
rect 30 14699 86 14705
rect 30 14511 60 14699
rect 115 14690 315 14715
rect 396 14705 400 14765
rect 344 14699 400 14705
rect 115 14670 185 14690
rect 90 14630 185 14670
rect 245 14670 315 14690
rect 245 14630 340 14670
rect 90 14580 340 14630
rect 90 14540 185 14580
rect 115 14520 185 14540
rect 245 14540 340 14580
rect 245 14520 315 14540
rect 30 14505 86 14511
rect 30 14445 34 14505
rect 115 14495 315 14520
rect 370 14511 400 14699
rect 344 14505 400 14511
rect 86 14445 344 14465
rect 396 14445 400 14505
rect 30 14435 400 14445
rect 430 14765 800 14775
rect 430 14705 434 14765
rect 486 14745 744 14765
rect 430 14699 486 14705
rect 430 14511 460 14699
rect 515 14690 715 14715
rect 796 14705 800 14765
rect 744 14699 800 14705
rect 515 14670 585 14690
rect 490 14630 585 14670
rect 645 14670 715 14690
rect 645 14630 740 14670
rect 490 14580 740 14630
rect 490 14540 585 14580
rect 515 14520 585 14540
rect 645 14540 740 14580
rect 645 14520 715 14540
rect 430 14505 486 14511
rect 430 14445 434 14505
rect 515 14495 715 14520
rect 770 14511 800 14699
rect 744 14505 800 14511
rect 486 14445 744 14465
rect 796 14445 800 14505
rect 430 14435 800 14445
rect 830 14765 1200 14775
rect 830 14705 834 14765
rect 886 14745 1144 14765
rect 830 14699 886 14705
rect 830 14511 860 14699
rect 915 14690 1115 14715
rect 1196 14705 1200 14765
rect 1144 14699 1200 14705
rect 915 14670 985 14690
rect 890 14630 985 14670
rect 1045 14670 1115 14690
rect 1045 14630 1140 14670
rect 890 14580 1140 14630
rect 890 14540 985 14580
rect 915 14520 985 14540
rect 1045 14540 1140 14580
rect 1045 14520 1115 14540
rect 830 14505 886 14511
rect 830 14445 834 14505
rect 915 14495 1115 14520
rect 1170 14511 1200 14699
rect 1144 14505 1200 14511
rect 886 14445 1144 14465
rect 1196 14445 1200 14505
rect 830 14435 1200 14445
rect 1230 14765 1600 14775
rect 1230 14705 1234 14765
rect 1286 14745 1544 14765
rect 1230 14699 1286 14705
rect 1230 14511 1260 14699
rect 1315 14690 1515 14715
rect 1596 14705 1600 14765
rect 1544 14699 1600 14705
rect 1315 14670 1385 14690
rect 1290 14630 1385 14670
rect 1445 14670 1515 14690
rect 1445 14630 1540 14670
rect 1290 14580 1540 14630
rect 1290 14540 1385 14580
rect 1315 14520 1385 14540
rect 1445 14540 1540 14580
rect 1445 14520 1515 14540
rect 1230 14505 1286 14511
rect 1230 14445 1234 14505
rect 1315 14495 1515 14520
rect 1570 14511 1600 14699
rect 1544 14505 1600 14511
rect 1286 14445 1544 14465
rect 1596 14445 1600 14505
rect 1230 14435 1600 14445
rect 1630 14765 2000 14775
rect 1630 14705 1634 14765
rect 1686 14745 1944 14765
rect 1630 14699 1686 14705
rect 1630 14511 1660 14699
rect 1715 14690 1915 14715
rect 1996 14705 2000 14765
rect 1944 14699 2000 14705
rect 1715 14670 1785 14690
rect 1690 14630 1785 14670
rect 1845 14670 1915 14690
rect 1845 14630 1940 14670
rect 1690 14580 1940 14630
rect 1690 14540 1785 14580
rect 1715 14520 1785 14540
rect 1845 14540 1940 14580
rect 1845 14520 1915 14540
rect 1630 14505 1686 14511
rect 1630 14445 1634 14505
rect 1715 14495 1915 14520
rect 1970 14511 2000 14699
rect 1944 14505 2000 14511
rect 1686 14445 1944 14465
rect 1996 14445 2000 14505
rect 1630 14435 2000 14445
rect 2030 14765 2400 14775
rect 2030 14705 2034 14765
rect 2086 14745 2344 14765
rect 2030 14699 2086 14705
rect 2030 14511 2060 14699
rect 2115 14690 2315 14715
rect 2396 14705 2400 14765
rect 2344 14699 2400 14705
rect 2115 14670 2185 14690
rect 2090 14630 2185 14670
rect 2245 14670 2315 14690
rect 2245 14630 2340 14670
rect 2090 14580 2340 14630
rect 2090 14540 2185 14580
rect 2115 14520 2185 14540
rect 2245 14540 2340 14580
rect 2245 14520 2315 14540
rect 2030 14505 2086 14511
rect 2030 14445 2034 14505
rect 2115 14495 2315 14520
rect 2370 14511 2400 14699
rect 2344 14505 2400 14511
rect 2086 14445 2344 14465
rect 2396 14445 2400 14505
rect 2030 14435 2400 14445
rect 2430 14765 2800 14775
rect 2430 14705 2434 14765
rect 2486 14745 2744 14765
rect 2430 14699 2486 14705
rect 2430 14511 2460 14699
rect 2515 14690 2715 14715
rect 2796 14705 2800 14765
rect 2744 14699 2800 14705
rect 2515 14670 2585 14690
rect 2490 14630 2585 14670
rect 2645 14670 2715 14690
rect 2645 14630 2740 14670
rect 2490 14580 2740 14630
rect 2490 14540 2585 14580
rect 2515 14520 2585 14540
rect 2645 14540 2740 14580
rect 2645 14520 2715 14540
rect 2430 14505 2486 14511
rect 2430 14445 2434 14505
rect 2515 14495 2715 14520
rect 2770 14511 2800 14699
rect 2744 14505 2800 14511
rect 2486 14445 2744 14465
rect 2796 14445 2800 14505
rect 2430 14435 2800 14445
rect 2830 14765 3200 14775
rect 2830 14705 2834 14765
rect 2886 14745 3144 14765
rect 2830 14699 2886 14705
rect 2830 14511 2860 14699
rect 2915 14690 3115 14715
rect 3196 14705 3200 14765
rect 3144 14699 3200 14705
rect 2915 14670 2985 14690
rect 2890 14630 2985 14670
rect 3045 14670 3115 14690
rect 3045 14630 3140 14670
rect 2890 14580 3140 14630
rect 2890 14540 2985 14580
rect 2915 14520 2985 14540
rect 3045 14540 3140 14580
rect 3045 14520 3115 14540
rect 2830 14505 2886 14511
rect 2830 14445 2834 14505
rect 2915 14495 3115 14520
rect 3170 14511 3200 14699
rect 3144 14505 3200 14511
rect 2886 14445 3144 14465
rect 3196 14445 3200 14505
rect 2830 14435 3200 14445
rect 3230 14765 3600 14775
rect 3230 14705 3234 14765
rect 3286 14745 3544 14765
rect 3230 14699 3286 14705
rect 3230 14511 3260 14699
rect 3315 14690 3515 14715
rect 3596 14705 3600 14765
rect 3544 14699 3600 14705
rect 3315 14670 3385 14690
rect 3290 14630 3385 14670
rect 3445 14670 3515 14690
rect 3445 14630 3540 14670
rect 3290 14580 3540 14630
rect 3290 14540 3385 14580
rect 3315 14520 3385 14540
rect 3445 14540 3540 14580
rect 3445 14520 3515 14540
rect 3230 14505 3286 14511
rect 3230 14445 3234 14505
rect 3315 14495 3515 14520
rect 3570 14511 3600 14699
rect 3544 14505 3600 14511
rect 3286 14445 3544 14465
rect 3596 14445 3600 14505
rect 3230 14435 3600 14445
rect 3630 14765 4000 14775
rect 3630 14705 3634 14765
rect 3686 14745 3944 14765
rect 3630 14699 3686 14705
rect 3630 14511 3660 14699
rect 3715 14690 3915 14715
rect 3996 14705 4000 14765
rect 3944 14699 4000 14705
rect 3715 14670 3785 14690
rect 3690 14630 3785 14670
rect 3845 14670 3915 14690
rect 3845 14630 3940 14670
rect 3690 14580 3940 14630
rect 3690 14540 3785 14580
rect 3715 14520 3785 14540
rect 3845 14540 3940 14580
rect 3845 14520 3915 14540
rect 3630 14505 3686 14511
rect 3630 14445 3634 14505
rect 3715 14495 3915 14520
rect 3970 14511 4000 14699
rect 3944 14505 4000 14511
rect 3686 14445 3944 14465
rect 3996 14445 4000 14505
rect 3630 14435 4000 14445
rect 4030 14765 4400 14775
rect 4030 14705 4034 14765
rect 4086 14745 4344 14765
rect 4030 14699 4086 14705
rect 4030 14511 4060 14699
rect 4115 14690 4315 14715
rect 4396 14705 4400 14765
rect 4344 14699 4400 14705
rect 4115 14670 4185 14690
rect 4090 14630 4185 14670
rect 4245 14670 4315 14690
rect 4245 14630 4340 14670
rect 4090 14580 4340 14630
rect 4090 14540 4185 14580
rect 4115 14520 4185 14540
rect 4245 14540 4340 14580
rect 4245 14520 4315 14540
rect 4030 14505 4086 14511
rect 4030 14445 4034 14505
rect 4115 14495 4315 14520
rect 4370 14511 4400 14699
rect 4344 14505 4400 14511
rect 4086 14445 4344 14465
rect 4396 14445 4400 14505
rect 4030 14435 4400 14445
rect 4430 14765 4800 14775
rect 4430 14705 4434 14765
rect 4486 14745 4744 14765
rect 4430 14699 4486 14705
rect 4430 14511 4460 14699
rect 4515 14690 4715 14715
rect 4796 14705 4800 14765
rect 4744 14699 4800 14705
rect 4515 14670 4585 14690
rect 4490 14630 4585 14670
rect 4645 14670 4715 14690
rect 4645 14630 4740 14670
rect 4490 14580 4740 14630
rect 4490 14540 4585 14580
rect 4515 14520 4585 14540
rect 4645 14540 4740 14580
rect 4645 14520 4715 14540
rect 4430 14505 4486 14511
rect 4430 14445 4434 14505
rect 4515 14495 4715 14520
rect 4770 14511 4800 14699
rect 4744 14505 4800 14511
rect 4486 14445 4744 14465
rect 4796 14445 4800 14505
rect 4430 14435 4800 14445
rect 4830 14765 5200 14775
rect 4830 14705 4834 14765
rect 4886 14745 5144 14765
rect 4830 14699 4886 14705
rect 4830 14511 4860 14699
rect 4915 14690 5115 14715
rect 5196 14705 5200 14765
rect 5144 14699 5200 14705
rect 4915 14670 4985 14690
rect 4890 14630 4985 14670
rect 5045 14670 5115 14690
rect 5045 14630 5140 14670
rect 4890 14580 5140 14630
rect 4890 14540 4985 14580
rect 4915 14520 4985 14540
rect 5045 14540 5140 14580
rect 5045 14520 5115 14540
rect 4830 14505 4886 14511
rect 4830 14445 4834 14505
rect 4915 14495 5115 14520
rect 5170 14511 5200 14699
rect 5144 14505 5200 14511
rect 4886 14445 5144 14465
rect 5196 14445 5200 14505
rect 4830 14435 5200 14445
rect 5230 14765 5600 14775
rect 5230 14705 5234 14765
rect 5286 14745 5544 14765
rect 5230 14699 5286 14705
rect 5230 14511 5260 14699
rect 5315 14690 5515 14715
rect 5596 14705 5600 14765
rect 5544 14699 5600 14705
rect 5315 14670 5385 14690
rect 5290 14630 5385 14670
rect 5445 14670 5515 14690
rect 5445 14630 5540 14670
rect 5290 14580 5540 14630
rect 5290 14540 5385 14580
rect 5315 14520 5385 14540
rect 5445 14540 5540 14580
rect 5445 14520 5515 14540
rect 5230 14505 5286 14511
rect 5230 14445 5234 14505
rect 5315 14495 5515 14520
rect 5570 14511 5600 14699
rect 5544 14505 5600 14511
rect 5286 14445 5544 14465
rect 5596 14445 5600 14505
rect 5230 14435 5600 14445
rect 5630 14765 6000 14775
rect 5630 14705 5634 14765
rect 5686 14745 5944 14765
rect 5630 14699 5686 14705
rect 5630 14511 5660 14699
rect 5715 14690 5915 14715
rect 5996 14705 6000 14765
rect 5944 14699 6000 14705
rect 5715 14670 5785 14690
rect 5690 14630 5785 14670
rect 5845 14670 5915 14690
rect 5845 14630 5940 14670
rect 5690 14580 5940 14630
rect 5690 14540 5785 14580
rect 5715 14520 5785 14540
rect 5845 14540 5940 14580
rect 5845 14520 5915 14540
rect 5630 14505 5686 14511
rect 5630 14445 5634 14505
rect 5715 14495 5915 14520
rect 5970 14511 6000 14699
rect 5944 14505 6000 14511
rect 5686 14445 5944 14465
rect 5996 14445 6000 14505
rect 5630 14435 6000 14445
rect 6030 14765 6400 14775
rect 6030 14705 6034 14765
rect 6086 14745 6344 14765
rect 6030 14699 6086 14705
rect 6030 14511 6060 14699
rect 6115 14690 6315 14715
rect 6396 14705 6400 14765
rect 6344 14699 6400 14705
rect 6115 14670 6185 14690
rect 6090 14630 6185 14670
rect 6245 14670 6315 14690
rect 6245 14630 6340 14670
rect 6090 14580 6340 14630
rect 6090 14540 6185 14580
rect 6115 14520 6185 14540
rect 6245 14540 6340 14580
rect 6245 14520 6315 14540
rect 6030 14505 6086 14511
rect 6030 14445 6034 14505
rect 6115 14495 6315 14520
rect 6370 14511 6400 14699
rect 6344 14505 6400 14511
rect 6086 14445 6344 14465
rect 6396 14445 6400 14505
rect 6030 14435 6400 14445
rect 6430 14765 6800 14775
rect 6430 14705 6434 14765
rect 6486 14745 6744 14765
rect 6430 14699 6486 14705
rect 6430 14511 6460 14699
rect 6515 14690 6715 14715
rect 6796 14705 6800 14765
rect 6744 14699 6800 14705
rect 6515 14670 6585 14690
rect 6490 14630 6585 14670
rect 6645 14670 6715 14690
rect 6645 14630 6740 14670
rect 6490 14580 6740 14630
rect 6490 14540 6585 14580
rect 6515 14520 6585 14540
rect 6645 14540 6740 14580
rect 6645 14520 6715 14540
rect 6430 14505 6486 14511
rect 6430 14445 6434 14505
rect 6515 14495 6715 14520
rect 6770 14511 6800 14699
rect 6744 14505 6800 14511
rect 6486 14445 6744 14465
rect 6796 14445 6800 14505
rect 6430 14435 6800 14445
rect 6830 14765 7200 14775
rect 6830 14705 6834 14765
rect 6886 14745 7144 14765
rect 6830 14699 6886 14705
rect 6830 14511 6860 14699
rect 6915 14690 7115 14715
rect 7196 14705 7200 14765
rect 7144 14699 7200 14705
rect 6915 14670 6985 14690
rect 6890 14630 6985 14670
rect 7045 14670 7115 14690
rect 7045 14630 7140 14670
rect 6890 14580 7140 14630
rect 6890 14540 6985 14580
rect 6915 14520 6985 14540
rect 7045 14540 7140 14580
rect 7045 14520 7115 14540
rect 6830 14505 6886 14511
rect 6830 14445 6834 14505
rect 6915 14495 7115 14520
rect 7170 14511 7200 14699
rect 7144 14505 7200 14511
rect 6886 14445 7144 14465
rect 7196 14445 7200 14505
rect 6830 14435 7200 14445
rect 7230 14765 7600 14775
rect 7230 14705 7234 14765
rect 7286 14745 7544 14765
rect 7230 14699 7286 14705
rect 7230 14511 7260 14699
rect 7315 14690 7515 14715
rect 7596 14705 7600 14765
rect 7544 14699 7600 14705
rect 7315 14670 7385 14690
rect 7290 14630 7385 14670
rect 7445 14670 7515 14690
rect 7445 14630 7540 14670
rect 7290 14580 7540 14630
rect 7290 14540 7385 14580
rect 7315 14520 7385 14540
rect 7445 14540 7540 14580
rect 7445 14520 7515 14540
rect 7230 14505 7286 14511
rect 7230 14445 7234 14505
rect 7315 14495 7515 14520
rect 7570 14511 7600 14699
rect 7544 14505 7600 14511
rect 7286 14445 7544 14465
rect 7596 14445 7600 14505
rect 7230 14435 7600 14445
rect 7630 14765 8000 14775
rect 7630 14705 7634 14765
rect 7686 14745 7944 14765
rect 7630 14699 7686 14705
rect 7630 14511 7660 14699
rect 7715 14690 7915 14715
rect 7996 14705 8000 14765
rect 7944 14699 8000 14705
rect 7715 14670 7785 14690
rect 7690 14630 7785 14670
rect 7845 14670 7915 14690
rect 7845 14630 7940 14670
rect 7690 14580 7940 14630
rect 7690 14540 7785 14580
rect 7715 14520 7785 14540
rect 7845 14540 7940 14580
rect 7845 14520 7915 14540
rect 7630 14505 7686 14511
rect 7630 14445 7634 14505
rect 7715 14495 7915 14520
rect 7970 14511 8000 14699
rect 7944 14505 8000 14511
rect 7686 14445 7944 14465
rect 7996 14445 8000 14505
rect 7630 14435 8000 14445
rect 8030 14765 8400 14775
rect 8030 14705 8034 14765
rect 8086 14745 8344 14765
rect 8030 14699 8086 14705
rect 8030 14511 8060 14699
rect 8115 14690 8315 14715
rect 8396 14705 8400 14765
rect 8344 14699 8400 14705
rect 8115 14670 8185 14690
rect 8090 14630 8185 14670
rect 8245 14670 8315 14690
rect 8245 14630 8340 14670
rect 8090 14580 8340 14630
rect 8090 14540 8185 14580
rect 8115 14520 8185 14540
rect 8245 14540 8340 14580
rect 8245 14520 8315 14540
rect 8030 14505 8086 14511
rect 8030 14445 8034 14505
rect 8115 14495 8315 14520
rect 8370 14511 8400 14699
rect 8344 14505 8400 14511
rect 8086 14445 8344 14465
rect 8396 14445 8400 14505
rect 8030 14435 8400 14445
rect 8430 14765 8800 14775
rect 8430 14705 8434 14765
rect 8486 14745 8744 14765
rect 8430 14699 8486 14705
rect 8430 14511 8460 14699
rect 8515 14690 8715 14715
rect 8796 14705 8800 14765
rect 8744 14699 8800 14705
rect 8515 14670 8585 14690
rect 8490 14630 8585 14670
rect 8645 14670 8715 14690
rect 8645 14630 8740 14670
rect 8490 14580 8740 14630
rect 8490 14540 8585 14580
rect 8515 14520 8585 14540
rect 8645 14540 8740 14580
rect 8645 14520 8715 14540
rect 8430 14505 8486 14511
rect 8430 14445 8434 14505
rect 8515 14495 8715 14520
rect 8770 14511 8800 14699
rect 8744 14505 8800 14511
rect 8486 14445 8744 14465
rect 8796 14445 8800 14505
rect 8430 14435 8800 14445
rect 8830 14765 9200 14775
rect 8830 14705 8834 14765
rect 8886 14745 9144 14765
rect 8830 14699 8886 14705
rect 8830 14511 8860 14699
rect 8915 14690 9115 14715
rect 9196 14705 9200 14765
rect 9144 14699 9200 14705
rect 8915 14670 8985 14690
rect 8890 14630 8985 14670
rect 9045 14670 9115 14690
rect 9045 14630 9140 14670
rect 8890 14580 9140 14630
rect 8890 14540 8985 14580
rect 8915 14520 8985 14540
rect 9045 14540 9140 14580
rect 9045 14520 9115 14540
rect 8830 14505 8886 14511
rect 8830 14445 8834 14505
rect 8915 14495 9115 14520
rect 9170 14511 9200 14699
rect 9144 14505 9200 14511
rect 8886 14445 9144 14465
rect 9196 14445 9200 14505
rect 8830 14435 9200 14445
rect 9230 14765 9600 14775
rect 9230 14705 9234 14765
rect 9286 14745 9544 14765
rect 9230 14699 9286 14705
rect 9230 14511 9260 14699
rect 9315 14690 9515 14715
rect 9596 14705 9600 14765
rect 9544 14699 9600 14705
rect 9315 14670 9385 14690
rect 9290 14630 9385 14670
rect 9445 14670 9515 14690
rect 9445 14630 9540 14670
rect 9290 14580 9540 14630
rect 9290 14540 9385 14580
rect 9315 14520 9385 14540
rect 9445 14540 9540 14580
rect 9445 14520 9515 14540
rect 9230 14505 9286 14511
rect 9230 14445 9234 14505
rect 9315 14495 9515 14520
rect 9570 14511 9600 14699
rect 9544 14505 9600 14511
rect 9286 14445 9544 14465
rect 9596 14445 9600 14505
rect 9230 14435 9600 14445
rect 9630 14765 10000 14775
rect 9630 14705 9634 14765
rect 9686 14745 9944 14765
rect 9630 14699 9686 14705
rect 9630 14511 9660 14699
rect 9715 14690 9915 14715
rect 9996 14705 10000 14765
rect 9944 14699 10000 14705
rect 9715 14670 9785 14690
rect 9690 14630 9785 14670
rect 9845 14670 9915 14690
rect 9845 14630 9940 14670
rect 9690 14580 9940 14630
rect 9690 14540 9785 14580
rect 9715 14520 9785 14540
rect 9845 14540 9940 14580
rect 9845 14520 9915 14540
rect 9630 14505 9686 14511
rect 9630 14445 9634 14505
rect 9715 14495 9915 14520
rect 9970 14511 10000 14699
rect 9944 14505 10000 14511
rect 9686 14445 9944 14465
rect 9996 14445 10000 14505
rect 9630 14435 10000 14445
rect 10030 14765 10400 14775
rect 10030 14705 10034 14765
rect 10086 14745 10344 14765
rect 10030 14699 10086 14705
rect 10030 14511 10060 14699
rect 10115 14690 10315 14715
rect 10396 14705 10400 14765
rect 10344 14699 10400 14705
rect 10115 14670 10185 14690
rect 10090 14630 10185 14670
rect 10245 14670 10315 14690
rect 10245 14630 10340 14670
rect 10090 14580 10340 14630
rect 10090 14540 10185 14580
rect 10115 14520 10185 14540
rect 10245 14540 10340 14580
rect 10245 14520 10315 14540
rect 10030 14505 10086 14511
rect 10030 14445 10034 14505
rect 10115 14495 10315 14520
rect 10370 14511 10400 14699
rect 10344 14505 10400 14511
rect 10086 14445 10344 14465
rect 10396 14445 10400 14505
rect 10030 14435 10400 14445
rect 10430 14765 10800 14775
rect 10430 14705 10434 14765
rect 10486 14745 10744 14765
rect 10430 14699 10486 14705
rect 10430 14511 10460 14699
rect 10515 14690 10715 14715
rect 10796 14705 10800 14765
rect 10744 14699 10800 14705
rect 10515 14670 10585 14690
rect 10490 14630 10585 14670
rect 10645 14670 10715 14690
rect 10645 14630 10740 14670
rect 10490 14580 10740 14630
rect 10490 14540 10585 14580
rect 10515 14520 10585 14540
rect 10645 14540 10740 14580
rect 10645 14520 10715 14540
rect 10430 14505 10486 14511
rect 10430 14445 10434 14505
rect 10515 14495 10715 14520
rect 10770 14511 10800 14699
rect 10744 14505 10800 14511
rect 10486 14445 10744 14465
rect 10796 14445 10800 14505
rect 10430 14435 10800 14445
rect 10830 14765 11200 14775
rect 10830 14705 10834 14765
rect 10886 14745 11144 14765
rect 10830 14699 10886 14705
rect 10830 14511 10860 14699
rect 10915 14690 11115 14715
rect 11196 14705 11200 14765
rect 11144 14699 11200 14705
rect 10915 14670 10985 14690
rect 10890 14630 10985 14670
rect 11045 14670 11115 14690
rect 11045 14630 11140 14670
rect 10890 14580 11140 14630
rect 10890 14540 10985 14580
rect 10915 14520 10985 14540
rect 11045 14540 11140 14580
rect 11045 14520 11115 14540
rect 10830 14505 10886 14511
rect 10830 14445 10834 14505
rect 10915 14495 11115 14520
rect 11170 14511 11200 14699
rect 11144 14505 11200 14511
rect 10886 14445 11144 14465
rect 11196 14445 11200 14505
rect 10830 14435 11200 14445
rect 11230 14765 11600 14775
rect 11230 14705 11234 14765
rect 11286 14745 11544 14765
rect 11230 14699 11286 14705
rect 11230 14511 11260 14699
rect 11315 14690 11515 14715
rect 11596 14705 11600 14765
rect 11544 14699 11600 14705
rect 11315 14670 11385 14690
rect 11290 14630 11385 14670
rect 11445 14670 11515 14690
rect 11445 14630 11540 14670
rect 11290 14580 11540 14630
rect 11290 14540 11385 14580
rect 11315 14520 11385 14540
rect 11445 14540 11540 14580
rect 11445 14520 11515 14540
rect 11230 14505 11286 14511
rect 11230 14445 11234 14505
rect 11315 14495 11515 14520
rect 11570 14511 11600 14699
rect 11544 14505 11600 14511
rect 11286 14445 11544 14465
rect 11596 14445 11600 14505
rect 11230 14435 11600 14445
rect 11630 14765 12000 14775
rect 11630 14705 11634 14765
rect 11686 14745 11944 14765
rect 11630 14699 11686 14705
rect 11630 14511 11660 14699
rect 11715 14690 11915 14715
rect 11996 14705 12000 14765
rect 11944 14699 12000 14705
rect 11715 14670 11785 14690
rect 11690 14630 11785 14670
rect 11845 14670 11915 14690
rect 11845 14630 11940 14670
rect 11690 14580 11940 14630
rect 11690 14540 11785 14580
rect 11715 14520 11785 14540
rect 11845 14540 11940 14580
rect 11845 14520 11915 14540
rect 11630 14505 11686 14511
rect 11630 14445 11634 14505
rect 11715 14495 11915 14520
rect 11970 14511 12000 14699
rect 11944 14505 12000 14511
rect 11686 14445 11944 14465
rect 11996 14445 12000 14505
rect 11630 14435 12000 14445
rect 12030 14765 12400 14775
rect 12030 14705 12034 14765
rect 12086 14745 12344 14765
rect 12030 14699 12086 14705
rect 12030 14511 12060 14699
rect 12115 14690 12315 14715
rect 12396 14705 12400 14765
rect 12344 14699 12400 14705
rect 12115 14670 12185 14690
rect 12090 14630 12185 14670
rect 12245 14670 12315 14690
rect 12245 14630 12340 14670
rect 12090 14580 12340 14630
rect 12090 14540 12185 14580
rect 12115 14520 12185 14540
rect 12245 14540 12340 14580
rect 12245 14520 12315 14540
rect 12030 14505 12086 14511
rect 12030 14445 12034 14505
rect 12115 14495 12315 14520
rect 12370 14511 12400 14699
rect 12344 14505 12400 14511
rect 12086 14445 12344 14465
rect 12396 14445 12400 14505
rect 12030 14435 12400 14445
rect 12430 14765 12800 14775
rect 12430 14705 12434 14765
rect 12486 14745 12744 14765
rect 12430 14699 12486 14705
rect 12430 14511 12460 14699
rect 12515 14690 12715 14715
rect 12796 14705 12800 14765
rect 12744 14699 12800 14705
rect 12515 14670 12585 14690
rect 12490 14630 12585 14670
rect 12645 14670 12715 14690
rect 12645 14630 12740 14670
rect 12490 14580 12740 14630
rect 12490 14540 12585 14580
rect 12515 14520 12585 14540
rect 12645 14540 12740 14580
rect 12645 14520 12715 14540
rect 12430 14505 12486 14511
rect 12430 14445 12434 14505
rect 12515 14495 12715 14520
rect 12770 14511 12800 14699
rect 12744 14505 12800 14511
rect 12486 14445 12744 14465
rect 12796 14445 12800 14505
rect 12430 14435 12800 14445
rect 12830 14765 13200 14775
rect 12830 14705 12834 14765
rect 12886 14745 13144 14765
rect 12830 14699 12886 14705
rect 12830 14511 12860 14699
rect 12915 14690 13115 14715
rect 13196 14705 13200 14765
rect 13144 14699 13200 14705
rect 12915 14670 12985 14690
rect 12890 14630 12985 14670
rect 13045 14670 13115 14690
rect 13045 14630 13140 14670
rect 12890 14580 13140 14630
rect 12890 14540 12985 14580
rect 12915 14520 12985 14540
rect 13045 14540 13140 14580
rect 13045 14520 13115 14540
rect 12830 14505 12886 14511
rect 12830 14445 12834 14505
rect 12915 14495 13115 14520
rect 13170 14511 13200 14699
rect 13144 14505 13200 14511
rect 12886 14445 13144 14465
rect 13196 14445 13200 14505
rect 12830 14435 13200 14445
rect -370 14395 0 14405
rect -370 14335 -366 14395
rect -314 14375 -56 14395
rect -370 14329 -314 14335
rect -370 14141 -340 14329
rect -285 14320 -85 14345
rect -4 14335 0 14395
rect -56 14329 0 14335
rect -285 14300 -215 14320
rect -310 14260 -215 14300
rect -155 14300 -85 14320
rect -155 14260 -60 14300
rect -310 14210 -60 14260
rect -310 14170 -215 14210
rect -285 14150 -215 14170
rect -155 14170 -60 14210
rect -155 14150 -85 14170
rect -370 14135 -314 14141
rect -370 14075 -366 14135
rect -285 14125 -85 14150
rect -30 14141 0 14329
rect -56 14135 0 14141
rect -314 14075 -56 14095
rect -4 14075 0 14135
rect -370 14065 0 14075
rect 30 14395 400 14405
rect 30 14335 34 14395
rect 86 14375 344 14395
rect 30 14329 86 14335
rect 30 14141 60 14329
rect 115 14320 315 14345
rect 396 14335 400 14395
rect 344 14329 400 14335
rect 115 14300 185 14320
rect 90 14260 185 14300
rect 245 14300 315 14320
rect 245 14260 340 14300
rect 90 14210 340 14260
rect 90 14170 185 14210
rect 115 14150 185 14170
rect 245 14170 340 14210
rect 245 14150 315 14170
rect 30 14135 86 14141
rect 30 14075 34 14135
rect 115 14125 315 14150
rect 370 14141 400 14329
rect 344 14135 400 14141
rect 86 14075 344 14095
rect 396 14075 400 14135
rect 30 14065 400 14075
rect 430 14395 800 14405
rect 430 14335 434 14395
rect 486 14375 744 14395
rect 430 14329 486 14335
rect 430 14141 460 14329
rect 515 14320 715 14345
rect 796 14335 800 14395
rect 744 14329 800 14335
rect 515 14300 585 14320
rect 490 14260 585 14300
rect 645 14300 715 14320
rect 645 14260 740 14300
rect 490 14210 740 14260
rect 490 14170 585 14210
rect 515 14150 585 14170
rect 645 14170 740 14210
rect 645 14150 715 14170
rect 430 14135 486 14141
rect 430 14075 434 14135
rect 515 14125 715 14150
rect 770 14141 800 14329
rect 744 14135 800 14141
rect 486 14075 744 14095
rect 796 14075 800 14135
rect 430 14065 800 14075
rect 830 14395 1200 14405
rect 830 14335 834 14395
rect 886 14375 1144 14395
rect 830 14329 886 14335
rect 830 14141 860 14329
rect 915 14320 1115 14345
rect 1196 14335 1200 14395
rect 1144 14329 1200 14335
rect 915 14300 985 14320
rect 890 14260 985 14300
rect 1045 14300 1115 14320
rect 1045 14260 1140 14300
rect 890 14210 1140 14260
rect 890 14170 985 14210
rect 915 14150 985 14170
rect 1045 14170 1140 14210
rect 1045 14150 1115 14170
rect 830 14135 886 14141
rect 830 14075 834 14135
rect 915 14125 1115 14150
rect 1170 14141 1200 14329
rect 1144 14135 1200 14141
rect 886 14075 1144 14095
rect 1196 14075 1200 14135
rect 830 14065 1200 14075
rect 1230 14395 1600 14405
rect 1230 14335 1234 14395
rect 1286 14375 1544 14395
rect 1230 14329 1286 14335
rect 1230 14141 1260 14329
rect 1315 14320 1515 14345
rect 1596 14335 1600 14395
rect 1544 14329 1600 14335
rect 1315 14300 1385 14320
rect 1290 14260 1385 14300
rect 1445 14300 1515 14320
rect 1445 14260 1540 14300
rect 1290 14210 1540 14260
rect 1290 14170 1385 14210
rect 1315 14150 1385 14170
rect 1445 14170 1540 14210
rect 1445 14150 1515 14170
rect 1230 14135 1286 14141
rect 1230 14075 1234 14135
rect 1315 14125 1515 14150
rect 1570 14141 1600 14329
rect 1544 14135 1600 14141
rect 1286 14075 1544 14095
rect 1596 14075 1600 14135
rect 1230 14065 1600 14075
rect 1630 14395 2000 14405
rect 1630 14335 1634 14395
rect 1686 14375 1944 14395
rect 1630 14329 1686 14335
rect 1630 14141 1660 14329
rect 1715 14320 1915 14345
rect 1996 14335 2000 14395
rect 1944 14329 2000 14335
rect 1715 14300 1785 14320
rect 1690 14260 1785 14300
rect 1845 14300 1915 14320
rect 1845 14260 1940 14300
rect 1690 14210 1940 14260
rect 1690 14170 1785 14210
rect 1715 14150 1785 14170
rect 1845 14170 1940 14210
rect 1845 14150 1915 14170
rect 1630 14135 1686 14141
rect 1630 14075 1634 14135
rect 1715 14125 1915 14150
rect 1970 14141 2000 14329
rect 1944 14135 2000 14141
rect 1686 14075 1944 14095
rect 1996 14075 2000 14135
rect 1630 14065 2000 14075
rect 2030 14395 2400 14405
rect 2030 14335 2034 14395
rect 2086 14375 2344 14395
rect 2030 14329 2086 14335
rect 2030 14141 2060 14329
rect 2115 14320 2315 14345
rect 2396 14335 2400 14395
rect 2344 14329 2400 14335
rect 2115 14300 2185 14320
rect 2090 14260 2185 14300
rect 2245 14300 2315 14320
rect 2245 14260 2340 14300
rect 2090 14210 2340 14260
rect 2090 14170 2185 14210
rect 2115 14150 2185 14170
rect 2245 14170 2340 14210
rect 2245 14150 2315 14170
rect 2030 14135 2086 14141
rect 2030 14075 2034 14135
rect 2115 14125 2315 14150
rect 2370 14141 2400 14329
rect 2344 14135 2400 14141
rect 2086 14075 2344 14095
rect 2396 14075 2400 14135
rect 2030 14065 2400 14075
rect 2430 14395 2800 14405
rect 2430 14335 2434 14395
rect 2486 14375 2744 14395
rect 2430 14329 2486 14335
rect 2430 14141 2460 14329
rect 2515 14320 2715 14345
rect 2796 14335 2800 14395
rect 2744 14329 2800 14335
rect 2515 14300 2585 14320
rect 2490 14260 2585 14300
rect 2645 14300 2715 14320
rect 2645 14260 2740 14300
rect 2490 14210 2740 14260
rect 2490 14170 2585 14210
rect 2515 14150 2585 14170
rect 2645 14170 2740 14210
rect 2645 14150 2715 14170
rect 2430 14135 2486 14141
rect 2430 14075 2434 14135
rect 2515 14125 2715 14150
rect 2770 14141 2800 14329
rect 2744 14135 2800 14141
rect 2486 14075 2744 14095
rect 2796 14075 2800 14135
rect 2430 14065 2800 14075
rect 2830 14395 3200 14405
rect 2830 14335 2834 14395
rect 2886 14375 3144 14395
rect 2830 14329 2886 14335
rect 2830 14141 2860 14329
rect 2915 14320 3115 14345
rect 3196 14335 3200 14395
rect 3144 14329 3200 14335
rect 2915 14300 2985 14320
rect 2890 14260 2985 14300
rect 3045 14300 3115 14320
rect 3045 14260 3140 14300
rect 2890 14210 3140 14260
rect 2890 14170 2985 14210
rect 2915 14150 2985 14170
rect 3045 14170 3140 14210
rect 3045 14150 3115 14170
rect 2830 14135 2886 14141
rect 2830 14075 2834 14135
rect 2915 14125 3115 14150
rect 3170 14141 3200 14329
rect 3144 14135 3200 14141
rect 2886 14075 3144 14095
rect 3196 14075 3200 14135
rect 2830 14065 3200 14075
rect 3230 14395 3600 14405
rect 3230 14335 3234 14395
rect 3286 14375 3544 14395
rect 3230 14329 3286 14335
rect 3230 14141 3260 14329
rect 3315 14320 3515 14345
rect 3596 14335 3600 14395
rect 3544 14329 3600 14335
rect 3315 14300 3385 14320
rect 3290 14260 3385 14300
rect 3445 14300 3515 14320
rect 3445 14260 3540 14300
rect 3290 14210 3540 14260
rect 3290 14170 3385 14210
rect 3315 14150 3385 14170
rect 3445 14170 3540 14210
rect 3445 14150 3515 14170
rect 3230 14135 3286 14141
rect 3230 14075 3234 14135
rect 3315 14125 3515 14150
rect 3570 14141 3600 14329
rect 3544 14135 3600 14141
rect 3286 14075 3544 14095
rect 3596 14075 3600 14135
rect 3230 14065 3600 14075
rect 3630 14395 4000 14405
rect 3630 14335 3634 14395
rect 3686 14375 3944 14395
rect 3630 14329 3686 14335
rect 3630 14141 3660 14329
rect 3715 14320 3915 14345
rect 3996 14335 4000 14395
rect 3944 14329 4000 14335
rect 3715 14300 3785 14320
rect 3690 14260 3785 14300
rect 3845 14300 3915 14320
rect 3845 14260 3940 14300
rect 3690 14210 3940 14260
rect 3690 14170 3785 14210
rect 3715 14150 3785 14170
rect 3845 14170 3940 14210
rect 3845 14150 3915 14170
rect 3630 14135 3686 14141
rect 3630 14075 3634 14135
rect 3715 14125 3915 14150
rect 3970 14141 4000 14329
rect 3944 14135 4000 14141
rect 3686 14075 3944 14095
rect 3996 14075 4000 14135
rect 3630 14065 4000 14075
rect 4030 14395 4400 14405
rect 4030 14335 4034 14395
rect 4086 14375 4344 14395
rect 4030 14329 4086 14335
rect 4030 14141 4060 14329
rect 4115 14320 4315 14345
rect 4396 14335 4400 14395
rect 4344 14329 4400 14335
rect 4115 14300 4185 14320
rect 4090 14260 4185 14300
rect 4245 14300 4315 14320
rect 4245 14260 4340 14300
rect 4090 14210 4340 14260
rect 4090 14170 4185 14210
rect 4115 14150 4185 14170
rect 4245 14170 4340 14210
rect 4245 14150 4315 14170
rect 4030 14135 4086 14141
rect 4030 14075 4034 14135
rect 4115 14125 4315 14150
rect 4370 14141 4400 14329
rect 4344 14135 4400 14141
rect 4086 14075 4344 14095
rect 4396 14075 4400 14135
rect 4030 14065 4400 14075
rect 4430 14395 4800 14405
rect 4430 14335 4434 14395
rect 4486 14375 4744 14395
rect 4430 14329 4486 14335
rect 4430 14141 4460 14329
rect 4515 14320 4715 14345
rect 4796 14335 4800 14395
rect 4744 14329 4800 14335
rect 4515 14300 4585 14320
rect 4490 14260 4585 14300
rect 4645 14300 4715 14320
rect 4645 14260 4740 14300
rect 4490 14210 4740 14260
rect 4490 14170 4585 14210
rect 4515 14150 4585 14170
rect 4645 14170 4740 14210
rect 4645 14150 4715 14170
rect 4430 14135 4486 14141
rect 4430 14075 4434 14135
rect 4515 14125 4715 14150
rect 4770 14141 4800 14329
rect 4744 14135 4800 14141
rect 4486 14075 4744 14095
rect 4796 14075 4800 14135
rect 4430 14065 4800 14075
rect 4830 14395 5200 14405
rect 4830 14335 4834 14395
rect 4886 14375 5144 14395
rect 4830 14329 4886 14335
rect 4830 14141 4860 14329
rect 4915 14320 5115 14345
rect 5196 14335 5200 14395
rect 5144 14329 5200 14335
rect 4915 14300 4985 14320
rect 4890 14260 4985 14300
rect 5045 14300 5115 14320
rect 5045 14260 5140 14300
rect 4890 14210 5140 14260
rect 4890 14170 4985 14210
rect 4915 14150 4985 14170
rect 5045 14170 5140 14210
rect 5045 14150 5115 14170
rect 4830 14135 4886 14141
rect 4830 14075 4834 14135
rect 4915 14125 5115 14150
rect 5170 14141 5200 14329
rect 5144 14135 5200 14141
rect 4886 14075 5144 14095
rect 5196 14075 5200 14135
rect 4830 14065 5200 14075
rect 5230 14395 5600 14405
rect 5230 14335 5234 14395
rect 5286 14375 5544 14395
rect 5230 14329 5286 14335
rect 5230 14141 5260 14329
rect 5315 14320 5515 14345
rect 5596 14335 5600 14395
rect 5544 14329 5600 14335
rect 5315 14300 5385 14320
rect 5290 14260 5385 14300
rect 5445 14300 5515 14320
rect 5445 14260 5540 14300
rect 5290 14210 5540 14260
rect 5290 14170 5385 14210
rect 5315 14150 5385 14170
rect 5445 14170 5540 14210
rect 5445 14150 5515 14170
rect 5230 14135 5286 14141
rect 5230 14075 5234 14135
rect 5315 14125 5515 14150
rect 5570 14141 5600 14329
rect 5544 14135 5600 14141
rect 5286 14075 5544 14095
rect 5596 14075 5600 14135
rect 5230 14065 5600 14075
rect 5630 14395 6000 14405
rect 5630 14335 5634 14395
rect 5686 14375 5944 14395
rect 5630 14329 5686 14335
rect 5630 14141 5660 14329
rect 5715 14320 5915 14345
rect 5996 14335 6000 14395
rect 5944 14329 6000 14335
rect 5715 14300 5785 14320
rect 5690 14260 5785 14300
rect 5845 14300 5915 14320
rect 5845 14260 5940 14300
rect 5690 14210 5940 14260
rect 5690 14170 5785 14210
rect 5715 14150 5785 14170
rect 5845 14170 5940 14210
rect 5845 14150 5915 14170
rect 5630 14135 5686 14141
rect 5630 14075 5634 14135
rect 5715 14125 5915 14150
rect 5970 14141 6000 14329
rect 5944 14135 6000 14141
rect 5686 14075 5944 14095
rect 5996 14075 6000 14135
rect 5630 14065 6000 14075
rect 6030 14395 6400 14405
rect 6030 14335 6034 14395
rect 6086 14375 6344 14395
rect 6030 14329 6086 14335
rect 6030 14141 6060 14329
rect 6115 14320 6315 14345
rect 6396 14335 6400 14395
rect 6344 14329 6400 14335
rect 6115 14300 6185 14320
rect 6090 14260 6185 14300
rect 6245 14300 6315 14320
rect 6245 14260 6340 14300
rect 6090 14210 6340 14260
rect 6090 14170 6185 14210
rect 6115 14150 6185 14170
rect 6245 14170 6340 14210
rect 6245 14150 6315 14170
rect 6030 14135 6086 14141
rect 6030 14075 6034 14135
rect 6115 14125 6315 14150
rect 6370 14141 6400 14329
rect 6344 14135 6400 14141
rect 6086 14075 6344 14095
rect 6396 14075 6400 14135
rect 6030 14065 6400 14075
rect 6430 14395 6800 14405
rect 6430 14335 6434 14395
rect 6486 14375 6744 14395
rect 6430 14329 6486 14335
rect 6430 14141 6460 14329
rect 6515 14320 6715 14345
rect 6796 14335 6800 14395
rect 6744 14329 6800 14335
rect 6515 14300 6585 14320
rect 6490 14260 6585 14300
rect 6645 14300 6715 14320
rect 6645 14260 6740 14300
rect 6490 14210 6740 14260
rect 6490 14170 6585 14210
rect 6515 14150 6585 14170
rect 6645 14170 6740 14210
rect 6645 14150 6715 14170
rect 6430 14135 6486 14141
rect 6430 14075 6434 14135
rect 6515 14125 6715 14150
rect 6770 14141 6800 14329
rect 6744 14135 6800 14141
rect 6486 14075 6744 14095
rect 6796 14075 6800 14135
rect 6430 14065 6800 14075
rect 6830 14395 7200 14405
rect 6830 14335 6834 14395
rect 6886 14375 7144 14395
rect 6830 14329 6886 14335
rect 6830 14141 6860 14329
rect 6915 14320 7115 14345
rect 7196 14335 7200 14395
rect 7144 14329 7200 14335
rect 6915 14300 6985 14320
rect 6890 14260 6985 14300
rect 7045 14300 7115 14320
rect 7045 14260 7140 14300
rect 6890 14210 7140 14260
rect 6890 14170 6985 14210
rect 6915 14150 6985 14170
rect 7045 14170 7140 14210
rect 7045 14150 7115 14170
rect 6830 14135 6886 14141
rect 6830 14075 6834 14135
rect 6915 14125 7115 14150
rect 7170 14141 7200 14329
rect 7144 14135 7200 14141
rect 6886 14075 7144 14095
rect 7196 14075 7200 14135
rect 6830 14065 7200 14075
rect 7230 14395 7600 14405
rect 7230 14335 7234 14395
rect 7286 14375 7544 14395
rect 7230 14329 7286 14335
rect 7230 14141 7260 14329
rect 7315 14320 7515 14345
rect 7596 14335 7600 14395
rect 7544 14329 7600 14335
rect 7315 14300 7385 14320
rect 7290 14260 7385 14300
rect 7445 14300 7515 14320
rect 7445 14260 7540 14300
rect 7290 14210 7540 14260
rect 7290 14170 7385 14210
rect 7315 14150 7385 14170
rect 7445 14170 7540 14210
rect 7445 14150 7515 14170
rect 7230 14135 7286 14141
rect 7230 14075 7234 14135
rect 7315 14125 7515 14150
rect 7570 14141 7600 14329
rect 7544 14135 7600 14141
rect 7286 14075 7544 14095
rect 7596 14075 7600 14135
rect 7230 14065 7600 14075
rect 7630 14395 8000 14405
rect 7630 14335 7634 14395
rect 7686 14375 7944 14395
rect 7630 14329 7686 14335
rect 7630 14141 7660 14329
rect 7715 14320 7915 14345
rect 7996 14335 8000 14395
rect 7944 14329 8000 14335
rect 7715 14300 7785 14320
rect 7690 14260 7785 14300
rect 7845 14300 7915 14320
rect 7845 14260 7940 14300
rect 7690 14210 7940 14260
rect 7690 14170 7785 14210
rect 7715 14150 7785 14170
rect 7845 14170 7940 14210
rect 7845 14150 7915 14170
rect 7630 14135 7686 14141
rect 7630 14075 7634 14135
rect 7715 14125 7915 14150
rect 7970 14141 8000 14329
rect 7944 14135 8000 14141
rect 7686 14075 7944 14095
rect 7996 14075 8000 14135
rect 7630 14065 8000 14075
rect 8030 14395 8400 14405
rect 8030 14335 8034 14395
rect 8086 14375 8344 14395
rect 8030 14329 8086 14335
rect 8030 14141 8060 14329
rect 8115 14320 8315 14345
rect 8396 14335 8400 14395
rect 8344 14329 8400 14335
rect 8115 14300 8185 14320
rect 8090 14260 8185 14300
rect 8245 14300 8315 14320
rect 8245 14260 8340 14300
rect 8090 14210 8340 14260
rect 8090 14170 8185 14210
rect 8115 14150 8185 14170
rect 8245 14170 8340 14210
rect 8245 14150 8315 14170
rect 8030 14135 8086 14141
rect 8030 14075 8034 14135
rect 8115 14125 8315 14150
rect 8370 14141 8400 14329
rect 8344 14135 8400 14141
rect 8086 14075 8344 14095
rect 8396 14075 8400 14135
rect 8030 14065 8400 14075
rect 8430 14395 8800 14405
rect 8430 14335 8434 14395
rect 8486 14375 8744 14395
rect 8430 14329 8486 14335
rect 8430 14141 8460 14329
rect 8515 14320 8715 14345
rect 8796 14335 8800 14395
rect 8744 14329 8800 14335
rect 8515 14300 8585 14320
rect 8490 14260 8585 14300
rect 8645 14300 8715 14320
rect 8645 14260 8740 14300
rect 8490 14210 8740 14260
rect 8490 14170 8585 14210
rect 8515 14150 8585 14170
rect 8645 14170 8740 14210
rect 8645 14150 8715 14170
rect 8430 14135 8486 14141
rect 8430 14075 8434 14135
rect 8515 14125 8715 14150
rect 8770 14141 8800 14329
rect 8744 14135 8800 14141
rect 8486 14075 8744 14095
rect 8796 14075 8800 14135
rect 8430 14065 8800 14075
rect 8830 14395 9200 14405
rect 8830 14335 8834 14395
rect 8886 14375 9144 14395
rect 8830 14329 8886 14335
rect 8830 14141 8860 14329
rect 8915 14320 9115 14345
rect 9196 14335 9200 14395
rect 9144 14329 9200 14335
rect 8915 14300 8985 14320
rect 8890 14260 8985 14300
rect 9045 14300 9115 14320
rect 9045 14260 9140 14300
rect 8890 14210 9140 14260
rect 8890 14170 8985 14210
rect 8915 14150 8985 14170
rect 9045 14170 9140 14210
rect 9045 14150 9115 14170
rect 8830 14135 8886 14141
rect 8830 14075 8834 14135
rect 8915 14125 9115 14150
rect 9170 14141 9200 14329
rect 9144 14135 9200 14141
rect 8886 14075 9144 14095
rect 9196 14075 9200 14135
rect 8830 14065 9200 14075
rect 9230 14395 9600 14405
rect 9230 14335 9234 14395
rect 9286 14375 9544 14395
rect 9230 14329 9286 14335
rect 9230 14141 9260 14329
rect 9315 14320 9515 14345
rect 9596 14335 9600 14395
rect 9544 14329 9600 14335
rect 9315 14300 9385 14320
rect 9290 14260 9385 14300
rect 9445 14300 9515 14320
rect 9445 14260 9540 14300
rect 9290 14210 9540 14260
rect 9290 14170 9385 14210
rect 9315 14150 9385 14170
rect 9445 14170 9540 14210
rect 9445 14150 9515 14170
rect 9230 14135 9286 14141
rect 9230 14075 9234 14135
rect 9315 14125 9515 14150
rect 9570 14141 9600 14329
rect 9544 14135 9600 14141
rect 9286 14075 9544 14095
rect 9596 14075 9600 14135
rect 9230 14065 9600 14075
rect 9630 14395 10000 14405
rect 9630 14335 9634 14395
rect 9686 14375 9944 14395
rect 9630 14329 9686 14335
rect 9630 14141 9660 14329
rect 9715 14320 9915 14345
rect 9996 14335 10000 14395
rect 9944 14329 10000 14335
rect 9715 14300 9785 14320
rect 9690 14260 9785 14300
rect 9845 14300 9915 14320
rect 9845 14260 9940 14300
rect 9690 14210 9940 14260
rect 9690 14170 9785 14210
rect 9715 14150 9785 14170
rect 9845 14170 9940 14210
rect 9845 14150 9915 14170
rect 9630 14135 9686 14141
rect 9630 14075 9634 14135
rect 9715 14125 9915 14150
rect 9970 14141 10000 14329
rect 9944 14135 10000 14141
rect 9686 14075 9944 14095
rect 9996 14075 10000 14135
rect 9630 14065 10000 14075
rect 10030 14395 10400 14405
rect 10030 14335 10034 14395
rect 10086 14375 10344 14395
rect 10030 14329 10086 14335
rect 10030 14141 10060 14329
rect 10115 14320 10315 14345
rect 10396 14335 10400 14395
rect 10344 14329 10400 14335
rect 10115 14300 10185 14320
rect 10090 14260 10185 14300
rect 10245 14300 10315 14320
rect 10245 14260 10340 14300
rect 10090 14210 10340 14260
rect 10090 14170 10185 14210
rect 10115 14150 10185 14170
rect 10245 14170 10340 14210
rect 10245 14150 10315 14170
rect 10030 14135 10086 14141
rect 10030 14075 10034 14135
rect 10115 14125 10315 14150
rect 10370 14141 10400 14329
rect 10344 14135 10400 14141
rect 10086 14075 10344 14095
rect 10396 14075 10400 14135
rect 10030 14065 10400 14075
rect 10430 14395 10800 14405
rect 10430 14335 10434 14395
rect 10486 14375 10744 14395
rect 10430 14329 10486 14335
rect 10430 14141 10460 14329
rect 10515 14320 10715 14345
rect 10796 14335 10800 14395
rect 10744 14329 10800 14335
rect 10515 14300 10585 14320
rect 10490 14260 10585 14300
rect 10645 14300 10715 14320
rect 10645 14260 10740 14300
rect 10490 14210 10740 14260
rect 10490 14170 10585 14210
rect 10515 14150 10585 14170
rect 10645 14170 10740 14210
rect 10645 14150 10715 14170
rect 10430 14135 10486 14141
rect 10430 14075 10434 14135
rect 10515 14125 10715 14150
rect 10770 14141 10800 14329
rect 10744 14135 10800 14141
rect 10486 14075 10744 14095
rect 10796 14075 10800 14135
rect 10430 14065 10800 14075
rect 10830 14395 11200 14405
rect 10830 14335 10834 14395
rect 10886 14375 11144 14395
rect 10830 14329 10886 14335
rect 10830 14141 10860 14329
rect 10915 14320 11115 14345
rect 11196 14335 11200 14395
rect 11144 14329 11200 14335
rect 10915 14300 10985 14320
rect 10890 14260 10985 14300
rect 11045 14300 11115 14320
rect 11045 14260 11140 14300
rect 10890 14210 11140 14260
rect 10890 14170 10985 14210
rect 10915 14150 10985 14170
rect 11045 14170 11140 14210
rect 11045 14150 11115 14170
rect 10830 14135 10886 14141
rect 10830 14075 10834 14135
rect 10915 14125 11115 14150
rect 11170 14141 11200 14329
rect 11144 14135 11200 14141
rect 10886 14075 11144 14095
rect 11196 14075 11200 14135
rect 10830 14065 11200 14075
rect 11230 14395 11600 14405
rect 11230 14335 11234 14395
rect 11286 14375 11544 14395
rect 11230 14329 11286 14335
rect 11230 14141 11260 14329
rect 11315 14320 11515 14345
rect 11596 14335 11600 14395
rect 11544 14329 11600 14335
rect 11315 14300 11385 14320
rect 11290 14260 11385 14300
rect 11445 14300 11515 14320
rect 11445 14260 11540 14300
rect 11290 14210 11540 14260
rect 11290 14170 11385 14210
rect 11315 14150 11385 14170
rect 11445 14170 11540 14210
rect 11445 14150 11515 14170
rect 11230 14135 11286 14141
rect 11230 14075 11234 14135
rect 11315 14125 11515 14150
rect 11570 14141 11600 14329
rect 11544 14135 11600 14141
rect 11286 14075 11544 14095
rect 11596 14075 11600 14135
rect 11230 14065 11600 14075
rect 11630 14395 12000 14405
rect 11630 14335 11634 14395
rect 11686 14375 11944 14395
rect 11630 14329 11686 14335
rect 11630 14141 11660 14329
rect 11715 14320 11915 14345
rect 11996 14335 12000 14395
rect 11944 14329 12000 14335
rect 11715 14300 11785 14320
rect 11690 14260 11785 14300
rect 11845 14300 11915 14320
rect 11845 14260 11940 14300
rect 11690 14210 11940 14260
rect 11690 14170 11785 14210
rect 11715 14150 11785 14170
rect 11845 14170 11940 14210
rect 11845 14150 11915 14170
rect 11630 14135 11686 14141
rect 11630 14075 11634 14135
rect 11715 14125 11915 14150
rect 11970 14141 12000 14329
rect 11944 14135 12000 14141
rect 11686 14075 11944 14095
rect 11996 14075 12000 14135
rect 11630 14065 12000 14075
rect 12030 14395 12400 14405
rect 12030 14335 12034 14395
rect 12086 14375 12344 14395
rect 12030 14329 12086 14335
rect 12030 14141 12060 14329
rect 12115 14320 12315 14345
rect 12396 14335 12400 14395
rect 12344 14329 12400 14335
rect 12115 14300 12185 14320
rect 12090 14260 12185 14300
rect 12245 14300 12315 14320
rect 12245 14260 12340 14300
rect 12090 14210 12340 14260
rect 12090 14170 12185 14210
rect 12115 14150 12185 14170
rect 12245 14170 12340 14210
rect 12245 14150 12315 14170
rect 12030 14135 12086 14141
rect 12030 14075 12034 14135
rect 12115 14125 12315 14150
rect 12370 14141 12400 14329
rect 12344 14135 12400 14141
rect 12086 14075 12344 14095
rect 12396 14075 12400 14135
rect 12030 14065 12400 14075
rect 12430 14395 12800 14405
rect 12430 14335 12434 14395
rect 12486 14375 12744 14395
rect 12430 14329 12486 14335
rect 12430 14141 12460 14329
rect 12515 14320 12715 14345
rect 12796 14335 12800 14395
rect 12744 14329 12800 14335
rect 12515 14300 12585 14320
rect 12490 14260 12585 14300
rect 12645 14300 12715 14320
rect 12645 14260 12740 14300
rect 12490 14210 12740 14260
rect 12490 14170 12585 14210
rect 12515 14150 12585 14170
rect 12645 14170 12740 14210
rect 12645 14150 12715 14170
rect 12430 14135 12486 14141
rect 12430 14075 12434 14135
rect 12515 14125 12715 14150
rect 12770 14141 12800 14329
rect 12744 14135 12800 14141
rect 12486 14075 12744 14095
rect 12796 14075 12800 14135
rect 12430 14065 12800 14075
rect 12830 14395 13200 14405
rect 12830 14335 12834 14395
rect 12886 14375 13144 14395
rect 12830 14329 12886 14335
rect 12830 14141 12860 14329
rect 12915 14320 13115 14345
rect 13196 14335 13200 14395
rect 13144 14329 13200 14335
rect 12915 14300 12985 14320
rect 12890 14260 12985 14300
rect 13045 14300 13115 14320
rect 13045 14260 13140 14300
rect 12890 14210 13140 14260
rect 12890 14170 12985 14210
rect 12915 14150 12985 14170
rect 13045 14170 13140 14210
rect 13045 14150 13115 14170
rect 12830 14135 12886 14141
rect 12830 14075 12834 14135
rect 12915 14125 13115 14150
rect 13170 14141 13200 14329
rect 13144 14135 13200 14141
rect 12886 14075 13144 14095
rect 13196 14075 13200 14135
rect 12830 14065 13200 14075
rect -370 14025 0 14035
rect -370 13965 -366 14025
rect -314 14005 -56 14025
rect -370 13959 -314 13965
rect -370 13771 -340 13959
rect -285 13950 -85 13975
rect -4 13965 0 14025
rect -56 13959 0 13965
rect -285 13930 -215 13950
rect -310 13890 -215 13930
rect -155 13930 -85 13950
rect -155 13890 -60 13930
rect -310 13840 -60 13890
rect -310 13800 -215 13840
rect -285 13780 -215 13800
rect -155 13800 -60 13840
rect -155 13780 -85 13800
rect -370 13765 -314 13771
rect -370 13705 -366 13765
rect -285 13755 -85 13780
rect -30 13771 0 13959
rect -56 13765 0 13771
rect -314 13705 -56 13725
rect -4 13705 0 13765
rect -370 13695 0 13705
rect 30 14025 400 14035
rect 30 13965 34 14025
rect 86 14005 344 14025
rect 30 13959 86 13965
rect 30 13771 60 13959
rect 115 13950 315 13975
rect 396 13965 400 14025
rect 344 13959 400 13965
rect 115 13930 185 13950
rect 90 13890 185 13930
rect 245 13930 315 13950
rect 245 13890 340 13930
rect 90 13840 340 13890
rect 90 13800 185 13840
rect 115 13780 185 13800
rect 245 13800 340 13840
rect 245 13780 315 13800
rect 30 13765 86 13771
rect 30 13705 34 13765
rect 115 13755 315 13780
rect 370 13771 400 13959
rect 344 13765 400 13771
rect 86 13705 344 13725
rect 396 13705 400 13765
rect 30 13695 400 13705
rect 430 14025 800 14035
rect 430 13965 434 14025
rect 486 14005 744 14025
rect 430 13959 486 13965
rect 430 13771 460 13959
rect 515 13950 715 13975
rect 796 13965 800 14025
rect 744 13959 800 13965
rect 515 13930 585 13950
rect 490 13890 585 13930
rect 645 13930 715 13950
rect 645 13890 740 13930
rect 490 13840 740 13890
rect 490 13800 585 13840
rect 515 13780 585 13800
rect 645 13800 740 13840
rect 645 13780 715 13800
rect 430 13765 486 13771
rect 430 13705 434 13765
rect 515 13755 715 13780
rect 770 13771 800 13959
rect 744 13765 800 13771
rect 486 13705 744 13725
rect 796 13705 800 13765
rect 430 13695 800 13705
rect 830 14025 1200 14035
rect 830 13965 834 14025
rect 886 14005 1144 14025
rect 830 13959 886 13965
rect 830 13771 860 13959
rect 915 13950 1115 13975
rect 1196 13965 1200 14025
rect 1144 13959 1200 13965
rect 915 13930 985 13950
rect 890 13890 985 13930
rect 1045 13930 1115 13950
rect 1045 13890 1140 13930
rect 890 13840 1140 13890
rect 890 13800 985 13840
rect 915 13780 985 13800
rect 1045 13800 1140 13840
rect 1045 13780 1115 13800
rect 830 13765 886 13771
rect 830 13705 834 13765
rect 915 13755 1115 13780
rect 1170 13771 1200 13959
rect 1144 13765 1200 13771
rect 886 13705 1144 13725
rect 1196 13705 1200 13765
rect 830 13695 1200 13705
rect 1230 14025 1600 14035
rect 1230 13965 1234 14025
rect 1286 14005 1544 14025
rect 1230 13959 1286 13965
rect 1230 13771 1260 13959
rect 1315 13950 1515 13975
rect 1596 13965 1600 14025
rect 1544 13959 1600 13965
rect 1315 13930 1385 13950
rect 1290 13890 1385 13930
rect 1445 13930 1515 13950
rect 1445 13890 1540 13930
rect 1290 13840 1540 13890
rect 1290 13800 1385 13840
rect 1315 13780 1385 13800
rect 1445 13800 1540 13840
rect 1445 13780 1515 13800
rect 1230 13765 1286 13771
rect 1230 13705 1234 13765
rect 1315 13755 1515 13780
rect 1570 13771 1600 13959
rect 1544 13765 1600 13771
rect 1286 13705 1544 13725
rect 1596 13705 1600 13765
rect 1230 13695 1600 13705
rect 1630 14025 2000 14035
rect 1630 13965 1634 14025
rect 1686 14005 1944 14025
rect 1630 13959 1686 13965
rect 1630 13771 1660 13959
rect 1715 13950 1915 13975
rect 1996 13965 2000 14025
rect 1944 13959 2000 13965
rect 1715 13930 1785 13950
rect 1690 13890 1785 13930
rect 1845 13930 1915 13950
rect 1845 13890 1940 13930
rect 1690 13840 1940 13890
rect 1690 13800 1785 13840
rect 1715 13780 1785 13800
rect 1845 13800 1940 13840
rect 1845 13780 1915 13800
rect 1630 13765 1686 13771
rect 1630 13705 1634 13765
rect 1715 13755 1915 13780
rect 1970 13771 2000 13959
rect 1944 13765 2000 13771
rect 1686 13705 1944 13725
rect 1996 13705 2000 13765
rect 1630 13695 2000 13705
rect 2030 14025 2400 14035
rect 2030 13965 2034 14025
rect 2086 14005 2344 14025
rect 2030 13959 2086 13965
rect 2030 13771 2060 13959
rect 2115 13950 2315 13975
rect 2396 13965 2400 14025
rect 2344 13959 2400 13965
rect 2115 13930 2185 13950
rect 2090 13890 2185 13930
rect 2245 13930 2315 13950
rect 2245 13890 2340 13930
rect 2090 13840 2340 13890
rect 2090 13800 2185 13840
rect 2115 13780 2185 13800
rect 2245 13800 2340 13840
rect 2245 13780 2315 13800
rect 2030 13765 2086 13771
rect 2030 13705 2034 13765
rect 2115 13755 2315 13780
rect 2370 13771 2400 13959
rect 2344 13765 2400 13771
rect 2086 13705 2344 13725
rect 2396 13705 2400 13765
rect 2030 13695 2400 13705
rect 2430 14025 2800 14035
rect 2430 13965 2434 14025
rect 2486 14005 2744 14025
rect 2430 13959 2486 13965
rect 2430 13771 2460 13959
rect 2515 13950 2715 13975
rect 2796 13965 2800 14025
rect 2744 13959 2800 13965
rect 2515 13930 2585 13950
rect 2490 13890 2585 13930
rect 2645 13930 2715 13950
rect 2645 13890 2740 13930
rect 2490 13840 2740 13890
rect 2490 13800 2585 13840
rect 2515 13780 2585 13800
rect 2645 13800 2740 13840
rect 2645 13780 2715 13800
rect 2430 13765 2486 13771
rect 2430 13705 2434 13765
rect 2515 13755 2715 13780
rect 2770 13771 2800 13959
rect 2744 13765 2800 13771
rect 2486 13705 2744 13725
rect 2796 13705 2800 13765
rect 2430 13695 2800 13705
rect 2830 14025 3200 14035
rect 2830 13965 2834 14025
rect 2886 14005 3144 14025
rect 2830 13959 2886 13965
rect 2830 13771 2860 13959
rect 2915 13950 3115 13975
rect 3196 13965 3200 14025
rect 3144 13959 3200 13965
rect 2915 13930 2985 13950
rect 2890 13890 2985 13930
rect 3045 13930 3115 13950
rect 3045 13890 3140 13930
rect 2890 13840 3140 13890
rect 2890 13800 2985 13840
rect 2915 13780 2985 13800
rect 3045 13800 3140 13840
rect 3045 13780 3115 13800
rect 2830 13765 2886 13771
rect 2830 13705 2834 13765
rect 2915 13755 3115 13780
rect 3170 13771 3200 13959
rect 3144 13765 3200 13771
rect 2886 13705 3144 13725
rect 3196 13705 3200 13765
rect 2830 13695 3200 13705
rect 3230 14025 3600 14035
rect 3230 13965 3234 14025
rect 3286 14005 3544 14025
rect 3230 13959 3286 13965
rect 3230 13771 3260 13959
rect 3315 13950 3515 13975
rect 3596 13965 3600 14025
rect 3544 13959 3600 13965
rect 3315 13930 3385 13950
rect 3290 13890 3385 13930
rect 3445 13930 3515 13950
rect 3445 13890 3540 13930
rect 3290 13840 3540 13890
rect 3290 13800 3385 13840
rect 3315 13780 3385 13800
rect 3445 13800 3540 13840
rect 3445 13780 3515 13800
rect 3230 13765 3286 13771
rect 3230 13705 3234 13765
rect 3315 13755 3515 13780
rect 3570 13771 3600 13959
rect 3544 13765 3600 13771
rect 3286 13705 3544 13725
rect 3596 13705 3600 13765
rect 3230 13695 3600 13705
rect 3630 14025 4000 14035
rect 3630 13965 3634 14025
rect 3686 14005 3944 14025
rect 3630 13959 3686 13965
rect 3630 13771 3660 13959
rect 3715 13950 3915 13975
rect 3996 13965 4000 14025
rect 3944 13959 4000 13965
rect 3715 13930 3785 13950
rect 3690 13890 3785 13930
rect 3845 13930 3915 13950
rect 3845 13890 3940 13930
rect 3690 13840 3940 13890
rect 3690 13800 3785 13840
rect 3715 13780 3785 13800
rect 3845 13800 3940 13840
rect 3845 13780 3915 13800
rect 3630 13765 3686 13771
rect 3630 13705 3634 13765
rect 3715 13755 3915 13780
rect 3970 13771 4000 13959
rect 3944 13765 4000 13771
rect 3686 13705 3944 13725
rect 3996 13705 4000 13765
rect 3630 13695 4000 13705
rect 4030 14025 4400 14035
rect 4030 13965 4034 14025
rect 4086 14005 4344 14025
rect 4030 13959 4086 13965
rect 4030 13771 4060 13959
rect 4115 13950 4315 13975
rect 4396 13965 4400 14025
rect 4344 13959 4400 13965
rect 4115 13930 4185 13950
rect 4090 13890 4185 13930
rect 4245 13930 4315 13950
rect 4245 13890 4340 13930
rect 4090 13840 4340 13890
rect 4090 13800 4185 13840
rect 4115 13780 4185 13800
rect 4245 13800 4340 13840
rect 4245 13780 4315 13800
rect 4030 13765 4086 13771
rect 4030 13705 4034 13765
rect 4115 13755 4315 13780
rect 4370 13771 4400 13959
rect 4344 13765 4400 13771
rect 4086 13705 4344 13725
rect 4396 13705 4400 13765
rect 4030 13695 4400 13705
rect 4430 14025 4800 14035
rect 4430 13965 4434 14025
rect 4486 14005 4744 14025
rect 4430 13959 4486 13965
rect 4430 13771 4460 13959
rect 4515 13950 4715 13975
rect 4796 13965 4800 14025
rect 4744 13959 4800 13965
rect 4515 13930 4585 13950
rect 4490 13890 4585 13930
rect 4645 13930 4715 13950
rect 4645 13890 4740 13930
rect 4490 13840 4740 13890
rect 4490 13800 4585 13840
rect 4515 13780 4585 13800
rect 4645 13800 4740 13840
rect 4645 13780 4715 13800
rect 4430 13765 4486 13771
rect 4430 13705 4434 13765
rect 4515 13755 4715 13780
rect 4770 13771 4800 13959
rect 4744 13765 4800 13771
rect 4486 13705 4744 13725
rect 4796 13705 4800 13765
rect 4430 13695 4800 13705
rect 4830 14025 5200 14035
rect 4830 13965 4834 14025
rect 4886 14005 5144 14025
rect 4830 13959 4886 13965
rect 4830 13771 4860 13959
rect 4915 13950 5115 13975
rect 5196 13965 5200 14025
rect 5144 13959 5200 13965
rect 4915 13930 4985 13950
rect 4890 13890 4985 13930
rect 5045 13930 5115 13950
rect 5045 13890 5140 13930
rect 4890 13840 5140 13890
rect 4890 13800 4985 13840
rect 4915 13780 4985 13800
rect 5045 13800 5140 13840
rect 5045 13780 5115 13800
rect 4830 13765 4886 13771
rect 4830 13705 4834 13765
rect 4915 13755 5115 13780
rect 5170 13771 5200 13959
rect 5144 13765 5200 13771
rect 4886 13705 5144 13725
rect 5196 13705 5200 13765
rect 4830 13695 5200 13705
rect 5230 14025 5600 14035
rect 5230 13965 5234 14025
rect 5286 14005 5544 14025
rect 5230 13959 5286 13965
rect 5230 13771 5260 13959
rect 5315 13950 5515 13975
rect 5596 13965 5600 14025
rect 5544 13959 5600 13965
rect 5315 13930 5385 13950
rect 5290 13890 5385 13930
rect 5445 13930 5515 13950
rect 5445 13890 5540 13930
rect 5290 13840 5540 13890
rect 5290 13800 5385 13840
rect 5315 13780 5385 13800
rect 5445 13800 5540 13840
rect 5445 13780 5515 13800
rect 5230 13765 5286 13771
rect 5230 13705 5234 13765
rect 5315 13755 5515 13780
rect 5570 13771 5600 13959
rect 5544 13765 5600 13771
rect 5286 13705 5544 13725
rect 5596 13705 5600 13765
rect 5230 13695 5600 13705
rect 5630 14025 6000 14035
rect 5630 13965 5634 14025
rect 5686 14005 5944 14025
rect 5630 13959 5686 13965
rect 5630 13771 5660 13959
rect 5715 13950 5915 13975
rect 5996 13965 6000 14025
rect 5944 13959 6000 13965
rect 5715 13930 5785 13950
rect 5690 13890 5785 13930
rect 5845 13930 5915 13950
rect 5845 13890 5940 13930
rect 5690 13840 5940 13890
rect 5690 13800 5785 13840
rect 5715 13780 5785 13800
rect 5845 13800 5940 13840
rect 5845 13780 5915 13800
rect 5630 13765 5686 13771
rect 5630 13705 5634 13765
rect 5715 13755 5915 13780
rect 5970 13771 6000 13959
rect 5944 13765 6000 13771
rect 5686 13705 5944 13725
rect 5996 13705 6000 13765
rect 5630 13695 6000 13705
rect 6030 14025 6400 14035
rect 6030 13965 6034 14025
rect 6086 14005 6344 14025
rect 6030 13959 6086 13965
rect 6030 13771 6060 13959
rect 6115 13950 6315 13975
rect 6396 13965 6400 14025
rect 6344 13959 6400 13965
rect 6115 13930 6185 13950
rect 6090 13890 6185 13930
rect 6245 13930 6315 13950
rect 6245 13890 6340 13930
rect 6090 13840 6340 13890
rect 6090 13800 6185 13840
rect 6115 13780 6185 13800
rect 6245 13800 6340 13840
rect 6245 13780 6315 13800
rect 6030 13765 6086 13771
rect 6030 13705 6034 13765
rect 6115 13755 6315 13780
rect 6370 13771 6400 13959
rect 6344 13765 6400 13771
rect 6086 13705 6344 13725
rect 6396 13705 6400 13765
rect 6030 13695 6400 13705
rect 6430 14025 6800 14035
rect 6430 13965 6434 14025
rect 6486 14005 6744 14025
rect 6430 13959 6486 13965
rect 6430 13771 6460 13959
rect 6515 13950 6715 13975
rect 6796 13965 6800 14025
rect 6744 13959 6800 13965
rect 6515 13930 6585 13950
rect 6490 13890 6585 13930
rect 6645 13930 6715 13950
rect 6645 13890 6740 13930
rect 6490 13840 6740 13890
rect 6490 13800 6585 13840
rect 6515 13780 6585 13800
rect 6645 13800 6740 13840
rect 6645 13780 6715 13800
rect 6430 13765 6486 13771
rect 6430 13705 6434 13765
rect 6515 13755 6715 13780
rect 6770 13771 6800 13959
rect 6744 13765 6800 13771
rect 6486 13705 6744 13725
rect 6796 13705 6800 13765
rect 6430 13695 6800 13705
rect 6830 14025 7200 14035
rect 6830 13965 6834 14025
rect 6886 14005 7144 14025
rect 6830 13959 6886 13965
rect 6830 13771 6860 13959
rect 6915 13950 7115 13975
rect 7196 13965 7200 14025
rect 7144 13959 7200 13965
rect 6915 13930 6985 13950
rect 6890 13890 6985 13930
rect 7045 13930 7115 13950
rect 7045 13890 7140 13930
rect 6890 13840 7140 13890
rect 6890 13800 6985 13840
rect 6915 13780 6985 13800
rect 7045 13800 7140 13840
rect 7045 13780 7115 13800
rect 6830 13765 6886 13771
rect 6830 13705 6834 13765
rect 6915 13755 7115 13780
rect 7170 13771 7200 13959
rect 7144 13765 7200 13771
rect 6886 13705 7144 13725
rect 7196 13705 7200 13765
rect 6830 13695 7200 13705
rect 7230 14025 7600 14035
rect 7230 13965 7234 14025
rect 7286 14005 7544 14025
rect 7230 13959 7286 13965
rect 7230 13771 7260 13959
rect 7315 13950 7515 13975
rect 7596 13965 7600 14025
rect 7544 13959 7600 13965
rect 7315 13930 7385 13950
rect 7290 13890 7385 13930
rect 7445 13930 7515 13950
rect 7445 13890 7540 13930
rect 7290 13840 7540 13890
rect 7290 13800 7385 13840
rect 7315 13780 7385 13800
rect 7445 13800 7540 13840
rect 7445 13780 7515 13800
rect 7230 13765 7286 13771
rect 7230 13705 7234 13765
rect 7315 13755 7515 13780
rect 7570 13771 7600 13959
rect 7544 13765 7600 13771
rect 7286 13705 7544 13725
rect 7596 13705 7600 13765
rect 7230 13695 7600 13705
rect 7630 14025 8000 14035
rect 7630 13965 7634 14025
rect 7686 14005 7944 14025
rect 7630 13959 7686 13965
rect 7630 13771 7660 13959
rect 7715 13950 7915 13975
rect 7996 13965 8000 14025
rect 7944 13959 8000 13965
rect 7715 13930 7785 13950
rect 7690 13890 7785 13930
rect 7845 13930 7915 13950
rect 7845 13890 7940 13930
rect 7690 13840 7940 13890
rect 7690 13800 7785 13840
rect 7715 13780 7785 13800
rect 7845 13800 7940 13840
rect 7845 13780 7915 13800
rect 7630 13765 7686 13771
rect 7630 13705 7634 13765
rect 7715 13755 7915 13780
rect 7970 13771 8000 13959
rect 7944 13765 8000 13771
rect 7686 13705 7944 13725
rect 7996 13705 8000 13765
rect 7630 13695 8000 13705
rect 8030 14025 8400 14035
rect 8030 13965 8034 14025
rect 8086 14005 8344 14025
rect 8030 13959 8086 13965
rect 8030 13771 8060 13959
rect 8115 13950 8315 13975
rect 8396 13965 8400 14025
rect 8344 13959 8400 13965
rect 8115 13930 8185 13950
rect 8090 13890 8185 13930
rect 8245 13930 8315 13950
rect 8245 13890 8340 13930
rect 8090 13840 8340 13890
rect 8090 13800 8185 13840
rect 8115 13780 8185 13800
rect 8245 13800 8340 13840
rect 8245 13780 8315 13800
rect 8030 13765 8086 13771
rect 8030 13705 8034 13765
rect 8115 13755 8315 13780
rect 8370 13771 8400 13959
rect 8344 13765 8400 13771
rect 8086 13705 8344 13725
rect 8396 13705 8400 13765
rect 8030 13695 8400 13705
rect 8430 14025 8800 14035
rect 8430 13965 8434 14025
rect 8486 14005 8744 14025
rect 8430 13959 8486 13965
rect 8430 13771 8460 13959
rect 8515 13950 8715 13975
rect 8796 13965 8800 14025
rect 8744 13959 8800 13965
rect 8515 13930 8585 13950
rect 8490 13890 8585 13930
rect 8645 13930 8715 13950
rect 8645 13890 8740 13930
rect 8490 13840 8740 13890
rect 8490 13800 8585 13840
rect 8515 13780 8585 13800
rect 8645 13800 8740 13840
rect 8645 13780 8715 13800
rect 8430 13765 8486 13771
rect 8430 13705 8434 13765
rect 8515 13755 8715 13780
rect 8770 13771 8800 13959
rect 8744 13765 8800 13771
rect 8486 13705 8744 13725
rect 8796 13705 8800 13765
rect 8430 13695 8800 13705
rect 8830 14025 9200 14035
rect 8830 13965 8834 14025
rect 8886 14005 9144 14025
rect 8830 13959 8886 13965
rect 8830 13771 8860 13959
rect 8915 13950 9115 13975
rect 9196 13965 9200 14025
rect 9144 13959 9200 13965
rect 8915 13930 8985 13950
rect 8890 13890 8985 13930
rect 9045 13930 9115 13950
rect 9045 13890 9140 13930
rect 8890 13840 9140 13890
rect 8890 13800 8985 13840
rect 8915 13780 8985 13800
rect 9045 13800 9140 13840
rect 9045 13780 9115 13800
rect 8830 13765 8886 13771
rect 8830 13705 8834 13765
rect 8915 13755 9115 13780
rect 9170 13771 9200 13959
rect 9144 13765 9200 13771
rect 8886 13705 9144 13725
rect 9196 13705 9200 13765
rect 8830 13695 9200 13705
rect 9230 14025 9600 14035
rect 9230 13965 9234 14025
rect 9286 14005 9544 14025
rect 9230 13959 9286 13965
rect 9230 13771 9260 13959
rect 9315 13950 9515 13975
rect 9596 13965 9600 14025
rect 9544 13959 9600 13965
rect 9315 13930 9385 13950
rect 9290 13890 9385 13930
rect 9445 13930 9515 13950
rect 9445 13890 9540 13930
rect 9290 13840 9540 13890
rect 9290 13800 9385 13840
rect 9315 13780 9385 13800
rect 9445 13800 9540 13840
rect 9445 13780 9515 13800
rect 9230 13765 9286 13771
rect 9230 13705 9234 13765
rect 9315 13755 9515 13780
rect 9570 13771 9600 13959
rect 9544 13765 9600 13771
rect 9286 13705 9544 13725
rect 9596 13705 9600 13765
rect 9230 13695 9600 13705
rect 9630 14025 10000 14035
rect 9630 13965 9634 14025
rect 9686 14005 9944 14025
rect 9630 13959 9686 13965
rect 9630 13771 9660 13959
rect 9715 13950 9915 13975
rect 9996 13965 10000 14025
rect 9944 13959 10000 13965
rect 9715 13930 9785 13950
rect 9690 13890 9785 13930
rect 9845 13930 9915 13950
rect 9845 13890 9940 13930
rect 9690 13840 9940 13890
rect 9690 13800 9785 13840
rect 9715 13780 9785 13800
rect 9845 13800 9940 13840
rect 9845 13780 9915 13800
rect 9630 13765 9686 13771
rect 9630 13705 9634 13765
rect 9715 13755 9915 13780
rect 9970 13771 10000 13959
rect 9944 13765 10000 13771
rect 9686 13705 9944 13725
rect 9996 13705 10000 13765
rect 9630 13695 10000 13705
rect 10030 14025 10400 14035
rect 10030 13965 10034 14025
rect 10086 14005 10344 14025
rect 10030 13959 10086 13965
rect 10030 13771 10060 13959
rect 10115 13950 10315 13975
rect 10396 13965 10400 14025
rect 10344 13959 10400 13965
rect 10115 13930 10185 13950
rect 10090 13890 10185 13930
rect 10245 13930 10315 13950
rect 10245 13890 10340 13930
rect 10090 13840 10340 13890
rect 10090 13800 10185 13840
rect 10115 13780 10185 13800
rect 10245 13800 10340 13840
rect 10245 13780 10315 13800
rect 10030 13765 10086 13771
rect 10030 13705 10034 13765
rect 10115 13755 10315 13780
rect 10370 13771 10400 13959
rect 10344 13765 10400 13771
rect 10086 13705 10344 13725
rect 10396 13705 10400 13765
rect 10030 13695 10400 13705
rect 10430 14025 10800 14035
rect 10430 13965 10434 14025
rect 10486 14005 10744 14025
rect 10430 13959 10486 13965
rect 10430 13771 10460 13959
rect 10515 13950 10715 13975
rect 10796 13965 10800 14025
rect 10744 13959 10800 13965
rect 10515 13930 10585 13950
rect 10490 13890 10585 13930
rect 10645 13930 10715 13950
rect 10645 13890 10740 13930
rect 10490 13840 10740 13890
rect 10490 13800 10585 13840
rect 10515 13780 10585 13800
rect 10645 13800 10740 13840
rect 10645 13780 10715 13800
rect 10430 13765 10486 13771
rect 10430 13705 10434 13765
rect 10515 13755 10715 13780
rect 10770 13771 10800 13959
rect 10744 13765 10800 13771
rect 10486 13705 10744 13725
rect 10796 13705 10800 13765
rect 10430 13695 10800 13705
rect 10830 14025 11200 14035
rect 10830 13965 10834 14025
rect 10886 14005 11144 14025
rect 10830 13959 10886 13965
rect 10830 13771 10860 13959
rect 10915 13950 11115 13975
rect 11196 13965 11200 14025
rect 11144 13959 11200 13965
rect 10915 13930 10985 13950
rect 10890 13890 10985 13930
rect 11045 13930 11115 13950
rect 11045 13890 11140 13930
rect 10890 13840 11140 13890
rect 10890 13800 10985 13840
rect 10915 13780 10985 13800
rect 11045 13800 11140 13840
rect 11045 13780 11115 13800
rect 10830 13765 10886 13771
rect 10830 13705 10834 13765
rect 10915 13755 11115 13780
rect 11170 13771 11200 13959
rect 11144 13765 11200 13771
rect 10886 13705 11144 13725
rect 11196 13705 11200 13765
rect 10830 13695 11200 13705
rect 11230 14025 11600 14035
rect 11230 13965 11234 14025
rect 11286 14005 11544 14025
rect 11230 13959 11286 13965
rect 11230 13771 11260 13959
rect 11315 13950 11515 13975
rect 11596 13965 11600 14025
rect 11544 13959 11600 13965
rect 11315 13930 11385 13950
rect 11290 13890 11385 13930
rect 11445 13930 11515 13950
rect 11445 13890 11540 13930
rect 11290 13840 11540 13890
rect 11290 13800 11385 13840
rect 11315 13780 11385 13800
rect 11445 13800 11540 13840
rect 11445 13780 11515 13800
rect 11230 13765 11286 13771
rect 11230 13705 11234 13765
rect 11315 13755 11515 13780
rect 11570 13771 11600 13959
rect 11544 13765 11600 13771
rect 11286 13705 11544 13725
rect 11596 13705 11600 13765
rect 11230 13695 11600 13705
rect 11630 14025 12000 14035
rect 11630 13965 11634 14025
rect 11686 14005 11944 14025
rect 11630 13959 11686 13965
rect 11630 13771 11660 13959
rect 11715 13950 11915 13975
rect 11996 13965 12000 14025
rect 11944 13959 12000 13965
rect 11715 13930 11785 13950
rect 11690 13890 11785 13930
rect 11845 13930 11915 13950
rect 11845 13890 11940 13930
rect 11690 13840 11940 13890
rect 11690 13800 11785 13840
rect 11715 13780 11785 13800
rect 11845 13800 11940 13840
rect 11845 13780 11915 13800
rect 11630 13765 11686 13771
rect 11630 13705 11634 13765
rect 11715 13755 11915 13780
rect 11970 13771 12000 13959
rect 11944 13765 12000 13771
rect 11686 13705 11944 13725
rect 11996 13705 12000 13765
rect 11630 13695 12000 13705
rect 12030 14025 12400 14035
rect 12030 13965 12034 14025
rect 12086 14005 12344 14025
rect 12030 13959 12086 13965
rect 12030 13771 12060 13959
rect 12115 13950 12315 13975
rect 12396 13965 12400 14025
rect 12344 13959 12400 13965
rect 12115 13930 12185 13950
rect 12090 13890 12185 13930
rect 12245 13930 12315 13950
rect 12245 13890 12340 13930
rect 12090 13840 12340 13890
rect 12090 13800 12185 13840
rect 12115 13780 12185 13800
rect 12245 13800 12340 13840
rect 12245 13780 12315 13800
rect 12030 13765 12086 13771
rect 12030 13705 12034 13765
rect 12115 13755 12315 13780
rect 12370 13771 12400 13959
rect 12344 13765 12400 13771
rect 12086 13705 12344 13725
rect 12396 13705 12400 13765
rect 12030 13695 12400 13705
rect 12430 14025 12800 14035
rect 12430 13965 12434 14025
rect 12486 14005 12744 14025
rect 12430 13959 12486 13965
rect 12430 13771 12460 13959
rect 12515 13950 12715 13975
rect 12796 13965 12800 14025
rect 12744 13959 12800 13965
rect 12515 13930 12585 13950
rect 12490 13890 12585 13930
rect 12645 13930 12715 13950
rect 12645 13890 12740 13930
rect 12490 13840 12740 13890
rect 12490 13800 12585 13840
rect 12515 13780 12585 13800
rect 12645 13800 12740 13840
rect 12645 13780 12715 13800
rect 12430 13765 12486 13771
rect 12430 13705 12434 13765
rect 12515 13755 12715 13780
rect 12770 13771 12800 13959
rect 12744 13765 12800 13771
rect 12486 13705 12744 13725
rect 12796 13705 12800 13765
rect 12430 13695 12800 13705
rect 12830 14025 13200 14035
rect 12830 13965 12834 14025
rect 12886 14005 13144 14025
rect 12830 13959 12886 13965
rect 12830 13771 12860 13959
rect 12915 13950 13115 13975
rect 13196 13965 13200 14025
rect 13144 13959 13200 13965
rect 12915 13930 12985 13950
rect 12890 13890 12985 13930
rect 13045 13930 13115 13950
rect 13045 13890 13140 13930
rect 12890 13840 13140 13890
rect 12890 13800 12985 13840
rect 12915 13780 12985 13800
rect 13045 13800 13140 13840
rect 13045 13780 13115 13800
rect 12830 13765 12886 13771
rect 12830 13705 12834 13765
rect 12915 13755 13115 13780
rect 13170 13771 13200 13959
rect 13144 13765 13200 13771
rect 12886 13705 13144 13725
rect 13196 13705 13200 13765
rect 12830 13695 13200 13705
rect -370 13655 0 13665
rect -370 13595 -366 13655
rect -314 13635 -56 13655
rect -370 13589 -314 13595
rect -370 13401 -340 13589
rect -285 13580 -85 13605
rect -4 13595 0 13655
rect -56 13589 0 13595
rect -285 13560 -215 13580
rect -310 13520 -215 13560
rect -155 13560 -85 13580
rect -155 13520 -60 13560
rect -310 13470 -60 13520
rect -310 13430 -215 13470
rect -285 13410 -215 13430
rect -155 13430 -60 13470
rect -155 13410 -85 13430
rect -370 13395 -314 13401
rect -370 13335 -366 13395
rect -285 13385 -85 13410
rect -30 13401 0 13589
rect -56 13395 0 13401
rect -314 13335 -56 13355
rect -4 13335 0 13395
rect -370 13325 0 13335
rect 30 13655 400 13665
rect 30 13595 34 13655
rect 86 13635 344 13655
rect 30 13589 86 13595
rect 30 13401 60 13589
rect 115 13580 315 13605
rect 396 13595 400 13655
rect 344 13589 400 13595
rect 115 13560 185 13580
rect 90 13520 185 13560
rect 245 13560 315 13580
rect 245 13520 340 13560
rect 90 13470 340 13520
rect 90 13430 185 13470
rect 115 13410 185 13430
rect 245 13430 340 13470
rect 245 13410 315 13430
rect 30 13395 86 13401
rect 30 13335 34 13395
rect 115 13385 315 13410
rect 370 13401 400 13589
rect 344 13395 400 13401
rect 86 13335 344 13355
rect 396 13335 400 13395
rect 30 13325 400 13335
rect 430 13655 800 13665
rect 430 13595 434 13655
rect 486 13635 744 13655
rect 430 13589 486 13595
rect 430 13401 460 13589
rect 515 13580 715 13605
rect 796 13595 800 13655
rect 744 13589 800 13595
rect 515 13560 585 13580
rect 490 13520 585 13560
rect 645 13560 715 13580
rect 645 13520 740 13560
rect 490 13470 740 13520
rect 490 13430 585 13470
rect 515 13410 585 13430
rect 645 13430 740 13470
rect 645 13410 715 13430
rect 430 13395 486 13401
rect 430 13335 434 13395
rect 515 13385 715 13410
rect 770 13401 800 13589
rect 744 13395 800 13401
rect 486 13335 744 13355
rect 796 13335 800 13395
rect 430 13325 800 13335
rect 830 13655 1200 13665
rect 830 13595 834 13655
rect 886 13635 1144 13655
rect 830 13589 886 13595
rect 830 13401 860 13589
rect 915 13580 1115 13605
rect 1196 13595 1200 13655
rect 1144 13589 1200 13595
rect 915 13560 985 13580
rect 890 13520 985 13560
rect 1045 13560 1115 13580
rect 1045 13520 1140 13560
rect 890 13470 1140 13520
rect 890 13430 985 13470
rect 915 13410 985 13430
rect 1045 13430 1140 13470
rect 1045 13410 1115 13430
rect 830 13395 886 13401
rect 830 13335 834 13395
rect 915 13385 1115 13410
rect 1170 13401 1200 13589
rect 1144 13395 1200 13401
rect 886 13335 1144 13355
rect 1196 13335 1200 13395
rect 830 13325 1200 13335
rect 1230 13655 1600 13665
rect 1230 13595 1234 13655
rect 1286 13635 1544 13655
rect 1230 13589 1286 13595
rect 1230 13401 1260 13589
rect 1315 13580 1515 13605
rect 1596 13595 1600 13655
rect 1544 13589 1600 13595
rect 1315 13560 1385 13580
rect 1290 13520 1385 13560
rect 1445 13560 1515 13580
rect 1445 13520 1540 13560
rect 1290 13470 1540 13520
rect 1290 13430 1385 13470
rect 1315 13410 1385 13430
rect 1445 13430 1540 13470
rect 1445 13410 1515 13430
rect 1230 13395 1286 13401
rect 1230 13335 1234 13395
rect 1315 13385 1515 13410
rect 1570 13401 1600 13589
rect 1544 13395 1600 13401
rect 1286 13335 1544 13355
rect 1596 13335 1600 13395
rect 1230 13325 1600 13335
rect 1630 13655 2000 13665
rect 1630 13595 1634 13655
rect 1686 13635 1944 13655
rect 1630 13589 1686 13595
rect 1630 13401 1660 13589
rect 1715 13580 1915 13605
rect 1996 13595 2000 13655
rect 1944 13589 2000 13595
rect 1715 13560 1785 13580
rect 1690 13520 1785 13560
rect 1845 13560 1915 13580
rect 1845 13520 1940 13560
rect 1690 13470 1940 13520
rect 1690 13430 1785 13470
rect 1715 13410 1785 13430
rect 1845 13430 1940 13470
rect 1845 13410 1915 13430
rect 1630 13395 1686 13401
rect 1630 13335 1634 13395
rect 1715 13385 1915 13410
rect 1970 13401 2000 13589
rect 1944 13395 2000 13401
rect 1686 13335 1944 13355
rect 1996 13335 2000 13395
rect 1630 13325 2000 13335
rect 2030 13655 2400 13665
rect 2030 13595 2034 13655
rect 2086 13635 2344 13655
rect 2030 13589 2086 13595
rect 2030 13401 2060 13589
rect 2115 13580 2315 13605
rect 2396 13595 2400 13655
rect 2344 13589 2400 13595
rect 2115 13560 2185 13580
rect 2090 13520 2185 13560
rect 2245 13560 2315 13580
rect 2245 13520 2340 13560
rect 2090 13470 2340 13520
rect 2090 13430 2185 13470
rect 2115 13410 2185 13430
rect 2245 13430 2340 13470
rect 2245 13410 2315 13430
rect 2030 13395 2086 13401
rect 2030 13335 2034 13395
rect 2115 13385 2315 13410
rect 2370 13401 2400 13589
rect 2344 13395 2400 13401
rect 2086 13335 2344 13355
rect 2396 13335 2400 13395
rect 2030 13325 2400 13335
rect 2430 13655 2800 13665
rect 2430 13595 2434 13655
rect 2486 13635 2744 13655
rect 2430 13589 2486 13595
rect 2430 13401 2460 13589
rect 2515 13580 2715 13605
rect 2796 13595 2800 13655
rect 2744 13589 2800 13595
rect 2515 13560 2585 13580
rect 2490 13520 2585 13560
rect 2645 13560 2715 13580
rect 2645 13520 2740 13560
rect 2490 13470 2740 13520
rect 2490 13430 2585 13470
rect 2515 13410 2585 13430
rect 2645 13430 2740 13470
rect 2645 13410 2715 13430
rect 2430 13395 2486 13401
rect 2430 13335 2434 13395
rect 2515 13385 2715 13410
rect 2770 13401 2800 13589
rect 2744 13395 2800 13401
rect 2486 13335 2744 13355
rect 2796 13335 2800 13395
rect 2430 13325 2800 13335
rect 2830 13655 3200 13665
rect 2830 13595 2834 13655
rect 2886 13635 3144 13655
rect 2830 13589 2886 13595
rect 2830 13401 2860 13589
rect 2915 13580 3115 13605
rect 3196 13595 3200 13655
rect 3144 13589 3200 13595
rect 2915 13560 2985 13580
rect 2890 13520 2985 13560
rect 3045 13560 3115 13580
rect 3045 13520 3140 13560
rect 2890 13470 3140 13520
rect 2890 13430 2985 13470
rect 2915 13410 2985 13430
rect 3045 13430 3140 13470
rect 3045 13410 3115 13430
rect 2830 13395 2886 13401
rect 2830 13335 2834 13395
rect 2915 13385 3115 13410
rect 3170 13401 3200 13589
rect 3144 13395 3200 13401
rect 2886 13335 3144 13355
rect 3196 13335 3200 13395
rect 2830 13325 3200 13335
rect 3230 13655 3600 13665
rect 3230 13595 3234 13655
rect 3286 13635 3544 13655
rect 3230 13589 3286 13595
rect 3230 13401 3260 13589
rect 3315 13580 3515 13605
rect 3596 13595 3600 13655
rect 3544 13589 3600 13595
rect 3315 13560 3385 13580
rect 3290 13520 3385 13560
rect 3445 13560 3515 13580
rect 3445 13520 3540 13560
rect 3290 13470 3540 13520
rect 3290 13430 3385 13470
rect 3315 13410 3385 13430
rect 3445 13430 3540 13470
rect 3445 13410 3515 13430
rect 3230 13395 3286 13401
rect 3230 13335 3234 13395
rect 3315 13385 3515 13410
rect 3570 13401 3600 13589
rect 3544 13395 3600 13401
rect 3286 13335 3544 13355
rect 3596 13335 3600 13395
rect 3230 13325 3600 13335
rect 3630 13655 4000 13665
rect 3630 13595 3634 13655
rect 3686 13635 3944 13655
rect 3630 13589 3686 13595
rect 3630 13401 3660 13589
rect 3715 13580 3915 13605
rect 3996 13595 4000 13655
rect 3944 13589 4000 13595
rect 3715 13560 3785 13580
rect 3690 13520 3785 13560
rect 3845 13560 3915 13580
rect 3845 13520 3940 13560
rect 3690 13470 3940 13520
rect 3690 13430 3785 13470
rect 3715 13410 3785 13430
rect 3845 13430 3940 13470
rect 3845 13410 3915 13430
rect 3630 13395 3686 13401
rect 3630 13335 3634 13395
rect 3715 13385 3915 13410
rect 3970 13401 4000 13589
rect 3944 13395 4000 13401
rect 3686 13335 3944 13355
rect 3996 13335 4000 13395
rect 3630 13325 4000 13335
rect 4030 13655 4400 13665
rect 4030 13595 4034 13655
rect 4086 13635 4344 13655
rect 4030 13589 4086 13595
rect 4030 13401 4060 13589
rect 4115 13580 4315 13605
rect 4396 13595 4400 13655
rect 4344 13589 4400 13595
rect 4115 13560 4185 13580
rect 4090 13520 4185 13560
rect 4245 13560 4315 13580
rect 4245 13520 4340 13560
rect 4090 13470 4340 13520
rect 4090 13430 4185 13470
rect 4115 13410 4185 13430
rect 4245 13430 4340 13470
rect 4245 13410 4315 13430
rect 4030 13395 4086 13401
rect 4030 13335 4034 13395
rect 4115 13385 4315 13410
rect 4370 13401 4400 13589
rect 4344 13395 4400 13401
rect 4086 13335 4344 13355
rect 4396 13335 4400 13395
rect 4030 13325 4400 13335
rect 4430 13655 4800 13665
rect 4430 13595 4434 13655
rect 4486 13635 4744 13655
rect 4430 13589 4486 13595
rect 4430 13401 4460 13589
rect 4515 13580 4715 13605
rect 4796 13595 4800 13655
rect 4744 13589 4800 13595
rect 4515 13560 4585 13580
rect 4490 13520 4585 13560
rect 4645 13560 4715 13580
rect 4645 13520 4740 13560
rect 4490 13470 4740 13520
rect 4490 13430 4585 13470
rect 4515 13410 4585 13430
rect 4645 13430 4740 13470
rect 4645 13410 4715 13430
rect 4430 13395 4486 13401
rect 4430 13335 4434 13395
rect 4515 13385 4715 13410
rect 4770 13401 4800 13589
rect 4744 13395 4800 13401
rect 4486 13335 4744 13355
rect 4796 13335 4800 13395
rect 4430 13325 4800 13335
rect 4830 13655 5200 13665
rect 4830 13595 4834 13655
rect 4886 13635 5144 13655
rect 4830 13589 4886 13595
rect 4830 13401 4860 13589
rect 4915 13580 5115 13605
rect 5196 13595 5200 13655
rect 5144 13589 5200 13595
rect 4915 13560 4985 13580
rect 4890 13520 4985 13560
rect 5045 13560 5115 13580
rect 5045 13520 5140 13560
rect 4890 13470 5140 13520
rect 4890 13430 4985 13470
rect 4915 13410 4985 13430
rect 5045 13430 5140 13470
rect 5045 13410 5115 13430
rect 4830 13395 4886 13401
rect 4830 13335 4834 13395
rect 4915 13385 5115 13410
rect 5170 13401 5200 13589
rect 5144 13395 5200 13401
rect 4886 13335 5144 13355
rect 5196 13335 5200 13395
rect 4830 13325 5200 13335
rect 5230 13655 5600 13665
rect 5230 13595 5234 13655
rect 5286 13635 5544 13655
rect 5230 13589 5286 13595
rect 5230 13401 5260 13589
rect 5315 13580 5515 13605
rect 5596 13595 5600 13655
rect 5544 13589 5600 13595
rect 5315 13560 5385 13580
rect 5290 13520 5385 13560
rect 5445 13560 5515 13580
rect 5445 13520 5540 13560
rect 5290 13470 5540 13520
rect 5290 13430 5385 13470
rect 5315 13410 5385 13430
rect 5445 13430 5540 13470
rect 5445 13410 5515 13430
rect 5230 13395 5286 13401
rect 5230 13335 5234 13395
rect 5315 13385 5515 13410
rect 5570 13401 5600 13589
rect 5544 13395 5600 13401
rect 5286 13335 5544 13355
rect 5596 13335 5600 13395
rect 5230 13325 5600 13335
rect 5630 13655 6000 13665
rect 5630 13595 5634 13655
rect 5686 13635 5944 13655
rect 5630 13589 5686 13595
rect 5630 13401 5660 13589
rect 5715 13580 5915 13605
rect 5996 13595 6000 13655
rect 5944 13589 6000 13595
rect 5715 13560 5785 13580
rect 5690 13520 5785 13560
rect 5845 13560 5915 13580
rect 5845 13520 5940 13560
rect 5690 13470 5940 13520
rect 5690 13430 5785 13470
rect 5715 13410 5785 13430
rect 5845 13430 5940 13470
rect 5845 13410 5915 13430
rect 5630 13395 5686 13401
rect 5630 13335 5634 13395
rect 5715 13385 5915 13410
rect 5970 13401 6000 13589
rect 5944 13395 6000 13401
rect 5686 13335 5944 13355
rect 5996 13335 6000 13395
rect 5630 13325 6000 13335
rect 6030 13655 6400 13665
rect 6030 13595 6034 13655
rect 6086 13635 6344 13655
rect 6030 13589 6086 13595
rect 6030 13401 6060 13589
rect 6115 13580 6315 13605
rect 6396 13595 6400 13655
rect 6344 13589 6400 13595
rect 6115 13560 6185 13580
rect 6090 13520 6185 13560
rect 6245 13560 6315 13580
rect 6245 13520 6340 13560
rect 6090 13470 6340 13520
rect 6090 13430 6185 13470
rect 6115 13410 6185 13430
rect 6245 13430 6340 13470
rect 6245 13410 6315 13430
rect 6030 13395 6086 13401
rect 6030 13335 6034 13395
rect 6115 13385 6315 13410
rect 6370 13401 6400 13589
rect 6344 13395 6400 13401
rect 6086 13335 6344 13355
rect 6396 13335 6400 13395
rect 6030 13325 6400 13335
rect 6430 13655 6800 13665
rect 6430 13595 6434 13655
rect 6486 13635 6744 13655
rect 6430 13589 6486 13595
rect 6430 13401 6460 13589
rect 6515 13580 6715 13605
rect 6796 13595 6800 13655
rect 6744 13589 6800 13595
rect 6515 13560 6585 13580
rect 6490 13520 6585 13560
rect 6645 13560 6715 13580
rect 6645 13520 6740 13560
rect 6490 13470 6740 13520
rect 6490 13430 6585 13470
rect 6515 13410 6585 13430
rect 6645 13430 6740 13470
rect 6645 13410 6715 13430
rect 6430 13395 6486 13401
rect 6430 13335 6434 13395
rect 6515 13385 6715 13410
rect 6770 13401 6800 13589
rect 6744 13395 6800 13401
rect 6486 13335 6744 13355
rect 6796 13335 6800 13395
rect 6430 13325 6800 13335
rect 6830 13655 7200 13665
rect 6830 13595 6834 13655
rect 6886 13635 7144 13655
rect 6830 13589 6886 13595
rect 6830 13401 6860 13589
rect 6915 13580 7115 13605
rect 7196 13595 7200 13655
rect 7144 13589 7200 13595
rect 6915 13560 6985 13580
rect 6890 13520 6985 13560
rect 7045 13560 7115 13580
rect 7045 13520 7140 13560
rect 6890 13470 7140 13520
rect 6890 13430 6985 13470
rect 6915 13410 6985 13430
rect 7045 13430 7140 13470
rect 7045 13410 7115 13430
rect 6830 13395 6886 13401
rect 6830 13335 6834 13395
rect 6915 13385 7115 13410
rect 7170 13401 7200 13589
rect 7144 13395 7200 13401
rect 6886 13335 7144 13355
rect 7196 13335 7200 13395
rect 6830 13325 7200 13335
rect 7230 13655 7600 13665
rect 7230 13595 7234 13655
rect 7286 13635 7544 13655
rect 7230 13589 7286 13595
rect 7230 13401 7260 13589
rect 7315 13580 7515 13605
rect 7596 13595 7600 13655
rect 7544 13589 7600 13595
rect 7315 13560 7385 13580
rect 7290 13520 7385 13560
rect 7445 13560 7515 13580
rect 7445 13520 7540 13560
rect 7290 13470 7540 13520
rect 7290 13430 7385 13470
rect 7315 13410 7385 13430
rect 7445 13430 7540 13470
rect 7445 13410 7515 13430
rect 7230 13395 7286 13401
rect 7230 13335 7234 13395
rect 7315 13385 7515 13410
rect 7570 13401 7600 13589
rect 7544 13395 7600 13401
rect 7286 13335 7544 13355
rect 7596 13335 7600 13395
rect 7230 13325 7600 13335
rect 7630 13655 8000 13665
rect 7630 13595 7634 13655
rect 7686 13635 7944 13655
rect 7630 13589 7686 13595
rect 7630 13401 7660 13589
rect 7715 13580 7915 13605
rect 7996 13595 8000 13655
rect 7944 13589 8000 13595
rect 7715 13560 7785 13580
rect 7690 13520 7785 13560
rect 7845 13560 7915 13580
rect 7845 13520 7940 13560
rect 7690 13470 7940 13520
rect 7690 13430 7785 13470
rect 7715 13410 7785 13430
rect 7845 13430 7940 13470
rect 7845 13410 7915 13430
rect 7630 13395 7686 13401
rect 7630 13335 7634 13395
rect 7715 13385 7915 13410
rect 7970 13401 8000 13589
rect 7944 13395 8000 13401
rect 7686 13335 7944 13355
rect 7996 13335 8000 13395
rect 7630 13325 8000 13335
rect 8030 13655 8400 13665
rect 8030 13595 8034 13655
rect 8086 13635 8344 13655
rect 8030 13589 8086 13595
rect 8030 13401 8060 13589
rect 8115 13580 8315 13605
rect 8396 13595 8400 13655
rect 8344 13589 8400 13595
rect 8115 13560 8185 13580
rect 8090 13520 8185 13560
rect 8245 13560 8315 13580
rect 8245 13520 8340 13560
rect 8090 13470 8340 13520
rect 8090 13430 8185 13470
rect 8115 13410 8185 13430
rect 8245 13430 8340 13470
rect 8245 13410 8315 13430
rect 8030 13395 8086 13401
rect 8030 13335 8034 13395
rect 8115 13385 8315 13410
rect 8370 13401 8400 13589
rect 8344 13395 8400 13401
rect 8086 13335 8344 13355
rect 8396 13335 8400 13395
rect 8030 13325 8400 13335
rect 8430 13655 8800 13665
rect 8430 13595 8434 13655
rect 8486 13635 8744 13655
rect 8430 13589 8486 13595
rect 8430 13401 8460 13589
rect 8515 13580 8715 13605
rect 8796 13595 8800 13655
rect 8744 13589 8800 13595
rect 8515 13560 8585 13580
rect 8490 13520 8585 13560
rect 8645 13560 8715 13580
rect 8645 13520 8740 13560
rect 8490 13470 8740 13520
rect 8490 13430 8585 13470
rect 8515 13410 8585 13430
rect 8645 13430 8740 13470
rect 8645 13410 8715 13430
rect 8430 13395 8486 13401
rect 8430 13335 8434 13395
rect 8515 13385 8715 13410
rect 8770 13401 8800 13589
rect 8744 13395 8800 13401
rect 8486 13335 8744 13355
rect 8796 13335 8800 13395
rect 8430 13325 8800 13335
rect 8830 13655 9200 13665
rect 8830 13595 8834 13655
rect 8886 13635 9144 13655
rect 8830 13589 8886 13595
rect 8830 13401 8860 13589
rect 8915 13580 9115 13605
rect 9196 13595 9200 13655
rect 9144 13589 9200 13595
rect 8915 13560 8985 13580
rect 8890 13520 8985 13560
rect 9045 13560 9115 13580
rect 9045 13520 9140 13560
rect 8890 13470 9140 13520
rect 8890 13430 8985 13470
rect 8915 13410 8985 13430
rect 9045 13430 9140 13470
rect 9045 13410 9115 13430
rect 8830 13395 8886 13401
rect 8830 13335 8834 13395
rect 8915 13385 9115 13410
rect 9170 13401 9200 13589
rect 9144 13395 9200 13401
rect 8886 13335 9144 13355
rect 9196 13335 9200 13395
rect 8830 13325 9200 13335
rect 9230 13655 9600 13665
rect 9230 13595 9234 13655
rect 9286 13635 9544 13655
rect 9230 13589 9286 13595
rect 9230 13401 9260 13589
rect 9315 13580 9515 13605
rect 9596 13595 9600 13655
rect 9544 13589 9600 13595
rect 9315 13560 9385 13580
rect 9290 13520 9385 13560
rect 9445 13560 9515 13580
rect 9445 13520 9540 13560
rect 9290 13470 9540 13520
rect 9290 13430 9385 13470
rect 9315 13410 9385 13430
rect 9445 13430 9540 13470
rect 9445 13410 9515 13430
rect 9230 13395 9286 13401
rect 9230 13335 9234 13395
rect 9315 13385 9515 13410
rect 9570 13401 9600 13589
rect 9544 13395 9600 13401
rect 9286 13335 9544 13355
rect 9596 13335 9600 13395
rect 9230 13325 9600 13335
rect 9630 13655 10000 13665
rect 9630 13595 9634 13655
rect 9686 13635 9944 13655
rect 9630 13589 9686 13595
rect 9630 13401 9660 13589
rect 9715 13580 9915 13605
rect 9996 13595 10000 13655
rect 9944 13589 10000 13595
rect 9715 13560 9785 13580
rect 9690 13520 9785 13560
rect 9845 13560 9915 13580
rect 9845 13520 9940 13560
rect 9690 13470 9940 13520
rect 9690 13430 9785 13470
rect 9715 13410 9785 13430
rect 9845 13430 9940 13470
rect 9845 13410 9915 13430
rect 9630 13395 9686 13401
rect 9630 13335 9634 13395
rect 9715 13385 9915 13410
rect 9970 13401 10000 13589
rect 9944 13395 10000 13401
rect 9686 13335 9944 13355
rect 9996 13335 10000 13395
rect 9630 13325 10000 13335
rect 10030 13655 10400 13665
rect 10030 13595 10034 13655
rect 10086 13635 10344 13655
rect 10030 13589 10086 13595
rect 10030 13401 10060 13589
rect 10115 13580 10315 13605
rect 10396 13595 10400 13655
rect 10344 13589 10400 13595
rect 10115 13560 10185 13580
rect 10090 13520 10185 13560
rect 10245 13560 10315 13580
rect 10245 13520 10340 13560
rect 10090 13470 10340 13520
rect 10090 13430 10185 13470
rect 10115 13410 10185 13430
rect 10245 13430 10340 13470
rect 10245 13410 10315 13430
rect 10030 13395 10086 13401
rect 10030 13335 10034 13395
rect 10115 13385 10315 13410
rect 10370 13401 10400 13589
rect 10344 13395 10400 13401
rect 10086 13335 10344 13355
rect 10396 13335 10400 13395
rect 10030 13325 10400 13335
rect 10430 13655 10800 13665
rect 10430 13595 10434 13655
rect 10486 13635 10744 13655
rect 10430 13589 10486 13595
rect 10430 13401 10460 13589
rect 10515 13580 10715 13605
rect 10796 13595 10800 13655
rect 10744 13589 10800 13595
rect 10515 13560 10585 13580
rect 10490 13520 10585 13560
rect 10645 13560 10715 13580
rect 10645 13520 10740 13560
rect 10490 13470 10740 13520
rect 10490 13430 10585 13470
rect 10515 13410 10585 13430
rect 10645 13430 10740 13470
rect 10645 13410 10715 13430
rect 10430 13395 10486 13401
rect 10430 13335 10434 13395
rect 10515 13385 10715 13410
rect 10770 13401 10800 13589
rect 10744 13395 10800 13401
rect 10486 13335 10744 13355
rect 10796 13335 10800 13395
rect 10430 13325 10800 13335
rect 10830 13655 11200 13665
rect 10830 13595 10834 13655
rect 10886 13635 11144 13655
rect 10830 13589 10886 13595
rect 10830 13401 10860 13589
rect 10915 13580 11115 13605
rect 11196 13595 11200 13655
rect 11144 13589 11200 13595
rect 10915 13560 10985 13580
rect 10890 13520 10985 13560
rect 11045 13560 11115 13580
rect 11045 13520 11140 13560
rect 10890 13470 11140 13520
rect 10890 13430 10985 13470
rect 10915 13410 10985 13430
rect 11045 13430 11140 13470
rect 11045 13410 11115 13430
rect 10830 13395 10886 13401
rect 10830 13335 10834 13395
rect 10915 13385 11115 13410
rect 11170 13401 11200 13589
rect 11144 13395 11200 13401
rect 10886 13335 11144 13355
rect 11196 13335 11200 13395
rect 10830 13325 11200 13335
rect 11230 13655 11600 13665
rect 11230 13595 11234 13655
rect 11286 13635 11544 13655
rect 11230 13589 11286 13595
rect 11230 13401 11260 13589
rect 11315 13580 11515 13605
rect 11596 13595 11600 13655
rect 11544 13589 11600 13595
rect 11315 13560 11385 13580
rect 11290 13520 11385 13560
rect 11445 13560 11515 13580
rect 11445 13520 11540 13560
rect 11290 13470 11540 13520
rect 11290 13430 11385 13470
rect 11315 13410 11385 13430
rect 11445 13430 11540 13470
rect 11445 13410 11515 13430
rect 11230 13395 11286 13401
rect 11230 13335 11234 13395
rect 11315 13385 11515 13410
rect 11570 13401 11600 13589
rect 11544 13395 11600 13401
rect 11286 13335 11544 13355
rect 11596 13335 11600 13395
rect 11230 13325 11600 13335
rect 11630 13655 12000 13665
rect 11630 13595 11634 13655
rect 11686 13635 11944 13655
rect 11630 13589 11686 13595
rect 11630 13401 11660 13589
rect 11715 13580 11915 13605
rect 11996 13595 12000 13655
rect 11944 13589 12000 13595
rect 11715 13560 11785 13580
rect 11690 13520 11785 13560
rect 11845 13560 11915 13580
rect 11845 13520 11940 13560
rect 11690 13470 11940 13520
rect 11690 13430 11785 13470
rect 11715 13410 11785 13430
rect 11845 13430 11940 13470
rect 11845 13410 11915 13430
rect 11630 13395 11686 13401
rect 11630 13335 11634 13395
rect 11715 13385 11915 13410
rect 11970 13401 12000 13589
rect 11944 13395 12000 13401
rect 11686 13335 11944 13355
rect 11996 13335 12000 13395
rect 11630 13325 12000 13335
rect 12030 13655 12400 13665
rect 12030 13595 12034 13655
rect 12086 13635 12344 13655
rect 12030 13589 12086 13595
rect 12030 13401 12060 13589
rect 12115 13580 12315 13605
rect 12396 13595 12400 13655
rect 12344 13589 12400 13595
rect 12115 13560 12185 13580
rect 12090 13520 12185 13560
rect 12245 13560 12315 13580
rect 12245 13520 12340 13560
rect 12090 13470 12340 13520
rect 12090 13430 12185 13470
rect 12115 13410 12185 13430
rect 12245 13430 12340 13470
rect 12245 13410 12315 13430
rect 12030 13395 12086 13401
rect 12030 13335 12034 13395
rect 12115 13385 12315 13410
rect 12370 13401 12400 13589
rect 12344 13395 12400 13401
rect 12086 13335 12344 13355
rect 12396 13335 12400 13395
rect 12030 13325 12400 13335
rect 12430 13655 12800 13665
rect 12430 13595 12434 13655
rect 12486 13635 12744 13655
rect 12430 13589 12486 13595
rect 12430 13401 12460 13589
rect 12515 13580 12715 13605
rect 12796 13595 12800 13655
rect 12744 13589 12800 13595
rect 12515 13560 12585 13580
rect 12490 13520 12585 13560
rect 12645 13560 12715 13580
rect 12645 13520 12740 13560
rect 12490 13470 12740 13520
rect 12490 13430 12585 13470
rect 12515 13410 12585 13430
rect 12645 13430 12740 13470
rect 12645 13410 12715 13430
rect 12430 13395 12486 13401
rect 12430 13335 12434 13395
rect 12515 13385 12715 13410
rect 12770 13401 12800 13589
rect 12744 13395 12800 13401
rect 12486 13335 12744 13355
rect 12796 13335 12800 13395
rect 12430 13325 12800 13335
rect 12830 13655 13200 13665
rect 12830 13595 12834 13655
rect 12886 13635 13144 13655
rect 12830 13589 12886 13595
rect 12830 13401 12860 13589
rect 12915 13580 13115 13605
rect 13196 13595 13200 13655
rect 13144 13589 13200 13595
rect 12915 13560 12985 13580
rect 12890 13520 12985 13560
rect 13045 13560 13115 13580
rect 13045 13520 13140 13560
rect 12890 13470 13140 13520
rect 12890 13430 12985 13470
rect 12915 13410 12985 13430
rect 13045 13430 13140 13470
rect 13045 13410 13115 13430
rect 12830 13395 12886 13401
rect 12830 13335 12834 13395
rect 12915 13385 13115 13410
rect 13170 13401 13200 13589
rect 13144 13395 13200 13401
rect 12886 13335 13144 13355
rect 13196 13335 13200 13395
rect 12830 13325 13200 13335
rect -370 13285 0 13295
rect -370 13225 -366 13285
rect -314 13265 -56 13285
rect -370 13219 -314 13225
rect -370 13031 -340 13219
rect -285 13210 -85 13235
rect -4 13225 0 13285
rect -56 13219 0 13225
rect -285 13190 -215 13210
rect -310 13150 -215 13190
rect -155 13190 -85 13210
rect -155 13150 -60 13190
rect -310 13100 -60 13150
rect -310 13060 -215 13100
rect -285 13040 -215 13060
rect -155 13060 -60 13100
rect -155 13040 -85 13060
rect -370 13025 -314 13031
rect -370 12965 -366 13025
rect -285 13015 -85 13040
rect -30 13031 0 13219
rect -56 13025 0 13031
rect -314 12965 -56 12985
rect -4 12965 0 13025
rect -370 12955 0 12965
rect 30 13285 400 13295
rect 30 13225 34 13285
rect 86 13265 344 13285
rect 30 13219 86 13225
rect 30 13031 60 13219
rect 115 13210 315 13235
rect 396 13225 400 13285
rect 344 13219 400 13225
rect 115 13190 185 13210
rect 90 13150 185 13190
rect 245 13190 315 13210
rect 245 13150 340 13190
rect 90 13100 340 13150
rect 90 13060 185 13100
rect 115 13040 185 13060
rect 245 13060 340 13100
rect 245 13040 315 13060
rect 30 13025 86 13031
rect 30 12965 34 13025
rect 115 13015 315 13040
rect 370 13031 400 13219
rect 344 13025 400 13031
rect 86 12965 344 12985
rect 396 12965 400 13025
rect 30 12955 400 12965
rect 430 13285 800 13295
rect 430 13225 434 13285
rect 486 13265 744 13285
rect 430 13219 486 13225
rect 430 13031 460 13219
rect 515 13210 715 13235
rect 796 13225 800 13285
rect 744 13219 800 13225
rect 515 13190 585 13210
rect 490 13150 585 13190
rect 645 13190 715 13210
rect 645 13150 740 13190
rect 490 13100 740 13150
rect 490 13060 585 13100
rect 515 13040 585 13060
rect 645 13060 740 13100
rect 645 13040 715 13060
rect 430 13025 486 13031
rect 430 12965 434 13025
rect 515 13015 715 13040
rect 770 13031 800 13219
rect 744 13025 800 13031
rect 486 12965 744 12985
rect 796 12965 800 13025
rect 430 12955 800 12965
rect 830 13285 1200 13295
rect 830 13225 834 13285
rect 886 13265 1144 13285
rect 830 13219 886 13225
rect 830 13031 860 13219
rect 915 13210 1115 13235
rect 1196 13225 1200 13285
rect 1144 13219 1200 13225
rect 915 13190 985 13210
rect 890 13150 985 13190
rect 1045 13190 1115 13210
rect 1045 13150 1140 13190
rect 890 13100 1140 13150
rect 890 13060 985 13100
rect 915 13040 985 13060
rect 1045 13060 1140 13100
rect 1045 13040 1115 13060
rect 830 13025 886 13031
rect 830 12965 834 13025
rect 915 13015 1115 13040
rect 1170 13031 1200 13219
rect 1144 13025 1200 13031
rect 886 12965 1144 12985
rect 1196 12965 1200 13025
rect 830 12955 1200 12965
rect 1230 13285 1600 13295
rect 1230 13225 1234 13285
rect 1286 13265 1544 13285
rect 1230 13219 1286 13225
rect 1230 13031 1260 13219
rect 1315 13210 1515 13235
rect 1596 13225 1600 13285
rect 1544 13219 1600 13225
rect 1315 13190 1385 13210
rect 1290 13150 1385 13190
rect 1445 13190 1515 13210
rect 1445 13150 1540 13190
rect 1290 13100 1540 13150
rect 1290 13060 1385 13100
rect 1315 13040 1385 13060
rect 1445 13060 1540 13100
rect 1445 13040 1515 13060
rect 1230 13025 1286 13031
rect 1230 12965 1234 13025
rect 1315 13015 1515 13040
rect 1570 13031 1600 13219
rect 1544 13025 1600 13031
rect 1286 12965 1544 12985
rect 1596 12965 1600 13025
rect 1230 12955 1600 12965
rect 1630 13285 2000 13295
rect 1630 13225 1634 13285
rect 1686 13265 1944 13285
rect 1630 13219 1686 13225
rect 1630 13031 1660 13219
rect 1715 13210 1915 13235
rect 1996 13225 2000 13285
rect 1944 13219 2000 13225
rect 1715 13190 1785 13210
rect 1690 13150 1785 13190
rect 1845 13190 1915 13210
rect 1845 13150 1940 13190
rect 1690 13100 1940 13150
rect 1690 13060 1785 13100
rect 1715 13040 1785 13060
rect 1845 13060 1940 13100
rect 1845 13040 1915 13060
rect 1630 13025 1686 13031
rect 1630 12965 1634 13025
rect 1715 13015 1915 13040
rect 1970 13031 2000 13219
rect 1944 13025 2000 13031
rect 1686 12965 1944 12985
rect 1996 12965 2000 13025
rect 1630 12955 2000 12965
rect 2030 13285 2400 13295
rect 2030 13225 2034 13285
rect 2086 13265 2344 13285
rect 2030 13219 2086 13225
rect 2030 13031 2060 13219
rect 2115 13210 2315 13235
rect 2396 13225 2400 13285
rect 2344 13219 2400 13225
rect 2115 13190 2185 13210
rect 2090 13150 2185 13190
rect 2245 13190 2315 13210
rect 2245 13150 2340 13190
rect 2090 13100 2340 13150
rect 2090 13060 2185 13100
rect 2115 13040 2185 13060
rect 2245 13060 2340 13100
rect 2245 13040 2315 13060
rect 2030 13025 2086 13031
rect 2030 12965 2034 13025
rect 2115 13015 2315 13040
rect 2370 13031 2400 13219
rect 2344 13025 2400 13031
rect 2086 12965 2344 12985
rect 2396 12965 2400 13025
rect 2030 12955 2400 12965
rect 2430 13285 2800 13295
rect 2430 13225 2434 13285
rect 2486 13265 2744 13285
rect 2430 13219 2486 13225
rect 2430 13031 2460 13219
rect 2515 13210 2715 13235
rect 2796 13225 2800 13285
rect 2744 13219 2800 13225
rect 2515 13190 2585 13210
rect 2490 13150 2585 13190
rect 2645 13190 2715 13210
rect 2645 13150 2740 13190
rect 2490 13100 2740 13150
rect 2490 13060 2585 13100
rect 2515 13040 2585 13060
rect 2645 13060 2740 13100
rect 2645 13040 2715 13060
rect 2430 13025 2486 13031
rect 2430 12965 2434 13025
rect 2515 13015 2715 13040
rect 2770 13031 2800 13219
rect 2744 13025 2800 13031
rect 2486 12965 2744 12985
rect 2796 12965 2800 13025
rect 2430 12955 2800 12965
rect 2830 13285 3200 13295
rect 2830 13225 2834 13285
rect 2886 13265 3144 13285
rect 2830 13219 2886 13225
rect 2830 13031 2860 13219
rect 2915 13210 3115 13235
rect 3196 13225 3200 13285
rect 3144 13219 3200 13225
rect 2915 13190 2985 13210
rect 2890 13150 2985 13190
rect 3045 13190 3115 13210
rect 3045 13150 3140 13190
rect 2890 13100 3140 13150
rect 2890 13060 2985 13100
rect 2915 13040 2985 13060
rect 3045 13060 3140 13100
rect 3045 13040 3115 13060
rect 2830 13025 2886 13031
rect 2830 12965 2834 13025
rect 2915 13015 3115 13040
rect 3170 13031 3200 13219
rect 3144 13025 3200 13031
rect 2886 12965 3144 12985
rect 3196 12965 3200 13025
rect 2830 12955 3200 12965
rect 3230 13285 3600 13295
rect 3230 13225 3234 13285
rect 3286 13265 3544 13285
rect 3230 13219 3286 13225
rect 3230 13031 3260 13219
rect 3315 13210 3515 13235
rect 3596 13225 3600 13285
rect 3544 13219 3600 13225
rect 3315 13190 3385 13210
rect 3290 13150 3385 13190
rect 3445 13190 3515 13210
rect 3445 13150 3540 13190
rect 3290 13100 3540 13150
rect 3290 13060 3385 13100
rect 3315 13040 3385 13060
rect 3445 13060 3540 13100
rect 3445 13040 3515 13060
rect 3230 13025 3286 13031
rect 3230 12965 3234 13025
rect 3315 13015 3515 13040
rect 3570 13031 3600 13219
rect 3544 13025 3600 13031
rect 3286 12965 3544 12985
rect 3596 12965 3600 13025
rect 3230 12955 3600 12965
rect 3630 13285 4000 13295
rect 3630 13225 3634 13285
rect 3686 13265 3944 13285
rect 3630 13219 3686 13225
rect 3630 13031 3660 13219
rect 3715 13210 3915 13235
rect 3996 13225 4000 13285
rect 3944 13219 4000 13225
rect 3715 13190 3785 13210
rect 3690 13150 3785 13190
rect 3845 13190 3915 13210
rect 3845 13150 3940 13190
rect 3690 13100 3940 13150
rect 3690 13060 3785 13100
rect 3715 13040 3785 13060
rect 3845 13060 3940 13100
rect 3845 13040 3915 13060
rect 3630 13025 3686 13031
rect 3630 12965 3634 13025
rect 3715 13015 3915 13040
rect 3970 13031 4000 13219
rect 3944 13025 4000 13031
rect 3686 12965 3944 12985
rect 3996 12965 4000 13025
rect 3630 12955 4000 12965
rect 4030 13285 4400 13295
rect 4030 13225 4034 13285
rect 4086 13265 4344 13285
rect 4030 13219 4086 13225
rect 4030 13031 4060 13219
rect 4115 13210 4315 13235
rect 4396 13225 4400 13285
rect 4344 13219 4400 13225
rect 4115 13190 4185 13210
rect 4090 13150 4185 13190
rect 4245 13190 4315 13210
rect 4245 13150 4340 13190
rect 4090 13100 4340 13150
rect 4090 13060 4185 13100
rect 4115 13040 4185 13060
rect 4245 13060 4340 13100
rect 4245 13040 4315 13060
rect 4030 13025 4086 13031
rect 4030 12965 4034 13025
rect 4115 13015 4315 13040
rect 4370 13031 4400 13219
rect 4344 13025 4400 13031
rect 4086 12965 4344 12985
rect 4396 12965 4400 13025
rect 4030 12955 4400 12965
rect 4430 13285 4800 13295
rect 4430 13225 4434 13285
rect 4486 13265 4744 13285
rect 4430 13219 4486 13225
rect 4430 13031 4460 13219
rect 4515 13210 4715 13235
rect 4796 13225 4800 13285
rect 4744 13219 4800 13225
rect 4515 13190 4585 13210
rect 4490 13150 4585 13190
rect 4645 13190 4715 13210
rect 4645 13150 4740 13190
rect 4490 13100 4740 13150
rect 4490 13060 4585 13100
rect 4515 13040 4585 13060
rect 4645 13060 4740 13100
rect 4645 13040 4715 13060
rect 4430 13025 4486 13031
rect 4430 12965 4434 13025
rect 4515 13015 4715 13040
rect 4770 13031 4800 13219
rect 4744 13025 4800 13031
rect 4486 12965 4744 12985
rect 4796 12965 4800 13025
rect 4430 12955 4800 12965
rect 4830 13285 5200 13295
rect 4830 13225 4834 13285
rect 4886 13265 5144 13285
rect 4830 13219 4886 13225
rect 4830 13031 4860 13219
rect 4915 13210 5115 13235
rect 5196 13225 5200 13285
rect 5144 13219 5200 13225
rect 4915 13190 4985 13210
rect 4890 13150 4985 13190
rect 5045 13190 5115 13210
rect 5045 13150 5140 13190
rect 4890 13100 5140 13150
rect 4890 13060 4985 13100
rect 4915 13040 4985 13060
rect 5045 13060 5140 13100
rect 5045 13040 5115 13060
rect 4830 13025 4886 13031
rect 4830 12965 4834 13025
rect 4915 13015 5115 13040
rect 5170 13031 5200 13219
rect 5144 13025 5200 13031
rect 4886 12965 5144 12985
rect 5196 12965 5200 13025
rect 4830 12955 5200 12965
rect 5230 13285 5600 13295
rect 5230 13225 5234 13285
rect 5286 13265 5544 13285
rect 5230 13219 5286 13225
rect 5230 13031 5260 13219
rect 5315 13210 5515 13235
rect 5596 13225 5600 13285
rect 5544 13219 5600 13225
rect 5315 13190 5385 13210
rect 5290 13150 5385 13190
rect 5445 13190 5515 13210
rect 5445 13150 5540 13190
rect 5290 13100 5540 13150
rect 5290 13060 5385 13100
rect 5315 13040 5385 13060
rect 5445 13060 5540 13100
rect 5445 13040 5515 13060
rect 5230 13025 5286 13031
rect 5230 12965 5234 13025
rect 5315 13015 5515 13040
rect 5570 13031 5600 13219
rect 5544 13025 5600 13031
rect 5286 12965 5544 12985
rect 5596 12965 5600 13025
rect 5230 12955 5600 12965
rect 5630 13285 6000 13295
rect 5630 13225 5634 13285
rect 5686 13265 5944 13285
rect 5630 13219 5686 13225
rect 5630 13031 5660 13219
rect 5715 13210 5915 13235
rect 5996 13225 6000 13285
rect 5944 13219 6000 13225
rect 5715 13190 5785 13210
rect 5690 13150 5785 13190
rect 5845 13190 5915 13210
rect 5845 13150 5940 13190
rect 5690 13100 5940 13150
rect 5690 13060 5785 13100
rect 5715 13040 5785 13060
rect 5845 13060 5940 13100
rect 5845 13040 5915 13060
rect 5630 13025 5686 13031
rect 5630 12965 5634 13025
rect 5715 13015 5915 13040
rect 5970 13031 6000 13219
rect 5944 13025 6000 13031
rect 5686 12965 5944 12985
rect 5996 12965 6000 13025
rect 5630 12955 6000 12965
rect 6030 13285 6400 13295
rect 6030 13225 6034 13285
rect 6086 13265 6344 13285
rect 6030 13219 6086 13225
rect 6030 13031 6060 13219
rect 6115 13210 6315 13235
rect 6396 13225 6400 13285
rect 6344 13219 6400 13225
rect 6115 13190 6185 13210
rect 6090 13150 6185 13190
rect 6245 13190 6315 13210
rect 6245 13150 6340 13190
rect 6090 13100 6340 13150
rect 6090 13060 6185 13100
rect 6115 13040 6185 13060
rect 6245 13060 6340 13100
rect 6245 13040 6315 13060
rect 6030 13025 6086 13031
rect 6030 12965 6034 13025
rect 6115 13015 6315 13040
rect 6370 13031 6400 13219
rect 6344 13025 6400 13031
rect 6086 12965 6344 12985
rect 6396 12965 6400 13025
rect 6030 12955 6400 12965
rect 6430 13285 6800 13295
rect 6430 13225 6434 13285
rect 6486 13265 6744 13285
rect 6430 13219 6486 13225
rect 6430 13031 6460 13219
rect 6515 13210 6715 13235
rect 6796 13225 6800 13285
rect 6744 13219 6800 13225
rect 6515 13190 6585 13210
rect 6490 13150 6585 13190
rect 6645 13190 6715 13210
rect 6645 13150 6740 13190
rect 6490 13100 6740 13150
rect 6490 13060 6585 13100
rect 6515 13040 6585 13060
rect 6645 13060 6740 13100
rect 6645 13040 6715 13060
rect 6430 13025 6486 13031
rect 6430 12965 6434 13025
rect 6515 13015 6715 13040
rect 6770 13031 6800 13219
rect 6744 13025 6800 13031
rect 6486 12965 6744 12985
rect 6796 12965 6800 13025
rect 6430 12955 6800 12965
rect 6830 13285 7200 13295
rect 6830 13225 6834 13285
rect 6886 13265 7144 13285
rect 6830 13219 6886 13225
rect 6830 13031 6860 13219
rect 6915 13210 7115 13235
rect 7196 13225 7200 13285
rect 7144 13219 7200 13225
rect 6915 13190 6985 13210
rect 6890 13150 6985 13190
rect 7045 13190 7115 13210
rect 7045 13150 7140 13190
rect 6890 13100 7140 13150
rect 6890 13060 6985 13100
rect 6915 13040 6985 13060
rect 7045 13060 7140 13100
rect 7045 13040 7115 13060
rect 6830 13025 6886 13031
rect 6830 12965 6834 13025
rect 6915 13015 7115 13040
rect 7170 13031 7200 13219
rect 7144 13025 7200 13031
rect 6886 12965 7144 12985
rect 7196 12965 7200 13025
rect 6830 12955 7200 12965
rect 7230 13285 7600 13295
rect 7230 13225 7234 13285
rect 7286 13265 7544 13285
rect 7230 13219 7286 13225
rect 7230 13031 7260 13219
rect 7315 13210 7515 13235
rect 7596 13225 7600 13285
rect 7544 13219 7600 13225
rect 7315 13190 7385 13210
rect 7290 13150 7385 13190
rect 7445 13190 7515 13210
rect 7445 13150 7540 13190
rect 7290 13100 7540 13150
rect 7290 13060 7385 13100
rect 7315 13040 7385 13060
rect 7445 13060 7540 13100
rect 7445 13040 7515 13060
rect 7230 13025 7286 13031
rect 7230 12965 7234 13025
rect 7315 13015 7515 13040
rect 7570 13031 7600 13219
rect 7544 13025 7600 13031
rect 7286 12965 7544 12985
rect 7596 12965 7600 13025
rect 7230 12955 7600 12965
rect 7630 13285 8000 13295
rect 7630 13225 7634 13285
rect 7686 13265 7944 13285
rect 7630 13219 7686 13225
rect 7630 13031 7660 13219
rect 7715 13210 7915 13235
rect 7996 13225 8000 13285
rect 7944 13219 8000 13225
rect 7715 13190 7785 13210
rect 7690 13150 7785 13190
rect 7845 13190 7915 13210
rect 7845 13150 7940 13190
rect 7690 13100 7940 13150
rect 7690 13060 7785 13100
rect 7715 13040 7785 13060
rect 7845 13060 7940 13100
rect 7845 13040 7915 13060
rect 7630 13025 7686 13031
rect 7630 12965 7634 13025
rect 7715 13015 7915 13040
rect 7970 13031 8000 13219
rect 7944 13025 8000 13031
rect 7686 12965 7944 12985
rect 7996 12965 8000 13025
rect 7630 12955 8000 12965
rect 8030 13285 8400 13295
rect 8030 13225 8034 13285
rect 8086 13265 8344 13285
rect 8030 13219 8086 13225
rect 8030 13031 8060 13219
rect 8115 13210 8315 13235
rect 8396 13225 8400 13285
rect 8344 13219 8400 13225
rect 8115 13190 8185 13210
rect 8090 13150 8185 13190
rect 8245 13190 8315 13210
rect 8245 13150 8340 13190
rect 8090 13100 8340 13150
rect 8090 13060 8185 13100
rect 8115 13040 8185 13060
rect 8245 13060 8340 13100
rect 8245 13040 8315 13060
rect 8030 13025 8086 13031
rect 8030 12965 8034 13025
rect 8115 13015 8315 13040
rect 8370 13031 8400 13219
rect 8344 13025 8400 13031
rect 8086 12965 8344 12985
rect 8396 12965 8400 13025
rect 8030 12955 8400 12965
rect 8430 13285 8800 13295
rect 8430 13225 8434 13285
rect 8486 13265 8744 13285
rect 8430 13219 8486 13225
rect 8430 13031 8460 13219
rect 8515 13210 8715 13235
rect 8796 13225 8800 13285
rect 8744 13219 8800 13225
rect 8515 13190 8585 13210
rect 8490 13150 8585 13190
rect 8645 13190 8715 13210
rect 8645 13150 8740 13190
rect 8490 13100 8740 13150
rect 8490 13060 8585 13100
rect 8515 13040 8585 13060
rect 8645 13060 8740 13100
rect 8645 13040 8715 13060
rect 8430 13025 8486 13031
rect 8430 12965 8434 13025
rect 8515 13015 8715 13040
rect 8770 13031 8800 13219
rect 8744 13025 8800 13031
rect 8486 12965 8744 12985
rect 8796 12965 8800 13025
rect 8430 12955 8800 12965
rect 8830 13285 9200 13295
rect 8830 13225 8834 13285
rect 8886 13265 9144 13285
rect 8830 13219 8886 13225
rect 8830 13031 8860 13219
rect 8915 13210 9115 13235
rect 9196 13225 9200 13285
rect 9144 13219 9200 13225
rect 8915 13190 8985 13210
rect 8890 13150 8985 13190
rect 9045 13190 9115 13210
rect 9045 13150 9140 13190
rect 8890 13100 9140 13150
rect 8890 13060 8985 13100
rect 8915 13040 8985 13060
rect 9045 13060 9140 13100
rect 9045 13040 9115 13060
rect 8830 13025 8886 13031
rect 8830 12965 8834 13025
rect 8915 13015 9115 13040
rect 9170 13031 9200 13219
rect 9144 13025 9200 13031
rect 8886 12965 9144 12985
rect 9196 12965 9200 13025
rect 8830 12955 9200 12965
rect 9230 13285 9600 13295
rect 9230 13225 9234 13285
rect 9286 13265 9544 13285
rect 9230 13219 9286 13225
rect 9230 13031 9260 13219
rect 9315 13210 9515 13235
rect 9596 13225 9600 13285
rect 9544 13219 9600 13225
rect 9315 13190 9385 13210
rect 9290 13150 9385 13190
rect 9445 13190 9515 13210
rect 9445 13150 9540 13190
rect 9290 13100 9540 13150
rect 9290 13060 9385 13100
rect 9315 13040 9385 13060
rect 9445 13060 9540 13100
rect 9445 13040 9515 13060
rect 9230 13025 9286 13031
rect 9230 12965 9234 13025
rect 9315 13015 9515 13040
rect 9570 13031 9600 13219
rect 9544 13025 9600 13031
rect 9286 12965 9544 12985
rect 9596 12965 9600 13025
rect 9230 12955 9600 12965
rect 9630 13285 10000 13295
rect 9630 13225 9634 13285
rect 9686 13265 9944 13285
rect 9630 13219 9686 13225
rect 9630 13031 9660 13219
rect 9715 13210 9915 13235
rect 9996 13225 10000 13285
rect 9944 13219 10000 13225
rect 9715 13190 9785 13210
rect 9690 13150 9785 13190
rect 9845 13190 9915 13210
rect 9845 13150 9940 13190
rect 9690 13100 9940 13150
rect 9690 13060 9785 13100
rect 9715 13040 9785 13060
rect 9845 13060 9940 13100
rect 9845 13040 9915 13060
rect 9630 13025 9686 13031
rect 9630 12965 9634 13025
rect 9715 13015 9915 13040
rect 9970 13031 10000 13219
rect 9944 13025 10000 13031
rect 9686 12965 9944 12985
rect 9996 12965 10000 13025
rect 9630 12955 10000 12965
rect 10030 13285 10400 13295
rect 10030 13225 10034 13285
rect 10086 13265 10344 13285
rect 10030 13219 10086 13225
rect 10030 13031 10060 13219
rect 10115 13210 10315 13235
rect 10396 13225 10400 13285
rect 10344 13219 10400 13225
rect 10115 13190 10185 13210
rect 10090 13150 10185 13190
rect 10245 13190 10315 13210
rect 10245 13150 10340 13190
rect 10090 13100 10340 13150
rect 10090 13060 10185 13100
rect 10115 13040 10185 13060
rect 10245 13060 10340 13100
rect 10245 13040 10315 13060
rect 10030 13025 10086 13031
rect 10030 12965 10034 13025
rect 10115 13015 10315 13040
rect 10370 13031 10400 13219
rect 10344 13025 10400 13031
rect 10086 12965 10344 12985
rect 10396 12965 10400 13025
rect 10030 12955 10400 12965
rect 10430 13285 10800 13295
rect 10430 13225 10434 13285
rect 10486 13265 10744 13285
rect 10430 13219 10486 13225
rect 10430 13031 10460 13219
rect 10515 13210 10715 13235
rect 10796 13225 10800 13285
rect 10744 13219 10800 13225
rect 10515 13190 10585 13210
rect 10490 13150 10585 13190
rect 10645 13190 10715 13210
rect 10645 13150 10740 13190
rect 10490 13100 10740 13150
rect 10490 13060 10585 13100
rect 10515 13040 10585 13060
rect 10645 13060 10740 13100
rect 10645 13040 10715 13060
rect 10430 13025 10486 13031
rect 10430 12965 10434 13025
rect 10515 13015 10715 13040
rect 10770 13031 10800 13219
rect 10744 13025 10800 13031
rect 10486 12965 10744 12985
rect 10796 12965 10800 13025
rect 10430 12955 10800 12965
rect 10830 13285 11200 13295
rect 10830 13225 10834 13285
rect 10886 13265 11144 13285
rect 10830 13219 10886 13225
rect 10830 13031 10860 13219
rect 10915 13210 11115 13235
rect 11196 13225 11200 13285
rect 11144 13219 11200 13225
rect 10915 13190 10985 13210
rect 10890 13150 10985 13190
rect 11045 13190 11115 13210
rect 11045 13150 11140 13190
rect 10890 13100 11140 13150
rect 10890 13060 10985 13100
rect 10915 13040 10985 13060
rect 11045 13060 11140 13100
rect 11045 13040 11115 13060
rect 10830 13025 10886 13031
rect 10830 12965 10834 13025
rect 10915 13015 11115 13040
rect 11170 13031 11200 13219
rect 11144 13025 11200 13031
rect 10886 12965 11144 12985
rect 11196 12965 11200 13025
rect 10830 12955 11200 12965
rect 11230 13285 11600 13295
rect 11230 13225 11234 13285
rect 11286 13265 11544 13285
rect 11230 13219 11286 13225
rect 11230 13031 11260 13219
rect 11315 13210 11515 13235
rect 11596 13225 11600 13285
rect 11544 13219 11600 13225
rect 11315 13190 11385 13210
rect 11290 13150 11385 13190
rect 11445 13190 11515 13210
rect 11445 13150 11540 13190
rect 11290 13100 11540 13150
rect 11290 13060 11385 13100
rect 11315 13040 11385 13060
rect 11445 13060 11540 13100
rect 11445 13040 11515 13060
rect 11230 13025 11286 13031
rect 11230 12965 11234 13025
rect 11315 13015 11515 13040
rect 11570 13031 11600 13219
rect 11544 13025 11600 13031
rect 11286 12965 11544 12985
rect 11596 12965 11600 13025
rect 11230 12955 11600 12965
rect 11630 13285 12000 13295
rect 11630 13225 11634 13285
rect 11686 13265 11944 13285
rect 11630 13219 11686 13225
rect 11630 13031 11660 13219
rect 11715 13210 11915 13235
rect 11996 13225 12000 13285
rect 11944 13219 12000 13225
rect 11715 13190 11785 13210
rect 11690 13150 11785 13190
rect 11845 13190 11915 13210
rect 11845 13150 11940 13190
rect 11690 13100 11940 13150
rect 11690 13060 11785 13100
rect 11715 13040 11785 13060
rect 11845 13060 11940 13100
rect 11845 13040 11915 13060
rect 11630 13025 11686 13031
rect 11630 12965 11634 13025
rect 11715 13015 11915 13040
rect 11970 13031 12000 13219
rect 11944 13025 12000 13031
rect 11686 12965 11944 12985
rect 11996 12965 12000 13025
rect 11630 12955 12000 12965
rect 12030 13285 12400 13295
rect 12030 13225 12034 13285
rect 12086 13265 12344 13285
rect 12030 13219 12086 13225
rect 12030 13031 12060 13219
rect 12115 13210 12315 13235
rect 12396 13225 12400 13285
rect 12344 13219 12400 13225
rect 12115 13190 12185 13210
rect 12090 13150 12185 13190
rect 12245 13190 12315 13210
rect 12245 13150 12340 13190
rect 12090 13100 12340 13150
rect 12090 13060 12185 13100
rect 12115 13040 12185 13060
rect 12245 13060 12340 13100
rect 12245 13040 12315 13060
rect 12030 13025 12086 13031
rect 12030 12965 12034 13025
rect 12115 13015 12315 13040
rect 12370 13031 12400 13219
rect 12344 13025 12400 13031
rect 12086 12965 12344 12985
rect 12396 12965 12400 13025
rect 12030 12955 12400 12965
rect 12430 13285 12800 13295
rect 12430 13225 12434 13285
rect 12486 13265 12744 13285
rect 12430 13219 12486 13225
rect 12430 13031 12460 13219
rect 12515 13210 12715 13235
rect 12796 13225 12800 13285
rect 12744 13219 12800 13225
rect 12515 13190 12585 13210
rect 12490 13150 12585 13190
rect 12645 13190 12715 13210
rect 12645 13150 12740 13190
rect 12490 13100 12740 13150
rect 12490 13060 12585 13100
rect 12515 13040 12585 13060
rect 12645 13060 12740 13100
rect 12645 13040 12715 13060
rect 12430 13025 12486 13031
rect 12430 12965 12434 13025
rect 12515 13015 12715 13040
rect 12770 13031 12800 13219
rect 12744 13025 12800 13031
rect 12486 12965 12744 12985
rect 12796 12965 12800 13025
rect 12430 12955 12800 12965
rect 12830 13285 13200 13295
rect 12830 13225 12834 13285
rect 12886 13265 13144 13285
rect 12830 13219 12886 13225
rect 12830 13031 12860 13219
rect 12915 13210 13115 13235
rect 13196 13225 13200 13285
rect 13144 13219 13200 13225
rect 12915 13190 12985 13210
rect 12890 13150 12985 13190
rect 13045 13190 13115 13210
rect 13045 13150 13140 13190
rect 12890 13100 13140 13150
rect 12890 13060 12985 13100
rect 12915 13040 12985 13060
rect 13045 13060 13140 13100
rect 13045 13040 13115 13060
rect 12830 13025 12886 13031
rect 12830 12965 12834 13025
rect 12915 13015 13115 13040
rect 13170 13031 13200 13219
rect 13144 13025 13200 13031
rect 12886 12965 13144 12985
rect 13196 12965 13200 13025
rect 12830 12955 13200 12965
rect -370 12915 0 12925
rect -370 12855 -366 12915
rect -314 12895 -56 12915
rect -370 12849 -314 12855
rect -370 12661 -340 12849
rect -285 12840 -85 12865
rect -4 12855 0 12915
rect -56 12849 0 12855
rect -285 12820 -215 12840
rect -310 12780 -215 12820
rect -155 12820 -85 12840
rect -155 12780 -60 12820
rect -310 12730 -60 12780
rect -310 12690 -215 12730
rect -285 12670 -215 12690
rect -155 12690 -60 12730
rect -155 12670 -85 12690
rect -370 12655 -314 12661
rect -370 12595 -366 12655
rect -285 12645 -85 12670
rect -30 12661 0 12849
rect -56 12655 0 12661
rect -314 12595 -56 12615
rect -4 12595 0 12655
rect -370 12585 0 12595
rect 30 12915 400 12925
rect 30 12855 34 12915
rect 86 12895 344 12915
rect 30 12849 86 12855
rect 30 12661 60 12849
rect 115 12840 315 12865
rect 396 12855 400 12915
rect 344 12849 400 12855
rect 115 12820 185 12840
rect 90 12780 185 12820
rect 245 12820 315 12840
rect 245 12780 340 12820
rect 90 12730 340 12780
rect 90 12690 185 12730
rect 115 12670 185 12690
rect 245 12690 340 12730
rect 245 12670 315 12690
rect 30 12655 86 12661
rect 30 12595 34 12655
rect 115 12645 315 12670
rect 370 12661 400 12849
rect 344 12655 400 12661
rect 86 12595 344 12615
rect 396 12595 400 12655
rect 30 12585 400 12595
rect 430 12915 800 12925
rect 430 12855 434 12915
rect 486 12895 744 12915
rect 430 12849 486 12855
rect 430 12661 460 12849
rect 515 12840 715 12865
rect 796 12855 800 12915
rect 744 12849 800 12855
rect 515 12820 585 12840
rect 490 12780 585 12820
rect 645 12820 715 12840
rect 645 12780 740 12820
rect 490 12730 740 12780
rect 490 12690 585 12730
rect 515 12670 585 12690
rect 645 12690 740 12730
rect 645 12670 715 12690
rect 430 12655 486 12661
rect 430 12595 434 12655
rect 515 12645 715 12670
rect 770 12661 800 12849
rect 744 12655 800 12661
rect 486 12595 744 12615
rect 796 12595 800 12655
rect 430 12585 800 12595
rect 830 12915 1200 12925
rect 830 12855 834 12915
rect 886 12895 1144 12915
rect 830 12849 886 12855
rect 830 12661 860 12849
rect 915 12840 1115 12865
rect 1196 12855 1200 12915
rect 1144 12849 1200 12855
rect 915 12820 985 12840
rect 890 12780 985 12820
rect 1045 12820 1115 12840
rect 1045 12780 1140 12820
rect 890 12730 1140 12780
rect 890 12690 985 12730
rect 915 12670 985 12690
rect 1045 12690 1140 12730
rect 1045 12670 1115 12690
rect 830 12655 886 12661
rect 830 12595 834 12655
rect 915 12645 1115 12670
rect 1170 12661 1200 12849
rect 1144 12655 1200 12661
rect 886 12595 1144 12615
rect 1196 12595 1200 12655
rect 830 12585 1200 12595
rect 1230 12915 1600 12925
rect 1230 12855 1234 12915
rect 1286 12895 1544 12915
rect 1230 12849 1286 12855
rect 1230 12661 1260 12849
rect 1315 12840 1515 12865
rect 1596 12855 1600 12915
rect 1544 12849 1600 12855
rect 1315 12820 1385 12840
rect 1290 12780 1385 12820
rect 1445 12820 1515 12840
rect 1445 12780 1540 12820
rect 1290 12730 1540 12780
rect 1290 12690 1385 12730
rect 1315 12670 1385 12690
rect 1445 12690 1540 12730
rect 1445 12670 1515 12690
rect 1230 12655 1286 12661
rect 1230 12595 1234 12655
rect 1315 12645 1515 12670
rect 1570 12661 1600 12849
rect 1544 12655 1600 12661
rect 1286 12595 1544 12615
rect 1596 12595 1600 12655
rect 1230 12585 1600 12595
rect 1630 12915 2000 12925
rect 1630 12855 1634 12915
rect 1686 12895 1944 12915
rect 1630 12849 1686 12855
rect 1630 12661 1660 12849
rect 1715 12840 1915 12865
rect 1996 12855 2000 12915
rect 1944 12849 2000 12855
rect 1715 12820 1785 12840
rect 1690 12780 1785 12820
rect 1845 12820 1915 12840
rect 1845 12780 1940 12820
rect 1690 12730 1940 12780
rect 1690 12690 1785 12730
rect 1715 12670 1785 12690
rect 1845 12690 1940 12730
rect 1845 12670 1915 12690
rect 1630 12655 1686 12661
rect 1630 12595 1634 12655
rect 1715 12645 1915 12670
rect 1970 12661 2000 12849
rect 1944 12655 2000 12661
rect 1686 12595 1944 12615
rect 1996 12595 2000 12655
rect 1630 12585 2000 12595
rect 2030 12915 2400 12925
rect 2030 12855 2034 12915
rect 2086 12895 2344 12915
rect 2030 12849 2086 12855
rect 2030 12661 2060 12849
rect 2115 12840 2315 12865
rect 2396 12855 2400 12915
rect 2344 12849 2400 12855
rect 2115 12820 2185 12840
rect 2090 12780 2185 12820
rect 2245 12820 2315 12840
rect 2245 12780 2340 12820
rect 2090 12730 2340 12780
rect 2090 12690 2185 12730
rect 2115 12670 2185 12690
rect 2245 12690 2340 12730
rect 2245 12670 2315 12690
rect 2030 12655 2086 12661
rect 2030 12595 2034 12655
rect 2115 12645 2315 12670
rect 2370 12661 2400 12849
rect 2344 12655 2400 12661
rect 2086 12595 2344 12615
rect 2396 12595 2400 12655
rect 2030 12585 2400 12595
rect 2430 12915 2800 12925
rect 2430 12855 2434 12915
rect 2486 12895 2744 12915
rect 2430 12849 2486 12855
rect 2430 12661 2460 12849
rect 2515 12840 2715 12865
rect 2796 12855 2800 12915
rect 2744 12849 2800 12855
rect 2515 12820 2585 12840
rect 2490 12780 2585 12820
rect 2645 12820 2715 12840
rect 2645 12780 2740 12820
rect 2490 12730 2740 12780
rect 2490 12690 2585 12730
rect 2515 12670 2585 12690
rect 2645 12690 2740 12730
rect 2645 12670 2715 12690
rect 2430 12655 2486 12661
rect 2430 12595 2434 12655
rect 2515 12645 2715 12670
rect 2770 12661 2800 12849
rect 2744 12655 2800 12661
rect 2486 12595 2744 12615
rect 2796 12595 2800 12655
rect 2430 12585 2800 12595
rect 2830 12915 3200 12925
rect 2830 12855 2834 12915
rect 2886 12895 3144 12915
rect 2830 12849 2886 12855
rect 2830 12661 2860 12849
rect 2915 12840 3115 12865
rect 3196 12855 3200 12915
rect 3144 12849 3200 12855
rect 2915 12820 2985 12840
rect 2890 12780 2985 12820
rect 3045 12820 3115 12840
rect 3045 12780 3140 12820
rect 2890 12730 3140 12780
rect 2890 12690 2985 12730
rect 2915 12670 2985 12690
rect 3045 12690 3140 12730
rect 3045 12670 3115 12690
rect 2830 12655 2886 12661
rect 2830 12595 2834 12655
rect 2915 12645 3115 12670
rect 3170 12661 3200 12849
rect 3144 12655 3200 12661
rect 2886 12595 3144 12615
rect 3196 12595 3200 12655
rect 2830 12585 3200 12595
rect 3230 12915 3600 12925
rect 3230 12855 3234 12915
rect 3286 12895 3544 12915
rect 3230 12849 3286 12855
rect 3230 12661 3260 12849
rect 3315 12840 3515 12865
rect 3596 12855 3600 12915
rect 3544 12849 3600 12855
rect 3315 12820 3385 12840
rect 3290 12780 3385 12820
rect 3445 12820 3515 12840
rect 3445 12780 3540 12820
rect 3290 12730 3540 12780
rect 3290 12690 3385 12730
rect 3315 12670 3385 12690
rect 3445 12690 3540 12730
rect 3445 12670 3515 12690
rect 3230 12655 3286 12661
rect 3230 12595 3234 12655
rect 3315 12645 3515 12670
rect 3570 12661 3600 12849
rect 3544 12655 3600 12661
rect 3286 12595 3544 12615
rect 3596 12595 3600 12655
rect 3230 12585 3600 12595
rect 3630 12915 4000 12925
rect 3630 12855 3634 12915
rect 3686 12895 3944 12915
rect 3630 12849 3686 12855
rect 3630 12661 3660 12849
rect 3715 12840 3915 12865
rect 3996 12855 4000 12915
rect 3944 12849 4000 12855
rect 3715 12820 3785 12840
rect 3690 12780 3785 12820
rect 3845 12820 3915 12840
rect 3845 12780 3940 12820
rect 3690 12730 3940 12780
rect 3690 12690 3785 12730
rect 3715 12670 3785 12690
rect 3845 12690 3940 12730
rect 3845 12670 3915 12690
rect 3630 12655 3686 12661
rect 3630 12595 3634 12655
rect 3715 12645 3915 12670
rect 3970 12661 4000 12849
rect 3944 12655 4000 12661
rect 3686 12595 3944 12615
rect 3996 12595 4000 12655
rect 3630 12585 4000 12595
rect 4030 12915 4400 12925
rect 4030 12855 4034 12915
rect 4086 12895 4344 12915
rect 4030 12849 4086 12855
rect 4030 12661 4060 12849
rect 4115 12840 4315 12865
rect 4396 12855 4400 12915
rect 4344 12849 4400 12855
rect 4115 12820 4185 12840
rect 4090 12780 4185 12820
rect 4245 12820 4315 12840
rect 4245 12780 4340 12820
rect 4090 12730 4340 12780
rect 4090 12690 4185 12730
rect 4115 12670 4185 12690
rect 4245 12690 4340 12730
rect 4245 12670 4315 12690
rect 4030 12655 4086 12661
rect 4030 12595 4034 12655
rect 4115 12645 4315 12670
rect 4370 12661 4400 12849
rect 4344 12655 4400 12661
rect 4086 12595 4344 12615
rect 4396 12595 4400 12655
rect 4030 12585 4400 12595
rect 4430 12915 4800 12925
rect 4430 12855 4434 12915
rect 4486 12895 4744 12915
rect 4430 12849 4486 12855
rect 4430 12661 4460 12849
rect 4515 12840 4715 12865
rect 4796 12855 4800 12915
rect 4744 12849 4800 12855
rect 4515 12820 4585 12840
rect 4490 12780 4585 12820
rect 4645 12820 4715 12840
rect 4645 12780 4740 12820
rect 4490 12730 4740 12780
rect 4490 12690 4585 12730
rect 4515 12670 4585 12690
rect 4645 12690 4740 12730
rect 4645 12670 4715 12690
rect 4430 12655 4486 12661
rect 4430 12595 4434 12655
rect 4515 12645 4715 12670
rect 4770 12661 4800 12849
rect 4744 12655 4800 12661
rect 4486 12595 4744 12615
rect 4796 12595 4800 12655
rect 4430 12585 4800 12595
rect 4830 12915 5200 12925
rect 4830 12855 4834 12915
rect 4886 12895 5144 12915
rect 4830 12849 4886 12855
rect 4830 12661 4860 12849
rect 4915 12840 5115 12865
rect 5196 12855 5200 12915
rect 5144 12849 5200 12855
rect 4915 12820 4985 12840
rect 4890 12780 4985 12820
rect 5045 12820 5115 12840
rect 5045 12780 5140 12820
rect 4890 12730 5140 12780
rect 4890 12690 4985 12730
rect 4915 12670 4985 12690
rect 5045 12690 5140 12730
rect 5045 12670 5115 12690
rect 4830 12655 4886 12661
rect 4830 12595 4834 12655
rect 4915 12645 5115 12670
rect 5170 12661 5200 12849
rect 5144 12655 5200 12661
rect 4886 12595 5144 12615
rect 5196 12595 5200 12655
rect 4830 12585 5200 12595
rect 5230 12915 5600 12925
rect 5230 12855 5234 12915
rect 5286 12895 5544 12915
rect 5230 12849 5286 12855
rect 5230 12661 5260 12849
rect 5315 12840 5515 12865
rect 5596 12855 5600 12915
rect 5544 12849 5600 12855
rect 5315 12820 5385 12840
rect 5290 12780 5385 12820
rect 5445 12820 5515 12840
rect 5445 12780 5540 12820
rect 5290 12730 5540 12780
rect 5290 12690 5385 12730
rect 5315 12670 5385 12690
rect 5445 12690 5540 12730
rect 5445 12670 5515 12690
rect 5230 12655 5286 12661
rect 5230 12595 5234 12655
rect 5315 12645 5515 12670
rect 5570 12661 5600 12849
rect 5544 12655 5600 12661
rect 5286 12595 5544 12615
rect 5596 12595 5600 12655
rect 5230 12585 5600 12595
rect 5630 12915 6000 12925
rect 5630 12855 5634 12915
rect 5686 12895 5944 12915
rect 5630 12849 5686 12855
rect 5630 12661 5660 12849
rect 5715 12840 5915 12865
rect 5996 12855 6000 12915
rect 5944 12849 6000 12855
rect 5715 12820 5785 12840
rect 5690 12780 5785 12820
rect 5845 12820 5915 12840
rect 5845 12780 5940 12820
rect 5690 12730 5940 12780
rect 5690 12690 5785 12730
rect 5715 12670 5785 12690
rect 5845 12690 5940 12730
rect 5845 12670 5915 12690
rect 5630 12655 5686 12661
rect 5630 12595 5634 12655
rect 5715 12645 5915 12670
rect 5970 12661 6000 12849
rect 5944 12655 6000 12661
rect 5686 12595 5944 12615
rect 5996 12595 6000 12655
rect 5630 12585 6000 12595
rect 6030 12915 6400 12925
rect 6030 12855 6034 12915
rect 6086 12895 6344 12915
rect 6030 12849 6086 12855
rect 6030 12661 6060 12849
rect 6115 12840 6315 12865
rect 6396 12855 6400 12915
rect 6344 12849 6400 12855
rect 6115 12820 6185 12840
rect 6090 12780 6185 12820
rect 6245 12820 6315 12840
rect 6245 12780 6340 12820
rect 6090 12730 6340 12780
rect 6090 12690 6185 12730
rect 6115 12670 6185 12690
rect 6245 12690 6340 12730
rect 6245 12670 6315 12690
rect 6030 12655 6086 12661
rect 6030 12595 6034 12655
rect 6115 12645 6315 12670
rect 6370 12661 6400 12849
rect 6344 12655 6400 12661
rect 6086 12595 6344 12615
rect 6396 12595 6400 12655
rect 6030 12585 6400 12595
rect 6430 12915 6800 12925
rect 6430 12855 6434 12915
rect 6486 12895 6744 12915
rect 6430 12849 6486 12855
rect 6430 12661 6460 12849
rect 6515 12840 6715 12865
rect 6796 12855 6800 12915
rect 6744 12849 6800 12855
rect 6515 12820 6585 12840
rect 6490 12780 6585 12820
rect 6645 12820 6715 12840
rect 6645 12780 6740 12820
rect 6490 12730 6740 12780
rect 6490 12690 6585 12730
rect 6515 12670 6585 12690
rect 6645 12690 6740 12730
rect 6645 12670 6715 12690
rect 6430 12655 6486 12661
rect 6430 12595 6434 12655
rect 6515 12645 6715 12670
rect 6770 12661 6800 12849
rect 6744 12655 6800 12661
rect 6486 12595 6744 12615
rect 6796 12595 6800 12655
rect 6430 12585 6800 12595
rect 6830 12915 7200 12925
rect 6830 12855 6834 12915
rect 6886 12895 7144 12915
rect 6830 12849 6886 12855
rect 6830 12661 6860 12849
rect 6915 12840 7115 12865
rect 7196 12855 7200 12915
rect 7144 12849 7200 12855
rect 6915 12820 6985 12840
rect 6890 12780 6985 12820
rect 7045 12820 7115 12840
rect 7045 12780 7140 12820
rect 6890 12730 7140 12780
rect 6890 12690 6985 12730
rect 6915 12670 6985 12690
rect 7045 12690 7140 12730
rect 7045 12670 7115 12690
rect 6830 12655 6886 12661
rect 6830 12595 6834 12655
rect 6915 12645 7115 12670
rect 7170 12661 7200 12849
rect 7144 12655 7200 12661
rect 6886 12595 7144 12615
rect 7196 12595 7200 12655
rect 6830 12585 7200 12595
rect 7230 12915 7600 12925
rect 7230 12855 7234 12915
rect 7286 12895 7544 12915
rect 7230 12849 7286 12855
rect 7230 12661 7260 12849
rect 7315 12840 7515 12865
rect 7596 12855 7600 12915
rect 7544 12849 7600 12855
rect 7315 12820 7385 12840
rect 7290 12780 7385 12820
rect 7445 12820 7515 12840
rect 7445 12780 7540 12820
rect 7290 12730 7540 12780
rect 7290 12690 7385 12730
rect 7315 12670 7385 12690
rect 7445 12690 7540 12730
rect 7445 12670 7515 12690
rect 7230 12655 7286 12661
rect 7230 12595 7234 12655
rect 7315 12645 7515 12670
rect 7570 12661 7600 12849
rect 7544 12655 7600 12661
rect 7286 12595 7544 12615
rect 7596 12595 7600 12655
rect 7230 12585 7600 12595
rect 7630 12915 8000 12925
rect 7630 12855 7634 12915
rect 7686 12895 7944 12915
rect 7630 12849 7686 12855
rect 7630 12661 7660 12849
rect 7715 12840 7915 12865
rect 7996 12855 8000 12915
rect 7944 12849 8000 12855
rect 7715 12820 7785 12840
rect 7690 12780 7785 12820
rect 7845 12820 7915 12840
rect 7845 12780 7940 12820
rect 7690 12730 7940 12780
rect 7690 12690 7785 12730
rect 7715 12670 7785 12690
rect 7845 12690 7940 12730
rect 7845 12670 7915 12690
rect 7630 12655 7686 12661
rect 7630 12595 7634 12655
rect 7715 12645 7915 12670
rect 7970 12661 8000 12849
rect 7944 12655 8000 12661
rect 7686 12595 7944 12615
rect 7996 12595 8000 12655
rect 7630 12585 8000 12595
rect 8030 12915 8400 12925
rect 8030 12855 8034 12915
rect 8086 12895 8344 12915
rect 8030 12849 8086 12855
rect 8030 12661 8060 12849
rect 8115 12840 8315 12865
rect 8396 12855 8400 12915
rect 8344 12849 8400 12855
rect 8115 12820 8185 12840
rect 8090 12780 8185 12820
rect 8245 12820 8315 12840
rect 8245 12780 8340 12820
rect 8090 12730 8340 12780
rect 8090 12690 8185 12730
rect 8115 12670 8185 12690
rect 8245 12690 8340 12730
rect 8245 12670 8315 12690
rect 8030 12655 8086 12661
rect 8030 12595 8034 12655
rect 8115 12645 8315 12670
rect 8370 12661 8400 12849
rect 8344 12655 8400 12661
rect 8086 12595 8344 12615
rect 8396 12595 8400 12655
rect 8030 12585 8400 12595
rect 8430 12915 8800 12925
rect 8430 12855 8434 12915
rect 8486 12895 8744 12915
rect 8430 12849 8486 12855
rect 8430 12661 8460 12849
rect 8515 12840 8715 12865
rect 8796 12855 8800 12915
rect 8744 12849 8800 12855
rect 8515 12820 8585 12840
rect 8490 12780 8585 12820
rect 8645 12820 8715 12840
rect 8645 12780 8740 12820
rect 8490 12730 8740 12780
rect 8490 12690 8585 12730
rect 8515 12670 8585 12690
rect 8645 12690 8740 12730
rect 8645 12670 8715 12690
rect 8430 12655 8486 12661
rect 8430 12595 8434 12655
rect 8515 12645 8715 12670
rect 8770 12661 8800 12849
rect 8744 12655 8800 12661
rect 8486 12595 8744 12615
rect 8796 12595 8800 12655
rect 8430 12585 8800 12595
rect 8830 12915 9200 12925
rect 8830 12855 8834 12915
rect 8886 12895 9144 12915
rect 8830 12849 8886 12855
rect 8830 12661 8860 12849
rect 8915 12840 9115 12865
rect 9196 12855 9200 12915
rect 9144 12849 9200 12855
rect 8915 12820 8985 12840
rect 8890 12780 8985 12820
rect 9045 12820 9115 12840
rect 9045 12780 9140 12820
rect 8890 12730 9140 12780
rect 8890 12690 8985 12730
rect 8915 12670 8985 12690
rect 9045 12690 9140 12730
rect 9045 12670 9115 12690
rect 8830 12655 8886 12661
rect 8830 12595 8834 12655
rect 8915 12645 9115 12670
rect 9170 12661 9200 12849
rect 9144 12655 9200 12661
rect 8886 12595 9144 12615
rect 9196 12595 9200 12655
rect 8830 12585 9200 12595
rect 9230 12915 9600 12925
rect 9230 12855 9234 12915
rect 9286 12895 9544 12915
rect 9230 12849 9286 12855
rect 9230 12661 9260 12849
rect 9315 12840 9515 12865
rect 9596 12855 9600 12915
rect 9544 12849 9600 12855
rect 9315 12820 9385 12840
rect 9290 12780 9385 12820
rect 9445 12820 9515 12840
rect 9445 12780 9540 12820
rect 9290 12730 9540 12780
rect 9290 12690 9385 12730
rect 9315 12670 9385 12690
rect 9445 12690 9540 12730
rect 9445 12670 9515 12690
rect 9230 12655 9286 12661
rect 9230 12595 9234 12655
rect 9315 12645 9515 12670
rect 9570 12661 9600 12849
rect 9544 12655 9600 12661
rect 9286 12595 9544 12615
rect 9596 12595 9600 12655
rect 9230 12585 9600 12595
rect 9630 12915 10000 12925
rect 9630 12855 9634 12915
rect 9686 12895 9944 12915
rect 9630 12849 9686 12855
rect 9630 12661 9660 12849
rect 9715 12840 9915 12865
rect 9996 12855 10000 12915
rect 9944 12849 10000 12855
rect 9715 12820 9785 12840
rect 9690 12780 9785 12820
rect 9845 12820 9915 12840
rect 9845 12780 9940 12820
rect 9690 12730 9940 12780
rect 9690 12690 9785 12730
rect 9715 12670 9785 12690
rect 9845 12690 9940 12730
rect 9845 12670 9915 12690
rect 9630 12655 9686 12661
rect 9630 12595 9634 12655
rect 9715 12645 9915 12670
rect 9970 12661 10000 12849
rect 9944 12655 10000 12661
rect 9686 12595 9944 12615
rect 9996 12595 10000 12655
rect 9630 12585 10000 12595
rect 10030 12915 10400 12925
rect 10030 12855 10034 12915
rect 10086 12895 10344 12915
rect 10030 12849 10086 12855
rect 10030 12661 10060 12849
rect 10115 12840 10315 12865
rect 10396 12855 10400 12915
rect 10344 12849 10400 12855
rect 10115 12820 10185 12840
rect 10090 12780 10185 12820
rect 10245 12820 10315 12840
rect 10245 12780 10340 12820
rect 10090 12730 10340 12780
rect 10090 12690 10185 12730
rect 10115 12670 10185 12690
rect 10245 12690 10340 12730
rect 10245 12670 10315 12690
rect 10030 12655 10086 12661
rect 10030 12595 10034 12655
rect 10115 12645 10315 12670
rect 10370 12661 10400 12849
rect 10344 12655 10400 12661
rect 10086 12595 10344 12615
rect 10396 12595 10400 12655
rect 10030 12585 10400 12595
rect 10430 12915 10800 12925
rect 10430 12855 10434 12915
rect 10486 12895 10744 12915
rect 10430 12849 10486 12855
rect 10430 12661 10460 12849
rect 10515 12840 10715 12865
rect 10796 12855 10800 12915
rect 10744 12849 10800 12855
rect 10515 12820 10585 12840
rect 10490 12780 10585 12820
rect 10645 12820 10715 12840
rect 10645 12780 10740 12820
rect 10490 12730 10740 12780
rect 10490 12690 10585 12730
rect 10515 12670 10585 12690
rect 10645 12690 10740 12730
rect 10645 12670 10715 12690
rect 10430 12655 10486 12661
rect 10430 12595 10434 12655
rect 10515 12645 10715 12670
rect 10770 12661 10800 12849
rect 10744 12655 10800 12661
rect 10486 12595 10744 12615
rect 10796 12595 10800 12655
rect 10430 12585 10800 12595
rect 10830 12915 11200 12925
rect 10830 12855 10834 12915
rect 10886 12895 11144 12915
rect 10830 12849 10886 12855
rect 10830 12661 10860 12849
rect 10915 12840 11115 12865
rect 11196 12855 11200 12915
rect 11144 12849 11200 12855
rect 10915 12820 10985 12840
rect 10890 12780 10985 12820
rect 11045 12820 11115 12840
rect 11045 12780 11140 12820
rect 10890 12730 11140 12780
rect 10890 12690 10985 12730
rect 10915 12670 10985 12690
rect 11045 12690 11140 12730
rect 11045 12670 11115 12690
rect 10830 12655 10886 12661
rect 10830 12595 10834 12655
rect 10915 12645 11115 12670
rect 11170 12661 11200 12849
rect 11144 12655 11200 12661
rect 10886 12595 11144 12615
rect 11196 12595 11200 12655
rect 10830 12585 11200 12595
rect 11230 12915 11600 12925
rect 11230 12855 11234 12915
rect 11286 12895 11544 12915
rect 11230 12849 11286 12855
rect 11230 12661 11260 12849
rect 11315 12840 11515 12865
rect 11596 12855 11600 12915
rect 11544 12849 11600 12855
rect 11315 12820 11385 12840
rect 11290 12780 11385 12820
rect 11445 12820 11515 12840
rect 11445 12780 11540 12820
rect 11290 12730 11540 12780
rect 11290 12690 11385 12730
rect 11315 12670 11385 12690
rect 11445 12690 11540 12730
rect 11445 12670 11515 12690
rect 11230 12655 11286 12661
rect 11230 12595 11234 12655
rect 11315 12645 11515 12670
rect 11570 12661 11600 12849
rect 11544 12655 11600 12661
rect 11286 12595 11544 12615
rect 11596 12595 11600 12655
rect 11230 12585 11600 12595
rect 11630 12915 12000 12925
rect 11630 12855 11634 12915
rect 11686 12895 11944 12915
rect 11630 12849 11686 12855
rect 11630 12661 11660 12849
rect 11715 12840 11915 12865
rect 11996 12855 12000 12915
rect 11944 12849 12000 12855
rect 11715 12820 11785 12840
rect 11690 12780 11785 12820
rect 11845 12820 11915 12840
rect 11845 12780 11940 12820
rect 11690 12730 11940 12780
rect 11690 12690 11785 12730
rect 11715 12670 11785 12690
rect 11845 12690 11940 12730
rect 11845 12670 11915 12690
rect 11630 12655 11686 12661
rect 11630 12595 11634 12655
rect 11715 12645 11915 12670
rect 11970 12661 12000 12849
rect 11944 12655 12000 12661
rect 11686 12595 11944 12615
rect 11996 12595 12000 12655
rect 11630 12585 12000 12595
rect 12030 12915 12400 12925
rect 12030 12855 12034 12915
rect 12086 12895 12344 12915
rect 12030 12849 12086 12855
rect 12030 12661 12060 12849
rect 12115 12840 12315 12865
rect 12396 12855 12400 12915
rect 12344 12849 12400 12855
rect 12115 12820 12185 12840
rect 12090 12780 12185 12820
rect 12245 12820 12315 12840
rect 12245 12780 12340 12820
rect 12090 12730 12340 12780
rect 12090 12690 12185 12730
rect 12115 12670 12185 12690
rect 12245 12690 12340 12730
rect 12245 12670 12315 12690
rect 12030 12655 12086 12661
rect 12030 12595 12034 12655
rect 12115 12645 12315 12670
rect 12370 12661 12400 12849
rect 12344 12655 12400 12661
rect 12086 12595 12344 12615
rect 12396 12595 12400 12655
rect 12030 12585 12400 12595
rect 12430 12915 12800 12925
rect 12430 12855 12434 12915
rect 12486 12895 12744 12915
rect 12430 12849 12486 12855
rect 12430 12661 12460 12849
rect 12515 12840 12715 12865
rect 12796 12855 12800 12915
rect 12744 12849 12800 12855
rect 12515 12820 12585 12840
rect 12490 12780 12585 12820
rect 12645 12820 12715 12840
rect 12645 12780 12740 12820
rect 12490 12730 12740 12780
rect 12490 12690 12585 12730
rect 12515 12670 12585 12690
rect 12645 12690 12740 12730
rect 12645 12670 12715 12690
rect 12430 12655 12486 12661
rect 12430 12595 12434 12655
rect 12515 12645 12715 12670
rect 12770 12661 12800 12849
rect 12744 12655 12800 12661
rect 12486 12595 12744 12615
rect 12796 12595 12800 12655
rect 12430 12585 12800 12595
rect 12830 12915 13200 12925
rect 12830 12855 12834 12915
rect 12886 12895 13144 12915
rect 12830 12849 12886 12855
rect 12830 12661 12860 12849
rect 12915 12840 13115 12865
rect 13196 12855 13200 12915
rect 13144 12849 13200 12855
rect 12915 12820 12985 12840
rect 12890 12780 12985 12820
rect 13045 12820 13115 12840
rect 13045 12780 13140 12820
rect 12890 12730 13140 12780
rect 12890 12690 12985 12730
rect 12915 12670 12985 12690
rect 13045 12690 13140 12730
rect 13045 12670 13115 12690
rect 12830 12655 12886 12661
rect 12830 12595 12834 12655
rect 12915 12645 13115 12670
rect 13170 12661 13200 12849
rect 13144 12655 13200 12661
rect 12886 12595 13144 12615
rect 13196 12595 13200 12655
rect 12830 12585 13200 12595
rect -370 12545 0 12555
rect -370 12485 -366 12545
rect -314 12525 -56 12545
rect -370 12479 -314 12485
rect -370 12291 -340 12479
rect -285 12470 -85 12495
rect -4 12485 0 12545
rect -56 12479 0 12485
rect -285 12450 -215 12470
rect -310 12410 -215 12450
rect -155 12450 -85 12470
rect -155 12410 -60 12450
rect -310 12360 -60 12410
rect -310 12320 -215 12360
rect -285 12300 -215 12320
rect -155 12320 -60 12360
rect -155 12300 -85 12320
rect -370 12285 -314 12291
rect -370 12225 -366 12285
rect -285 12275 -85 12300
rect -30 12291 0 12479
rect -56 12285 0 12291
rect -314 12225 -56 12245
rect -4 12225 0 12285
rect -370 12215 0 12225
rect 30 12545 400 12555
rect 30 12485 34 12545
rect 86 12525 344 12545
rect 30 12479 86 12485
rect 30 12291 60 12479
rect 115 12470 315 12495
rect 396 12485 400 12545
rect 344 12479 400 12485
rect 115 12450 185 12470
rect 90 12410 185 12450
rect 245 12450 315 12470
rect 245 12410 340 12450
rect 90 12360 340 12410
rect 90 12320 185 12360
rect 115 12300 185 12320
rect 245 12320 340 12360
rect 245 12300 315 12320
rect 30 12285 86 12291
rect 30 12225 34 12285
rect 115 12275 315 12300
rect 370 12291 400 12479
rect 344 12285 400 12291
rect 86 12225 344 12245
rect 396 12225 400 12285
rect 30 12215 400 12225
rect 430 12545 800 12555
rect 430 12485 434 12545
rect 486 12525 744 12545
rect 430 12479 486 12485
rect 430 12291 460 12479
rect 515 12470 715 12495
rect 796 12485 800 12545
rect 744 12479 800 12485
rect 515 12450 585 12470
rect 490 12410 585 12450
rect 645 12450 715 12470
rect 645 12410 740 12450
rect 490 12360 740 12410
rect 490 12320 585 12360
rect 515 12300 585 12320
rect 645 12320 740 12360
rect 645 12300 715 12320
rect 430 12285 486 12291
rect 430 12225 434 12285
rect 515 12275 715 12300
rect 770 12291 800 12479
rect 744 12285 800 12291
rect 486 12225 744 12245
rect 796 12225 800 12285
rect 430 12215 800 12225
rect 830 12545 1200 12555
rect 830 12485 834 12545
rect 886 12525 1144 12545
rect 830 12479 886 12485
rect 830 12291 860 12479
rect 915 12470 1115 12495
rect 1196 12485 1200 12545
rect 1144 12479 1200 12485
rect 915 12450 985 12470
rect 890 12410 985 12450
rect 1045 12450 1115 12470
rect 1045 12410 1140 12450
rect 890 12360 1140 12410
rect 890 12320 985 12360
rect 915 12300 985 12320
rect 1045 12320 1140 12360
rect 1045 12300 1115 12320
rect 830 12285 886 12291
rect 830 12225 834 12285
rect 915 12275 1115 12300
rect 1170 12291 1200 12479
rect 1144 12285 1200 12291
rect 886 12225 1144 12245
rect 1196 12225 1200 12285
rect 830 12215 1200 12225
rect 1230 12545 1600 12555
rect 1230 12485 1234 12545
rect 1286 12525 1544 12545
rect 1230 12479 1286 12485
rect 1230 12291 1260 12479
rect 1315 12470 1515 12495
rect 1596 12485 1600 12545
rect 1544 12479 1600 12485
rect 1315 12450 1385 12470
rect 1290 12410 1385 12450
rect 1445 12450 1515 12470
rect 1445 12410 1540 12450
rect 1290 12360 1540 12410
rect 1290 12320 1385 12360
rect 1315 12300 1385 12320
rect 1445 12320 1540 12360
rect 1445 12300 1515 12320
rect 1230 12285 1286 12291
rect 1230 12225 1234 12285
rect 1315 12275 1515 12300
rect 1570 12291 1600 12479
rect 1544 12285 1600 12291
rect 1286 12225 1544 12245
rect 1596 12225 1600 12285
rect 1230 12215 1600 12225
rect 1630 12545 2000 12555
rect 1630 12485 1634 12545
rect 1686 12525 1944 12545
rect 1630 12479 1686 12485
rect 1630 12291 1660 12479
rect 1715 12470 1915 12495
rect 1996 12485 2000 12545
rect 1944 12479 2000 12485
rect 1715 12450 1785 12470
rect 1690 12410 1785 12450
rect 1845 12450 1915 12470
rect 1845 12410 1940 12450
rect 1690 12360 1940 12410
rect 1690 12320 1785 12360
rect 1715 12300 1785 12320
rect 1845 12320 1940 12360
rect 1845 12300 1915 12320
rect 1630 12285 1686 12291
rect 1630 12225 1634 12285
rect 1715 12275 1915 12300
rect 1970 12291 2000 12479
rect 1944 12285 2000 12291
rect 1686 12225 1944 12245
rect 1996 12225 2000 12285
rect 1630 12215 2000 12225
rect 2030 12545 2400 12555
rect 2030 12485 2034 12545
rect 2086 12525 2344 12545
rect 2030 12479 2086 12485
rect 2030 12291 2060 12479
rect 2115 12470 2315 12495
rect 2396 12485 2400 12545
rect 2344 12479 2400 12485
rect 2115 12450 2185 12470
rect 2090 12410 2185 12450
rect 2245 12450 2315 12470
rect 2245 12410 2340 12450
rect 2090 12360 2340 12410
rect 2090 12320 2185 12360
rect 2115 12300 2185 12320
rect 2245 12320 2340 12360
rect 2245 12300 2315 12320
rect 2030 12285 2086 12291
rect 2030 12225 2034 12285
rect 2115 12275 2315 12300
rect 2370 12291 2400 12479
rect 2344 12285 2400 12291
rect 2086 12225 2344 12245
rect 2396 12225 2400 12285
rect 2030 12215 2400 12225
rect 2430 12545 2800 12555
rect 2430 12485 2434 12545
rect 2486 12525 2744 12545
rect 2430 12479 2486 12485
rect 2430 12291 2460 12479
rect 2515 12470 2715 12495
rect 2796 12485 2800 12545
rect 2744 12479 2800 12485
rect 2515 12450 2585 12470
rect 2490 12410 2585 12450
rect 2645 12450 2715 12470
rect 2645 12410 2740 12450
rect 2490 12360 2740 12410
rect 2490 12320 2585 12360
rect 2515 12300 2585 12320
rect 2645 12320 2740 12360
rect 2645 12300 2715 12320
rect 2430 12285 2486 12291
rect 2430 12225 2434 12285
rect 2515 12275 2715 12300
rect 2770 12291 2800 12479
rect 2744 12285 2800 12291
rect 2486 12225 2744 12245
rect 2796 12225 2800 12285
rect 2430 12215 2800 12225
rect 2830 12545 3200 12555
rect 2830 12485 2834 12545
rect 2886 12525 3144 12545
rect 2830 12479 2886 12485
rect 2830 12291 2860 12479
rect 2915 12470 3115 12495
rect 3196 12485 3200 12545
rect 3144 12479 3200 12485
rect 2915 12450 2985 12470
rect 2890 12410 2985 12450
rect 3045 12450 3115 12470
rect 3045 12410 3140 12450
rect 2890 12360 3140 12410
rect 2890 12320 2985 12360
rect 2915 12300 2985 12320
rect 3045 12320 3140 12360
rect 3045 12300 3115 12320
rect 2830 12285 2886 12291
rect 2830 12225 2834 12285
rect 2915 12275 3115 12300
rect 3170 12291 3200 12479
rect 3144 12285 3200 12291
rect 2886 12225 3144 12245
rect 3196 12225 3200 12285
rect 2830 12215 3200 12225
rect 3230 12545 3600 12555
rect 3230 12485 3234 12545
rect 3286 12525 3544 12545
rect 3230 12479 3286 12485
rect 3230 12291 3260 12479
rect 3315 12470 3515 12495
rect 3596 12485 3600 12545
rect 3544 12479 3600 12485
rect 3315 12450 3385 12470
rect 3290 12410 3385 12450
rect 3445 12450 3515 12470
rect 3445 12410 3540 12450
rect 3290 12360 3540 12410
rect 3290 12320 3385 12360
rect 3315 12300 3385 12320
rect 3445 12320 3540 12360
rect 3445 12300 3515 12320
rect 3230 12285 3286 12291
rect 3230 12225 3234 12285
rect 3315 12275 3515 12300
rect 3570 12291 3600 12479
rect 3544 12285 3600 12291
rect 3286 12225 3544 12245
rect 3596 12225 3600 12285
rect 3230 12215 3600 12225
rect 3630 12545 4000 12555
rect 3630 12485 3634 12545
rect 3686 12525 3944 12545
rect 3630 12479 3686 12485
rect 3630 12291 3660 12479
rect 3715 12470 3915 12495
rect 3996 12485 4000 12545
rect 3944 12479 4000 12485
rect 3715 12450 3785 12470
rect 3690 12410 3785 12450
rect 3845 12450 3915 12470
rect 3845 12410 3940 12450
rect 3690 12360 3940 12410
rect 3690 12320 3785 12360
rect 3715 12300 3785 12320
rect 3845 12320 3940 12360
rect 3845 12300 3915 12320
rect 3630 12285 3686 12291
rect 3630 12225 3634 12285
rect 3715 12275 3915 12300
rect 3970 12291 4000 12479
rect 3944 12285 4000 12291
rect 3686 12225 3944 12245
rect 3996 12225 4000 12285
rect 3630 12215 4000 12225
rect 4030 12545 4400 12555
rect 4030 12485 4034 12545
rect 4086 12525 4344 12545
rect 4030 12479 4086 12485
rect 4030 12291 4060 12479
rect 4115 12470 4315 12495
rect 4396 12485 4400 12545
rect 4344 12479 4400 12485
rect 4115 12450 4185 12470
rect 4090 12410 4185 12450
rect 4245 12450 4315 12470
rect 4245 12410 4340 12450
rect 4090 12360 4340 12410
rect 4090 12320 4185 12360
rect 4115 12300 4185 12320
rect 4245 12320 4340 12360
rect 4245 12300 4315 12320
rect 4030 12285 4086 12291
rect 4030 12225 4034 12285
rect 4115 12275 4315 12300
rect 4370 12291 4400 12479
rect 4344 12285 4400 12291
rect 4086 12225 4344 12245
rect 4396 12225 4400 12285
rect 4030 12215 4400 12225
rect 4430 12545 4800 12555
rect 4430 12485 4434 12545
rect 4486 12525 4744 12545
rect 4430 12479 4486 12485
rect 4430 12291 4460 12479
rect 4515 12470 4715 12495
rect 4796 12485 4800 12545
rect 4744 12479 4800 12485
rect 4515 12450 4585 12470
rect 4490 12410 4585 12450
rect 4645 12450 4715 12470
rect 4645 12410 4740 12450
rect 4490 12360 4740 12410
rect 4490 12320 4585 12360
rect 4515 12300 4585 12320
rect 4645 12320 4740 12360
rect 4645 12300 4715 12320
rect 4430 12285 4486 12291
rect 4430 12225 4434 12285
rect 4515 12275 4715 12300
rect 4770 12291 4800 12479
rect 4744 12285 4800 12291
rect 4486 12225 4744 12245
rect 4796 12225 4800 12285
rect 4430 12215 4800 12225
rect 4830 12545 5200 12555
rect 4830 12485 4834 12545
rect 4886 12525 5144 12545
rect 4830 12479 4886 12485
rect 4830 12291 4860 12479
rect 4915 12470 5115 12495
rect 5196 12485 5200 12545
rect 5144 12479 5200 12485
rect 4915 12450 4985 12470
rect 4890 12410 4985 12450
rect 5045 12450 5115 12470
rect 5045 12410 5140 12450
rect 4890 12360 5140 12410
rect 4890 12320 4985 12360
rect 4915 12300 4985 12320
rect 5045 12320 5140 12360
rect 5045 12300 5115 12320
rect 4830 12285 4886 12291
rect 4830 12225 4834 12285
rect 4915 12275 5115 12300
rect 5170 12291 5200 12479
rect 5144 12285 5200 12291
rect 4886 12225 5144 12245
rect 5196 12225 5200 12285
rect 4830 12215 5200 12225
rect 5230 12545 5600 12555
rect 5230 12485 5234 12545
rect 5286 12525 5544 12545
rect 5230 12479 5286 12485
rect 5230 12291 5260 12479
rect 5315 12470 5515 12495
rect 5596 12485 5600 12545
rect 5544 12479 5600 12485
rect 5315 12450 5385 12470
rect 5290 12410 5385 12450
rect 5445 12450 5515 12470
rect 5445 12410 5540 12450
rect 5290 12360 5540 12410
rect 5290 12320 5385 12360
rect 5315 12300 5385 12320
rect 5445 12320 5540 12360
rect 5445 12300 5515 12320
rect 5230 12285 5286 12291
rect 5230 12225 5234 12285
rect 5315 12275 5515 12300
rect 5570 12291 5600 12479
rect 5544 12285 5600 12291
rect 5286 12225 5544 12245
rect 5596 12225 5600 12285
rect 5230 12215 5600 12225
rect 5630 12545 6000 12555
rect 5630 12485 5634 12545
rect 5686 12525 5944 12545
rect 5630 12479 5686 12485
rect 5630 12291 5660 12479
rect 5715 12470 5915 12495
rect 5996 12485 6000 12545
rect 5944 12479 6000 12485
rect 5715 12450 5785 12470
rect 5690 12410 5785 12450
rect 5845 12450 5915 12470
rect 5845 12410 5940 12450
rect 5690 12360 5940 12410
rect 5690 12320 5785 12360
rect 5715 12300 5785 12320
rect 5845 12320 5940 12360
rect 5845 12300 5915 12320
rect 5630 12285 5686 12291
rect 5630 12225 5634 12285
rect 5715 12275 5915 12300
rect 5970 12291 6000 12479
rect 5944 12285 6000 12291
rect 5686 12225 5944 12245
rect 5996 12225 6000 12285
rect 5630 12215 6000 12225
rect 6030 12545 6400 12555
rect 6030 12485 6034 12545
rect 6086 12525 6344 12545
rect 6030 12479 6086 12485
rect 6030 12291 6060 12479
rect 6115 12470 6315 12495
rect 6396 12485 6400 12545
rect 6344 12479 6400 12485
rect 6115 12450 6185 12470
rect 6090 12410 6185 12450
rect 6245 12450 6315 12470
rect 6245 12410 6340 12450
rect 6090 12360 6340 12410
rect 6090 12320 6185 12360
rect 6115 12300 6185 12320
rect 6245 12320 6340 12360
rect 6245 12300 6315 12320
rect 6030 12285 6086 12291
rect 6030 12225 6034 12285
rect 6115 12275 6315 12300
rect 6370 12291 6400 12479
rect 6344 12285 6400 12291
rect 6086 12225 6344 12245
rect 6396 12225 6400 12285
rect 6030 12215 6400 12225
rect 6430 12545 6800 12555
rect 6430 12485 6434 12545
rect 6486 12525 6744 12545
rect 6430 12479 6486 12485
rect 6430 12291 6460 12479
rect 6515 12470 6715 12495
rect 6796 12485 6800 12545
rect 6744 12479 6800 12485
rect 6515 12450 6585 12470
rect 6490 12410 6585 12450
rect 6645 12450 6715 12470
rect 6645 12410 6740 12450
rect 6490 12360 6740 12410
rect 6490 12320 6585 12360
rect 6515 12300 6585 12320
rect 6645 12320 6740 12360
rect 6645 12300 6715 12320
rect 6430 12285 6486 12291
rect 6430 12225 6434 12285
rect 6515 12275 6715 12300
rect 6770 12291 6800 12479
rect 6744 12285 6800 12291
rect 6486 12225 6744 12245
rect 6796 12225 6800 12285
rect 6430 12215 6800 12225
rect 6830 12545 7200 12555
rect 6830 12485 6834 12545
rect 6886 12525 7144 12545
rect 6830 12479 6886 12485
rect 6830 12291 6860 12479
rect 6915 12470 7115 12495
rect 7196 12485 7200 12545
rect 7144 12479 7200 12485
rect 6915 12450 6985 12470
rect 6890 12410 6985 12450
rect 7045 12450 7115 12470
rect 7045 12410 7140 12450
rect 6890 12360 7140 12410
rect 6890 12320 6985 12360
rect 6915 12300 6985 12320
rect 7045 12320 7140 12360
rect 7045 12300 7115 12320
rect 6830 12285 6886 12291
rect 6830 12225 6834 12285
rect 6915 12275 7115 12300
rect 7170 12291 7200 12479
rect 7144 12285 7200 12291
rect 6886 12225 7144 12245
rect 7196 12225 7200 12285
rect 6830 12215 7200 12225
rect 7230 12545 7600 12555
rect 7230 12485 7234 12545
rect 7286 12525 7544 12545
rect 7230 12479 7286 12485
rect 7230 12291 7260 12479
rect 7315 12470 7515 12495
rect 7596 12485 7600 12545
rect 7544 12479 7600 12485
rect 7315 12450 7385 12470
rect 7290 12410 7385 12450
rect 7445 12450 7515 12470
rect 7445 12410 7540 12450
rect 7290 12360 7540 12410
rect 7290 12320 7385 12360
rect 7315 12300 7385 12320
rect 7445 12320 7540 12360
rect 7445 12300 7515 12320
rect 7230 12285 7286 12291
rect 7230 12225 7234 12285
rect 7315 12275 7515 12300
rect 7570 12291 7600 12479
rect 7544 12285 7600 12291
rect 7286 12225 7544 12245
rect 7596 12225 7600 12285
rect 7230 12215 7600 12225
rect 7630 12545 8000 12555
rect 7630 12485 7634 12545
rect 7686 12525 7944 12545
rect 7630 12479 7686 12485
rect 7630 12291 7660 12479
rect 7715 12470 7915 12495
rect 7996 12485 8000 12545
rect 7944 12479 8000 12485
rect 7715 12450 7785 12470
rect 7690 12410 7785 12450
rect 7845 12450 7915 12470
rect 7845 12410 7940 12450
rect 7690 12360 7940 12410
rect 7690 12320 7785 12360
rect 7715 12300 7785 12320
rect 7845 12320 7940 12360
rect 7845 12300 7915 12320
rect 7630 12285 7686 12291
rect 7630 12225 7634 12285
rect 7715 12275 7915 12300
rect 7970 12291 8000 12479
rect 7944 12285 8000 12291
rect 7686 12225 7944 12245
rect 7996 12225 8000 12285
rect 7630 12215 8000 12225
rect 8030 12545 8400 12555
rect 8030 12485 8034 12545
rect 8086 12525 8344 12545
rect 8030 12479 8086 12485
rect 8030 12291 8060 12479
rect 8115 12470 8315 12495
rect 8396 12485 8400 12545
rect 8344 12479 8400 12485
rect 8115 12450 8185 12470
rect 8090 12410 8185 12450
rect 8245 12450 8315 12470
rect 8245 12410 8340 12450
rect 8090 12360 8340 12410
rect 8090 12320 8185 12360
rect 8115 12300 8185 12320
rect 8245 12320 8340 12360
rect 8245 12300 8315 12320
rect 8030 12285 8086 12291
rect 8030 12225 8034 12285
rect 8115 12275 8315 12300
rect 8370 12291 8400 12479
rect 8344 12285 8400 12291
rect 8086 12225 8344 12245
rect 8396 12225 8400 12285
rect 8030 12215 8400 12225
rect 8430 12545 8800 12555
rect 8430 12485 8434 12545
rect 8486 12525 8744 12545
rect 8430 12479 8486 12485
rect 8430 12291 8460 12479
rect 8515 12470 8715 12495
rect 8796 12485 8800 12545
rect 8744 12479 8800 12485
rect 8515 12450 8585 12470
rect 8490 12410 8585 12450
rect 8645 12450 8715 12470
rect 8645 12410 8740 12450
rect 8490 12360 8740 12410
rect 8490 12320 8585 12360
rect 8515 12300 8585 12320
rect 8645 12320 8740 12360
rect 8645 12300 8715 12320
rect 8430 12285 8486 12291
rect 8430 12225 8434 12285
rect 8515 12275 8715 12300
rect 8770 12291 8800 12479
rect 8744 12285 8800 12291
rect 8486 12225 8744 12245
rect 8796 12225 8800 12285
rect 8430 12215 8800 12225
rect 8830 12545 9200 12555
rect 8830 12485 8834 12545
rect 8886 12525 9144 12545
rect 8830 12479 8886 12485
rect 8830 12291 8860 12479
rect 8915 12470 9115 12495
rect 9196 12485 9200 12545
rect 9144 12479 9200 12485
rect 8915 12450 8985 12470
rect 8890 12410 8985 12450
rect 9045 12450 9115 12470
rect 9045 12410 9140 12450
rect 8890 12360 9140 12410
rect 8890 12320 8985 12360
rect 8915 12300 8985 12320
rect 9045 12320 9140 12360
rect 9045 12300 9115 12320
rect 8830 12285 8886 12291
rect 8830 12225 8834 12285
rect 8915 12275 9115 12300
rect 9170 12291 9200 12479
rect 9144 12285 9200 12291
rect 8886 12225 9144 12245
rect 9196 12225 9200 12285
rect 8830 12215 9200 12225
rect 9230 12545 9600 12555
rect 9230 12485 9234 12545
rect 9286 12525 9544 12545
rect 9230 12479 9286 12485
rect 9230 12291 9260 12479
rect 9315 12470 9515 12495
rect 9596 12485 9600 12545
rect 9544 12479 9600 12485
rect 9315 12450 9385 12470
rect 9290 12410 9385 12450
rect 9445 12450 9515 12470
rect 9445 12410 9540 12450
rect 9290 12360 9540 12410
rect 9290 12320 9385 12360
rect 9315 12300 9385 12320
rect 9445 12320 9540 12360
rect 9445 12300 9515 12320
rect 9230 12285 9286 12291
rect 9230 12225 9234 12285
rect 9315 12275 9515 12300
rect 9570 12291 9600 12479
rect 9544 12285 9600 12291
rect 9286 12225 9544 12245
rect 9596 12225 9600 12285
rect 9230 12215 9600 12225
rect 9630 12545 10000 12555
rect 9630 12485 9634 12545
rect 9686 12525 9944 12545
rect 9630 12479 9686 12485
rect 9630 12291 9660 12479
rect 9715 12470 9915 12495
rect 9996 12485 10000 12545
rect 9944 12479 10000 12485
rect 9715 12450 9785 12470
rect 9690 12410 9785 12450
rect 9845 12450 9915 12470
rect 9845 12410 9940 12450
rect 9690 12360 9940 12410
rect 9690 12320 9785 12360
rect 9715 12300 9785 12320
rect 9845 12320 9940 12360
rect 9845 12300 9915 12320
rect 9630 12285 9686 12291
rect 9630 12225 9634 12285
rect 9715 12275 9915 12300
rect 9970 12291 10000 12479
rect 9944 12285 10000 12291
rect 9686 12225 9944 12245
rect 9996 12225 10000 12285
rect 9630 12215 10000 12225
rect 10030 12545 10400 12555
rect 10030 12485 10034 12545
rect 10086 12525 10344 12545
rect 10030 12479 10086 12485
rect 10030 12291 10060 12479
rect 10115 12470 10315 12495
rect 10396 12485 10400 12545
rect 10344 12479 10400 12485
rect 10115 12450 10185 12470
rect 10090 12410 10185 12450
rect 10245 12450 10315 12470
rect 10245 12410 10340 12450
rect 10090 12360 10340 12410
rect 10090 12320 10185 12360
rect 10115 12300 10185 12320
rect 10245 12320 10340 12360
rect 10245 12300 10315 12320
rect 10030 12285 10086 12291
rect 10030 12225 10034 12285
rect 10115 12275 10315 12300
rect 10370 12291 10400 12479
rect 10344 12285 10400 12291
rect 10086 12225 10344 12245
rect 10396 12225 10400 12285
rect 10030 12215 10400 12225
rect 10430 12545 10800 12555
rect 10430 12485 10434 12545
rect 10486 12525 10744 12545
rect 10430 12479 10486 12485
rect 10430 12291 10460 12479
rect 10515 12470 10715 12495
rect 10796 12485 10800 12545
rect 10744 12479 10800 12485
rect 10515 12450 10585 12470
rect 10490 12410 10585 12450
rect 10645 12450 10715 12470
rect 10645 12410 10740 12450
rect 10490 12360 10740 12410
rect 10490 12320 10585 12360
rect 10515 12300 10585 12320
rect 10645 12320 10740 12360
rect 10645 12300 10715 12320
rect 10430 12285 10486 12291
rect 10430 12225 10434 12285
rect 10515 12275 10715 12300
rect 10770 12291 10800 12479
rect 10744 12285 10800 12291
rect 10486 12225 10744 12245
rect 10796 12225 10800 12285
rect 10430 12215 10800 12225
rect 10830 12545 11200 12555
rect 10830 12485 10834 12545
rect 10886 12525 11144 12545
rect 10830 12479 10886 12485
rect 10830 12291 10860 12479
rect 10915 12470 11115 12495
rect 11196 12485 11200 12545
rect 11144 12479 11200 12485
rect 10915 12450 10985 12470
rect 10890 12410 10985 12450
rect 11045 12450 11115 12470
rect 11045 12410 11140 12450
rect 10890 12360 11140 12410
rect 10890 12320 10985 12360
rect 10915 12300 10985 12320
rect 11045 12320 11140 12360
rect 11045 12300 11115 12320
rect 10830 12285 10886 12291
rect 10830 12225 10834 12285
rect 10915 12275 11115 12300
rect 11170 12291 11200 12479
rect 11144 12285 11200 12291
rect 10886 12225 11144 12245
rect 11196 12225 11200 12285
rect 10830 12215 11200 12225
rect 11230 12545 11600 12555
rect 11230 12485 11234 12545
rect 11286 12525 11544 12545
rect 11230 12479 11286 12485
rect 11230 12291 11260 12479
rect 11315 12470 11515 12495
rect 11596 12485 11600 12545
rect 11544 12479 11600 12485
rect 11315 12450 11385 12470
rect 11290 12410 11385 12450
rect 11445 12450 11515 12470
rect 11445 12410 11540 12450
rect 11290 12360 11540 12410
rect 11290 12320 11385 12360
rect 11315 12300 11385 12320
rect 11445 12320 11540 12360
rect 11445 12300 11515 12320
rect 11230 12285 11286 12291
rect 11230 12225 11234 12285
rect 11315 12275 11515 12300
rect 11570 12291 11600 12479
rect 11544 12285 11600 12291
rect 11286 12225 11544 12245
rect 11596 12225 11600 12285
rect 11230 12215 11600 12225
rect 11630 12545 12000 12555
rect 11630 12485 11634 12545
rect 11686 12525 11944 12545
rect 11630 12479 11686 12485
rect 11630 12291 11660 12479
rect 11715 12470 11915 12495
rect 11996 12485 12000 12545
rect 11944 12479 12000 12485
rect 11715 12450 11785 12470
rect 11690 12410 11785 12450
rect 11845 12450 11915 12470
rect 11845 12410 11940 12450
rect 11690 12360 11940 12410
rect 11690 12320 11785 12360
rect 11715 12300 11785 12320
rect 11845 12320 11940 12360
rect 11845 12300 11915 12320
rect 11630 12285 11686 12291
rect 11630 12225 11634 12285
rect 11715 12275 11915 12300
rect 11970 12291 12000 12479
rect 11944 12285 12000 12291
rect 11686 12225 11944 12245
rect 11996 12225 12000 12285
rect 11630 12215 12000 12225
rect 12030 12545 12400 12555
rect 12030 12485 12034 12545
rect 12086 12525 12344 12545
rect 12030 12479 12086 12485
rect 12030 12291 12060 12479
rect 12115 12470 12315 12495
rect 12396 12485 12400 12545
rect 12344 12479 12400 12485
rect 12115 12450 12185 12470
rect 12090 12410 12185 12450
rect 12245 12450 12315 12470
rect 12245 12410 12340 12450
rect 12090 12360 12340 12410
rect 12090 12320 12185 12360
rect 12115 12300 12185 12320
rect 12245 12320 12340 12360
rect 12245 12300 12315 12320
rect 12030 12285 12086 12291
rect 12030 12225 12034 12285
rect 12115 12275 12315 12300
rect 12370 12291 12400 12479
rect 12344 12285 12400 12291
rect 12086 12225 12344 12245
rect 12396 12225 12400 12285
rect 12030 12215 12400 12225
rect 12430 12545 12800 12555
rect 12430 12485 12434 12545
rect 12486 12525 12744 12545
rect 12430 12479 12486 12485
rect 12430 12291 12460 12479
rect 12515 12470 12715 12495
rect 12796 12485 12800 12545
rect 12744 12479 12800 12485
rect 12515 12450 12585 12470
rect 12490 12410 12585 12450
rect 12645 12450 12715 12470
rect 12645 12410 12740 12450
rect 12490 12360 12740 12410
rect 12490 12320 12585 12360
rect 12515 12300 12585 12320
rect 12645 12320 12740 12360
rect 12645 12300 12715 12320
rect 12430 12285 12486 12291
rect 12430 12225 12434 12285
rect 12515 12275 12715 12300
rect 12770 12291 12800 12479
rect 12744 12285 12800 12291
rect 12486 12225 12744 12245
rect 12796 12225 12800 12285
rect 12430 12215 12800 12225
rect 12830 12545 13200 12555
rect 12830 12485 12834 12545
rect 12886 12525 13144 12545
rect 12830 12479 12886 12485
rect 12830 12291 12860 12479
rect 12915 12470 13115 12495
rect 13196 12485 13200 12545
rect 13144 12479 13200 12485
rect 12915 12450 12985 12470
rect 12890 12410 12985 12450
rect 13045 12450 13115 12470
rect 13045 12410 13140 12450
rect 12890 12360 13140 12410
rect 12890 12320 12985 12360
rect 12915 12300 12985 12320
rect 13045 12320 13140 12360
rect 13045 12300 13115 12320
rect 12830 12285 12886 12291
rect 12830 12225 12834 12285
rect 12915 12275 13115 12300
rect 13170 12291 13200 12479
rect 13144 12285 13200 12291
rect 12886 12225 13144 12245
rect 13196 12225 13200 12285
rect 12830 12215 13200 12225
rect -370 12175 0 12185
rect -370 12115 -366 12175
rect -314 12155 -56 12175
rect -370 12109 -314 12115
rect -370 11921 -340 12109
rect -285 12100 -85 12125
rect -4 12115 0 12175
rect -56 12109 0 12115
rect -285 12080 -215 12100
rect -310 12040 -215 12080
rect -155 12080 -85 12100
rect -155 12040 -60 12080
rect -310 11990 -60 12040
rect -310 11950 -215 11990
rect -285 11930 -215 11950
rect -155 11950 -60 11990
rect -155 11930 -85 11950
rect -370 11915 -314 11921
rect -370 11855 -366 11915
rect -285 11905 -85 11930
rect -30 11921 0 12109
rect -56 11915 0 11921
rect -314 11855 -56 11875
rect -4 11855 0 11915
rect -370 11845 0 11855
rect 30 12175 400 12185
rect 30 12115 34 12175
rect 86 12155 344 12175
rect 30 12109 86 12115
rect 30 11921 60 12109
rect 115 12100 315 12125
rect 396 12115 400 12175
rect 344 12109 400 12115
rect 115 12080 185 12100
rect 90 12040 185 12080
rect 245 12080 315 12100
rect 245 12040 340 12080
rect 90 11990 340 12040
rect 90 11950 185 11990
rect 115 11930 185 11950
rect 245 11950 340 11990
rect 245 11930 315 11950
rect 30 11915 86 11921
rect 30 11855 34 11915
rect 115 11905 315 11930
rect 370 11921 400 12109
rect 344 11915 400 11921
rect 86 11855 344 11875
rect 396 11855 400 11915
rect 30 11845 400 11855
rect 430 12175 800 12185
rect 430 12115 434 12175
rect 486 12155 744 12175
rect 430 12109 486 12115
rect 430 11921 460 12109
rect 515 12100 715 12125
rect 796 12115 800 12175
rect 744 12109 800 12115
rect 515 12080 585 12100
rect 490 12040 585 12080
rect 645 12080 715 12100
rect 645 12040 740 12080
rect 490 11990 740 12040
rect 490 11950 585 11990
rect 515 11930 585 11950
rect 645 11950 740 11990
rect 645 11930 715 11950
rect 430 11915 486 11921
rect 430 11855 434 11915
rect 515 11905 715 11930
rect 770 11921 800 12109
rect 744 11915 800 11921
rect 486 11855 744 11875
rect 796 11855 800 11915
rect 430 11845 800 11855
rect 830 12175 1200 12185
rect 830 12115 834 12175
rect 886 12155 1144 12175
rect 830 12109 886 12115
rect 830 11921 860 12109
rect 915 12100 1115 12125
rect 1196 12115 1200 12175
rect 1144 12109 1200 12115
rect 915 12080 985 12100
rect 890 12040 985 12080
rect 1045 12080 1115 12100
rect 1045 12040 1140 12080
rect 890 11990 1140 12040
rect 890 11950 985 11990
rect 915 11930 985 11950
rect 1045 11950 1140 11990
rect 1045 11930 1115 11950
rect 830 11915 886 11921
rect 830 11855 834 11915
rect 915 11905 1115 11930
rect 1170 11921 1200 12109
rect 1144 11915 1200 11921
rect 886 11855 1144 11875
rect 1196 11855 1200 11915
rect 830 11845 1200 11855
rect 1230 12175 1600 12185
rect 1230 12115 1234 12175
rect 1286 12155 1544 12175
rect 1230 12109 1286 12115
rect 1230 11921 1260 12109
rect 1315 12100 1515 12125
rect 1596 12115 1600 12175
rect 1544 12109 1600 12115
rect 1315 12080 1385 12100
rect 1290 12040 1385 12080
rect 1445 12080 1515 12100
rect 1445 12040 1540 12080
rect 1290 11990 1540 12040
rect 1290 11950 1385 11990
rect 1315 11930 1385 11950
rect 1445 11950 1540 11990
rect 1445 11930 1515 11950
rect 1230 11915 1286 11921
rect 1230 11855 1234 11915
rect 1315 11905 1515 11930
rect 1570 11921 1600 12109
rect 1544 11915 1600 11921
rect 1286 11855 1544 11875
rect 1596 11855 1600 11915
rect 1230 11845 1600 11855
rect 1630 12175 2000 12185
rect 1630 12115 1634 12175
rect 1686 12155 1944 12175
rect 1630 12109 1686 12115
rect 1630 11921 1660 12109
rect 1715 12100 1915 12125
rect 1996 12115 2000 12175
rect 1944 12109 2000 12115
rect 1715 12080 1785 12100
rect 1690 12040 1785 12080
rect 1845 12080 1915 12100
rect 1845 12040 1940 12080
rect 1690 11990 1940 12040
rect 1690 11950 1785 11990
rect 1715 11930 1785 11950
rect 1845 11950 1940 11990
rect 1845 11930 1915 11950
rect 1630 11915 1686 11921
rect 1630 11855 1634 11915
rect 1715 11905 1915 11930
rect 1970 11921 2000 12109
rect 1944 11915 2000 11921
rect 1686 11855 1944 11875
rect 1996 11855 2000 11915
rect 1630 11845 2000 11855
rect 2030 12175 2400 12185
rect 2030 12115 2034 12175
rect 2086 12155 2344 12175
rect 2030 12109 2086 12115
rect 2030 11921 2060 12109
rect 2115 12100 2315 12125
rect 2396 12115 2400 12175
rect 2344 12109 2400 12115
rect 2115 12080 2185 12100
rect 2090 12040 2185 12080
rect 2245 12080 2315 12100
rect 2245 12040 2340 12080
rect 2090 11990 2340 12040
rect 2090 11950 2185 11990
rect 2115 11930 2185 11950
rect 2245 11950 2340 11990
rect 2245 11930 2315 11950
rect 2030 11915 2086 11921
rect 2030 11855 2034 11915
rect 2115 11905 2315 11930
rect 2370 11921 2400 12109
rect 2344 11915 2400 11921
rect 2086 11855 2344 11875
rect 2396 11855 2400 11915
rect 2030 11845 2400 11855
rect 2430 12175 2800 12185
rect 2430 12115 2434 12175
rect 2486 12155 2744 12175
rect 2430 12109 2486 12115
rect 2430 11921 2460 12109
rect 2515 12100 2715 12125
rect 2796 12115 2800 12175
rect 2744 12109 2800 12115
rect 2515 12080 2585 12100
rect 2490 12040 2585 12080
rect 2645 12080 2715 12100
rect 2645 12040 2740 12080
rect 2490 11990 2740 12040
rect 2490 11950 2585 11990
rect 2515 11930 2585 11950
rect 2645 11950 2740 11990
rect 2645 11930 2715 11950
rect 2430 11915 2486 11921
rect 2430 11855 2434 11915
rect 2515 11905 2715 11930
rect 2770 11921 2800 12109
rect 2744 11915 2800 11921
rect 2486 11855 2744 11875
rect 2796 11855 2800 11915
rect 2430 11845 2800 11855
rect 2830 12175 3200 12185
rect 2830 12115 2834 12175
rect 2886 12155 3144 12175
rect 2830 12109 2886 12115
rect 2830 11921 2860 12109
rect 2915 12100 3115 12125
rect 3196 12115 3200 12175
rect 3144 12109 3200 12115
rect 2915 12080 2985 12100
rect 2890 12040 2985 12080
rect 3045 12080 3115 12100
rect 3045 12040 3140 12080
rect 2890 11990 3140 12040
rect 2890 11950 2985 11990
rect 2915 11930 2985 11950
rect 3045 11950 3140 11990
rect 3045 11930 3115 11950
rect 2830 11915 2886 11921
rect 2830 11855 2834 11915
rect 2915 11905 3115 11930
rect 3170 11921 3200 12109
rect 3144 11915 3200 11921
rect 2886 11855 3144 11875
rect 3196 11855 3200 11915
rect 2830 11845 3200 11855
rect 3230 12175 3600 12185
rect 3230 12115 3234 12175
rect 3286 12155 3544 12175
rect 3230 12109 3286 12115
rect 3230 11921 3260 12109
rect 3315 12100 3515 12125
rect 3596 12115 3600 12175
rect 3544 12109 3600 12115
rect 3315 12080 3385 12100
rect 3290 12040 3385 12080
rect 3445 12080 3515 12100
rect 3445 12040 3540 12080
rect 3290 11990 3540 12040
rect 3290 11950 3385 11990
rect 3315 11930 3385 11950
rect 3445 11950 3540 11990
rect 3445 11930 3515 11950
rect 3230 11915 3286 11921
rect 3230 11855 3234 11915
rect 3315 11905 3515 11930
rect 3570 11921 3600 12109
rect 3544 11915 3600 11921
rect 3286 11855 3544 11875
rect 3596 11855 3600 11915
rect 3230 11845 3600 11855
rect 3630 12175 4000 12185
rect 3630 12115 3634 12175
rect 3686 12155 3944 12175
rect 3630 12109 3686 12115
rect 3630 11921 3660 12109
rect 3715 12100 3915 12125
rect 3996 12115 4000 12175
rect 3944 12109 4000 12115
rect 3715 12080 3785 12100
rect 3690 12040 3785 12080
rect 3845 12080 3915 12100
rect 3845 12040 3940 12080
rect 3690 11990 3940 12040
rect 3690 11950 3785 11990
rect 3715 11930 3785 11950
rect 3845 11950 3940 11990
rect 3845 11930 3915 11950
rect 3630 11915 3686 11921
rect 3630 11855 3634 11915
rect 3715 11905 3915 11930
rect 3970 11921 4000 12109
rect 3944 11915 4000 11921
rect 3686 11855 3944 11875
rect 3996 11855 4000 11915
rect 3630 11845 4000 11855
rect 4030 12175 4400 12185
rect 4030 12115 4034 12175
rect 4086 12155 4344 12175
rect 4030 12109 4086 12115
rect 4030 11921 4060 12109
rect 4115 12100 4315 12125
rect 4396 12115 4400 12175
rect 4344 12109 4400 12115
rect 4115 12080 4185 12100
rect 4090 12040 4185 12080
rect 4245 12080 4315 12100
rect 4245 12040 4340 12080
rect 4090 11990 4340 12040
rect 4090 11950 4185 11990
rect 4115 11930 4185 11950
rect 4245 11950 4340 11990
rect 4245 11930 4315 11950
rect 4030 11915 4086 11921
rect 4030 11855 4034 11915
rect 4115 11905 4315 11930
rect 4370 11921 4400 12109
rect 4344 11915 4400 11921
rect 4086 11855 4344 11875
rect 4396 11855 4400 11915
rect 4030 11845 4400 11855
rect 4430 12175 4800 12185
rect 4430 12115 4434 12175
rect 4486 12155 4744 12175
rect 4430 12109 4486 12115
rect 4430 11921 4460 12109
rect 4515 12100 4715 12125
rect 4796 12115 4800 12175
rect 4744 12109 4800 12115
rect 4515 12080 4585 12100
rect 4490 12040 4585 12080
rect 4645 12080 4715 12100
rect 4645 12040 4740 12080
rect 4490 11990 4740 12040
rect 4490 11950 4585 11990
rect 4515 11930 4585 11950
rect 4645 11950 4740 11990
rect 4645 11930 4715 11950
rect 4430 11915 4486 11921
rect 4430 11855 4434 11915
rect 4515 11905 4715 11930
rect 4770 11921 4800 12109
rect 4744 11915 4800 11921
rect 4486 11855 4744 11875
rect 4796 11855 4800 11915
rect 4430 11845 4800 11855
rect 4830 12175 5200 12185
rect 4830 12115 4834 12175
rect 4886 12155 5144 12175
rect 4830 12109 4886 12115
rect 4830 11921 4860 12109
rect 4915 12100 5115 12125
rect 5196 12115 5200 12175
rect 5144 12109 5200 12115
rect 4915 12080 4985 12100
rect 4890 12040 4985 12080
rect 5045 12080 5115 12100
rect 5045 12040 5140 12080
rect 4890 11990 5140 12040
rect 4890 11950 4985 11990
rect 4915 11930 4985 11950
rect 5045 11950 5140 11990
rect 5045 11930 5115 11950
rect 4830 11915 4886 11921
rect 4830 11855 4834 11915
rect 4915 11905 5115 11930
rect 5170 11921 5200 12109
rect 5144 11915 5200 11921
rect 4886 11855 5144 11875
rect 5196 11855 5200 11915
rect 4830 11845 5200 11855
rect 5230 12175 5600 12185
rect 5230 12115 5234 12175
rect 5286 12155 5544 12175
rect 5230 12109 5286 12115
rect 5230 11921 5260 12109
rect 5315 12100 5515 12125
rect 5596 12115 5600 12175
rect 5544 12109 5600 12115
rect 5315 12080 5385 12100
rect 5290 12040 5385 12080
rect 5445 12080 5515 12100
rect 5445 12040 5540 12080
rect 5290 11990 5540 12040
rect 5290 11950 5385 11990
rect 5315 11930 5385 11950
rect 5445 11950 5540 11990
rect 5445 11930 5515 11950
rect 5230 11915 5286 11921
rect 5230 11855 5234 11915
rect 5315 11905 5515 11930
rect 5570 11921 5600 12109
rect 5544 11915 5600 11921
rect 5286 11855 5544 11875
rect 5596 11855 5600 11915
rect 5230 11845 5600 11855
rect 5630 12175 6000 12185
rect 5630 12115 5634 12175
rect 5686 12155 5944 12175
rect 5630 12109 5686 12115
rect 5630 11921 5660 12109
rect 5715 12100 5915 12125
rect 5996 12115 6000 12175
rect 5944 12109 6000 12115
rect 5715 12080 5785 12100
rect 5690 12040 5785 12080
rect 5845 12080 5915 12100
rect 5845 12040 5940 12080
rect 5690 11990 5940 12040
rect 5690 11950 5785 11990
rect 5715 11930 5785 11950
rect 5845 11950 5940 11990
rect 5845 11930 5915 11950
rect 5630 11915 5686 11921
rect 5630 11855 5634 11915
rect 5715 11905 5915 11930
rect 5970 11921 6000 12109
rect 5944 11915 6000 11921
rect 5686 11855 5944 11875
rect 5996 11855 6000 11915
rect 5630 11845 6000 11855
rect 6030 12175 6400 12185
rect 6030 12115 6034 12175
rect 6086 12155 6344 12175
rect 6030 12109 6086 12115
rect 6030 11921 6060 12109
rect 6115 12100 6315 12125
rect 6396 12115 6400 12175
rect 6344 12109 6400 12115
rect 6115 12080 6185 12100
rect 6090 12040 6185 12080
rect 6245 12080 6315 12100
rect 6245 12040 6340 12080
rect 6090 11990 6340 12040
rect 6090 11950 6185 11990
rect 6115 11930 6185 11950
rect 6245 11950 6340 11990
rect 6245 11930 6315 11950
rect 6030 11915 6086 11921
rect 6030 11855 6034 11915
rect 6115 11905 6315 11930
rect 6370 11921 6400 12109
rect 6344 11915 6400 11921
rect 6086 11855 6344 11875
rect 6396 11855 6400 11915
rect 6030 11845 6400 11855
rect 6430 12175 6800 12185
rect 6430 12115 6434 12175
rect 6486 12155 6744 12175
rect 6430 12109 6486 12115
rect 6430 11921 6460 12109
rect 6515 12100 6715 12125
rect 6796 12115 6800 12175
rect 6744 12109 6800 12115
rect 6515 12080 6585 12100
rect 6490 12040 6585 12080
rect 6645 12080 6715 12100
rect 6645 12040 6740 12080
rect 6490 11990 6740 12040
rect 6490 11950 6585 11990
rect 6515 11930 6585 11950
rect 6645 11950 6740 11990
rect 6645 11930 6715 11950
rect 6430 11915 6486 11921
rect 6430 11855 6434 11915
rect 6515 11905 6715 11930
rect 6770 11921 6800 12109
rect 6744 11915 6800 11921
rect 6486 11855 6744 11875
rect 6796 11855 6800 11915
rect 6430 11845 6800 11855
rect 6830 12175 7200 12185
rect 6830 12115 6834 12175
rect 6886 12155 7144 12175
rect 6830 12109 6886 12115
rect 6830 11921 6860 12109
rect 6915 12100 7115 12125
rect 7196 12115 7200 12175
rect 7144 12109 7200 12115
rect 6915 12080 6985 12100
rect 6890 12040 6985 12080
rect 7045 12080 7115 12100
rect 7045 12040 7140 12080
rect 6890 11990 7140 12040
rect 6890 11950 6985 11990
rect 6915 11930 6985 11950
rect 7045 11950 7140 11990
rect 7045 11930 7115 11950
rect 6830 11915 6886 11921
rect 6830 11855 6834 11915
rect 6915 11905 7115 11930
rect 7170 11921 7200 12109
rect 7144 11915 7200 11921
rect 6886 11855 7144 11875
rect 7196 11855 7200 11915
rect 6830 11845 7200 11855
rect 7230 12175 7600 12185
rect 7230 12115 7234 12175
rect 7286 12155 7544 12175
rect 7230 12109 7286 12115
rect 7230 11921 7260 12109
rect 7315 12100 7515 12125
rect 7596 12115 7600 12175
rect 7544 12109 7600 12115
rect 7315 12080 7385 12100
rect 7290 12040 7385 12080
rect 7445 12080 7515 12100
rect 7445 12040 7540 12080
rect 7290 11990 7540 12040
rect 7290 11950 7385 11990
rect 7315 11930 7385 11950
rect 7445 11950 7540 11990
rect 7445 11930 7515 11950
rect 7230 11915 7286 11921
rect 7230 11855 7234 11915
rect 7315 11905 7515 11930
rect 7570 11921 7600 12109
rect 7544 11915 7600 11921
rect 7286 11855 7544 11875
rect 7596 11855 7600 11915
rect 7230 11845 7600 11855
rect 7630 12175 8000 12185
rect 7630 12115 7634 12175
rect 7686 12155 7944 12175
rect 7630 12109 7686 12115
rect 7630 11921 7660 12109
rect 7715 12100 7915 12125
rect 7996 12115 8000 12175
rect 7944 12109 8000 12115
rect 7715 12080 7785 12100
rect 7690 12040 7785 12080
rect 7845 12080 7915 12100
rect 7845 12040 7940 12080
rect 7690 11990 7940 12040
rect 7690 11950 7785 11990
rect 7715 11930 7785 11950
rect 7845 11950 7940 11990
rect 7845 11930 7915 11950
rect 7630 11915 7686 11921
rect 7630 11855 7634 11915
rect 7715 11905 7915 11930
rect 7970 11921 8000 12109
rect 7944 11915 8000 11921
rect 7686 11855 7944 11875
rect 7996 11855 8000 11915
rect 7630 11845 8000 11855
rect 8030 12175 8400 12185
rect 8030 12115 8034 12175
rect 8086 12155 8344 12175
rect 8030 12109 8086 12115
rect 8030 11921 8060 12109
rect 8115 12100 8315 12125
rect 8396 12115 8400 12175
rect 8344 12109 8400 12115
rect 8115 12080 8185 12100
rect 8090 12040 8185 12080
rect 8245 12080 8315 12100
rect 8245 12040 8340 12080
rect 8090 11990 8340 12040
rect 8090 11950 8185 11990
rect 8115 11930 8185 11950
rect 8245 11950 8340 11990
rect 8245 11930 8315 11950
rect 8030 11915 8086 11921
rect 8030 11855 8034 11915
rect 8115 11905 8315 11930
rect 8370 11921 8400 12109
rect 8344 11915 8400 11921
rect 8086 11855 8344 11875
rect 8396 11855 8400 11915
rect 8030 11845 8400 11855
rect 8430 12175 8800 12185
rect 8430 12115 8434 12175
rect 8486 12155 8744 12175
rect 8430 12109 8486 12115
rect 8430 11921 8460 12109
rect 8515 12100 8715 12125
rect 8796 12115 8800 12175
rect 8744 12109 8800 12115
rect 8515 12080 8585 12100
rect 8490 12040 8585 12080
rect 8645 12080 8715 12100
rect 8645 12040 8740 12080
rect 8490 11990 8740 12040
rect 8490 11950 8585 11990
rect 8515 11930 8585 11950
rect 8645 11950 8740 11990
rect 8645 11930 8715 11950
rect 8430 11915 8486 11921
rect 8430 11855 8434 11915
rect 8515 11905 8715 11930
rect 8770 11921 8800 12109
rect 8744 11915 8800 11921
rect 8486 11855 8744 11875
rect 8796 11855 8800 11915
rect 8430 11845 8800 11855
rect 8830 12175 9200 12185
rect 8830 12115 8834 12175
rect 8886 12155 9144 12175
rect 8830 12109 8886 12115
rect 8830 11921 8860 12109
rect 8915 12100 9115 12125
rect 9196 12115 9200 12175
rect 9144 12109 9200 12115
rect 8915 12080 8985 12100
rect 8890 12040 8985 12080
rect 9045 12080 9115 12100
rect 9045 12040 9140 12080
rect 8890 11990 9140 12040
rect 8890 11950 8985 11990
rect 8915 11930 8985 11950
rect 9045 11950 9140 11990
rect 9045 11930 9115 11950
rect 8830 11915 8886 11921
rect 8830 11855 8834 11915
rect 8915 11905 9115 11930
rect 9170 11921 9200 12109
rect 9144 11915 9200 11921
rect 8886 11855 9144 11875
rect 9196 11855 9200 11915
rect 8830 11845 9200 11855
rect 9230 12175 9600 12185
rect 9230 12115 9234 12175
rect 9286 12155 9544 12175
rect 9230 12109 9286 12115
rect 9230 11921 9260 12109
rect 9315 12100 9515 12125
rect 9596 12115 9600 12175
rect 9544 12109 9600 12115
rect 9315 12080 9385 12100
rect 9290 12040 9385 12080
rect 9445 12080 9515 12100
rect 9445 12040 9540 12080
rect 9290 11990 9540 12040
rect 9290 11950 9385 11990
rect 9315 11930 9385 11950
rect 9445 11950 9540 11990
rect 9445 11930 9515 11950
rect 9230 11915 9286 11921
rect 9230 11855 9234 11915
rect 9315 11905 9515 11930
rect 9570 11921 9600 12109
rect 9544 11915 9600 11921
rect 9286 11855 9544 11875
rect 9596 11855 9600 11915
rect 9230 11845 9600 11855
rect 9630 12175 10000 12185
rect 9630 12115 9634 12175
rect 9686 12155 9944 12175
rect 9630 12109 9686 12115
rect 9630 11921 9660 12109
rect 9715 12100 9915 12125
rect 9996 12115 10000 12175
rect 9944 12109 10000 12115
rect 9715 12080 9785 12100
rect 9690 12040 9785 12080
rect 9845 12080 9915 12100
rect 9845 12040 9940 12080
rect 9690 11990 9940 12040
rect 9690 11950 9785 11990
rect 9715 11930 9785 11950
rect 9845 11950 9940 11990
rect 9845 11930 9915 11950
rect 9630 11915 9686 11921
rect 9630 11855 9634 11915
rect 9715 11905 9915 11930
rect 9970 11921 10000 12109
rect 9944 11915 10000 11921
rect 9686 11855 9944 11875
rect 9996 11855 10000 11915
rect 9630 11845 10000 11855
rect 10030 12175 10400 12185
rect 10030 12115 10034 12175
rect 10086 12155 10344 12175
rect 10030 12109 10086 12115
rect 10030 11921 10060 12109
rect 10115 12100 10315 12125
rect 10396 12115 10400 12175
rect 10344 12109 10400 12115
rect 10115 12080 10185 12100
rect 10090 12040 10185 12080
rect 10245 12080 10315 12100
rect 10245 12040 10340 12080
rect 10090 11990 10340 12040
rect 10090 11950 10185 11990
rect 10115 11930 10185 11950
rect 10245 11950 10340 11990
rect 10245 11930 10315 11950
rect 10030 11915 10086 11921
rect 10030 11855 10034 11915
rect 10115 11905 10315 11930
rect 10370 11921 10400 12109
rect 10344 11915 10400 11921
rect 10086 11855 10344 11875
rect 10396 11855 10400 11915
rect 10030 11845 10400 11855
rect 10430 12175 10800 12185
rect 10430 12115 10434 12175
rect 10486 12155 10744 12175
rect 10430 12109 10486 12115
rect 10430 11921 10460 12109
rect 10515 12100 10715 12125
rect 10796 12115 10800 12175
rect 10744 12109 10800 12115
rect 10515 12080 10585 12100
rect 10490 12040 10585 12080
rect 10645 12080 10715 12100
rect 10645 12040 10740 12080
rect 10490 11990 10740 12040
rect 10490 11950 10585 11990
rect 10515 11930 10585 11950
rect 10645 11950 10740 11990
rect 10645 11930 10715 11950
rect 10430 11915 10486 11921
rect 10430 11855 10434 11915
rect 10515 11905 10715 11930
rect 10770 11921 10800 12109
rect 10744 11915 10800 11921
rect 10486 11855 10744 11875
rect 10796 11855 10800 11915
rect 10430 11845 10800 11855
rect 10830 12175 11200 12185
rect 10830 12115 10834 12175
rect 10886 12155 11144 12175
rect 10830 12109 10886 12115
rect 10830 11921 10860 12109
rect 10915 12100 11115 12125
rect 11196 12115 11200 12175
rect 11144 12109 11200 12115
rect 10915 12080 10985 12100
rect 10890 12040 10985 12080
rect 11045 12080 11115 12100
rect 11045 12040 11140 12080
rect 10890 11990 11140 12040
rect 10890 11950 10985 11990
rect 10915 11930 10985 11950
rect 11045 11950 11140 11990
rect 11045 11930 11115 11950
rect 10830 11915 10886 11921
rect 10830 11855 10834 11915
rect 10915 11905 11115 11930
rect 11170 11921 11200 12109
rect 11144 11915 11200 11921
rect 10886 11855 11144 11875
rect 11196 11855 11200 11915
rect 10830 11845 11200 11855
rect 11230 12175 11600 12185
rect 11230 12115 11234 12175
rect 11286 12155 11544 12175
rect 11230 12109 11286 12115
rect 11230 11921 11260 12109
rect 11315 12100 11515 12125
rect 11596 12115 11600 12175
rect 11544 12109 11600 12115
rect 11315 12080 11385 12100
rect 11290 12040 11385 12080
rect 11445 12080 11515 12100
rect 11445 12040 11540 12080
rect 11290 11990 11540 12040
rect 11290 11950 11385 11990
rect 11315 11930 11385 11950
rect 11445 11950 11540 11990
rect 11445 11930 11515 11950
rect 11230 11915 11286 11921
rect 11230 11855 11234 11915
rect 11315 11905 11515 11930
rect 11570 11921 11600 12109
rect 11544 11915 11600 11921
rect 11286 11855 11544 11875
rect 11596 11855 11600 11915
rect 11230 11845 11600 11855
rect 11630 12175 12000 12185
rect 11630 12115 11634 12175
rect 11686 12155 11944 12175
rect 11630 12109 11686 12115
rect 11630 11921 11660 12109
rect 11715 12100 11915 12125
rect 11996 12115 12000 12175
rect 11944 12109 12000 12115
rect 11715 12080 11785 12100
rect 11690 12040 11785 12080
rect 11845 12080 11915 12100
rect 11845 12040 11940 12080
rect 11690 11990 11940 12040
rect 11690 11950 11785 11990
rect 11715 11930 11785 11950
rect 11845 11950 11940 11990
rect 11845 11930 11915 11950
rect 11630 11915 11686 11921
rect 11630 11855 11634 11915
rect 11715 11905 11915 11930
rect 11970 11921 12000 12109
rect 11944 11915 12000 11921
rect 11686 11855 11944 11875
rect 11996 11855 12000 11915
rect 11630 11845 12000 11855
rect 12030 12175 12400 12185
rect 12030 12115 12034 12175
rect 12086 12155 12344 12175
rect 12030 12109 12086 12115
rect 12030 11921 12060 12109
rect 12115 12100 12315 12125
rect 12396 12115 12400 12175
rect 12344 12109 12400 12115
rect 12115 12080 12185 12100
rect 12090 12040 12185 12080
rect 12245 12080 12315 12100
rect 12245 12040 12340 12080
rect 12090 11990 12340 12040
rect 12090 11950 12185 11990
rect 12115 11930 12185 11950
rect 12245 11950 12340 11990
rect 12245 11930 12315 11950
rect 12030 11915 12086 11921
rect 12030 11855 12034 11915
rect 12115 11905 12315 11930
rect 12370 11921 12400 12109
rect 12344 11915 12400 11921
rect 12086 11855 12344 11875
rect 12396 11855 12400 11915
rect 12030 11845 12400 11855
rect 12430 12175 12800 12185
rect 12430 12115 12434 12175
rect 12486 12155 12744 12175
rect 12430 12109 12486 12115
rect 12430 11921 12460 12109
rect 12515 12100 12715 12125
rect 12796 12115 12800 12175
rect 12744 12109 12800 12115
rect 12515 12080 12585 12100
rect 12490 12040 12585 12080
rect 12645 12080 12715 12100
rect 12645 12040 12740 12080
rect 12490 11990 12740 12040
rect 12490 11950 12585 11990
rect 12515 11930 12585 11950
rect 12645 11950 12740 11990
rect 12645 11930 12715 11950
rect 12430 11915 12486 11921
rect 12430 11855 12434 11915
rect 12515 11905 12715 11930
rect 12770 11921 12800 12109
rect 12744 11915 12800 11921
rect 12486 11855 12744 11875
rect 12796 11855 12800 11915
rect 12430 11845 12800 11855
rect 12830 12175 13200 12185
rect 12830 12115 12834 12175
rect 12886 12155 13144 12175
rect 12830 12109 12886 12115
rect 12830 11921 12860 12109
rect 12915 12100 13115 12125
rect 13196 12115 13200 12175
rect 13144 12109 13200 12115
rect 12915 12080 12985 12100
rect 12890 12040 12985 12080
rect 13045 12080 13115 12100
rect 13045 12040 13140 12080
rect 12890 11990 13140 12040
rect 12890 11950 12985 11990
rect 12915 11930 12985 11950
rect 13045 11950 13140 11990
rect 13045 11930 13115 11950
rect 12830 11915 12886 11921
rect 12830 11855 12834 11915
rect 12915 11905 13115 11930
rect 13170 11921 13200 12109
rect 13144 11915 13200 11921
rect 12886 11855 13144 11875
rect 13196 11855 13200 11915
rect 12830 11845 13200 11855
rect -370 11805 0 11815
rect -370 11745 -366 11805
rect -314 11785 -56 11805
rect -370 11739 -314 11745
rect -370 11551 -340 11739
rect -285 11730 -85 11755
rect -4 11745 0 11805
rect -56 11739 0 11745
rect -285 11710 -215 11730
rect -310 11670 -215 11710
rect -155 11710 -85 11730
rect -155 11670 -60 11710
rect -310 11620 -60 11670
rect -310 11580 -215 11620
rect -285 11560 -215 11580
rect -155 11580 -60 11620
rect -155 11560 -85 11580
rect -370 11545 -314 11551
rect -370 11485 -366 11545
rect -285 11535 -85 11560
rect -30 11551 0 11739
rect -56 11545 0 11551
rect -314 11485 -56 11505
rect -4 11485 0 11545
rect -370 11475 0 11485
rect 30 11805 400 11815
rect 30 11745 34 11805
rect 86 11785 344 11805
rect 30 11739 86 11745
rect 30 11551 60 11739
rect 115 11730 315 11755
rect 396 11745 400 11805
rect 344 11739 400 11745
rect 115 11710 185 11730
rect 90 11670 185 11710
rect 245 11710 315 11730
rect 245 11670 340 11710
rect 90 11620 340 11670
rect 90 11580 185 11620
rect 115 11560 185 11580
rect 245 11580 340 11620
rect 245 11560 315 11580
rect 30 11545 86 11551
rect 30 11485 34 11545
rect 115 11535 315 11560
rect 370 11551 400 11739
rect 344 11545 400 11551
rect 86 11485 344 11505
rect 396 11485 400 11545
rect 30 11475 400 11485
rect 430 11805 800 11815
rect 430 11745 434 11805
rect 486 11785 744 11805
rect 430 11739 486 11745
rect 430 11551 460 11739
rect 515 11730 715 11755
rect 796 11745 800 11805
rect 744 11739 800 11745
rect 515 11710 585 11730
rect 490 11670 585 11710
rect 645 11710 715 11730
rect 645 11670 740 11710
rect 490 11620 740 11670
rect 490 11580 585 11620
rect 515 11560 585 11580
rect 645 11580 740 11620
rect 645 11560 715 11580
rect 430 11545 486 11551
rect 430 11485 434 11545
rect 515 11535 715 11560
rect 770 11551 800 11739
rect 744 11545 800 11551
rect 486 11485 744 11505
rect 796 11485 800 11545
rect 430 11475 800 11485
rect 830 11805 1200 11815
rect 830 11745 834 11805
rect 886 11785 1144 11805
rect 830 11739 886 11745
rect 830 11551 860 11739
rect 915 11730 1115 11755
rect 1196 11745 1200 11805
rect 1144 11739 1200 11745
rect 915 11710 985 11730
rect 890 11670 985 11710
rect 1045 11710 1115 11730
rect 1045 11670 1140 11710
rect 890 11620 1140 11670
rect 890 11580 985 11620
rect 915 11560 985 11580
rect 1045 11580 1140 11620
rect 1045 11560 1115 11580
rect 830 11545 886 11551
rect 830 11485 834 11545
rect 915 11535 1115 11560
rect 1170 11551 1200 11739
rect 1144 11545 1200 11551
rect 886 11485 1144 11505
rect 1196 11485 1200 11545
rect 830 11475 1200 11485
rect 1230 11805 1600 11815
rect 1230 11745 1234 11805
rect 1286 11785 1544 11805
rect 1230 11739 1286 11745
rect 1230 11551 1260 11739
rect 1315 11730 1515 11755
rect 1596 11745 1600 11805
rect 1544 11739 1600 11745
rect 1315 11710 1385 11730
rect 1290 11670 1385 11710
rect 1445 11710 1515 11730
rect 1445 11670 1540 11710
rect 1290 11620 1540 11670
rect 1290 11580 1385 11620
rect 1315 11560 1385 11580
rect 1445 11580 1540 11620
rect 1445 11560 1515 11580
rect 1230 11545 1286 11551
rect 1230 11485 1234 11545
rect 1315 11535 1515 11560
rect 1570 11551 1600 11739
rect 1544 11545 1600 11551
rect 1286 11485 1544 11505
rect 1596 11485 1600 11545
rect 1230 11475 1600 11485
rect 1630 11805 2000 11815
rect 1630 11745 1634 11805
rect 1686 11785 1944 11805
rect 1630 11739 1686 11745
rect 1630 11551 1660 11739
rect 1715 11730 1915 11755
rect 1996 11745 2000 11805
rect 1944 11739 2000 11745
rect 1715 11710 1785 11730
rect 1690 11670 1785 11710
rect 1845 11710 1915 11730
rect 1845 11670 1940 11710
rect 1690 11620 1940 11670
rect 1690 11580 1785 11620
rect 1715 11560 1785 11580
rect 1845 11580 1940 11620
rect 1845 11560 1915 11580
rect 1630 11545 1686 11551
rect 1630 11485 1634 11545
rect 1715 11535 1915 11560
rect 1970 11551 2000 11739
rect 1944 11545 2000 11551
rect 1686 11485 1944 11505
rect 1996 11485 2000 11545
rect 1630 11475 2000 11485
rect 2030 11805 2400 11815
rect 2030 11745 2034 11805
rect 2086 11785 2344 11805
rect 2030 11739 2086 11745
rect 2030 11551 2060 11739
rect 2115 11730 2315 11755
rect 2396 11745 2400 11805
rect 2344 11739 2400 11745
rect 2115 11710 2185 11730
rect 2090 11670 2185 11710
rect 2245 11710 2315 11730
rect 2245 11670 2340 11710
rect 2090 11620 2340 11670
rect 2090 11580 2185 11620
rect 2115 11560 2185 11580
rect 2245 11580 2340 11620
rect 2245 11560 2315 11580
rect 2030 11545 2086 11551
rect 2030 11485 2034 11545
rect 2115 11535 2315 11560
rect 2370 11551 2400 11739
rect 2344 11545 2400 11551
rect 2086 11485 2344 11505
rect 2396 11485 2400 11545
rect 2030 11475 2400 11485
rect 2430 11805 2800 11815
rect 2430 11745 2434 11805
rect 2486 11785 2744 11805
rect 2430 11739 2486 11745
rect 2430 11551 2460 11739
rect 2515 11730 2715 11755
rect 2796 11745 2800 11805
rect 2744 11739 2800 11745
rect 2515 11710 2585 11730
rect 2490 11670 2585 11710
rect 2645 11710 2715 11730
rect 2645 11670 2740 11710
rect 2490 11620 2740 11670
rect 2490 11580 2585 11620
rect 2515 11560 2585 11580
rect 2645 11580 2740 11620
rect 2645 11560 2715 11580
rect 2430 11545 2486 11551
rect 2430 11485 2434 11545
rect 2515 11535 2715 11560
rect 2770 11551 2800 11739
rect 2744 11545 2800 11551
rect 2486 11485 2744 11505
rect 2796 11485 2800 11545
rect 2430 11475 2800 11485
rect 2830 11805 3200 11815
rect 2830 11745 2834 11805
rect 2886 11785 3144 11805
rect 2830 11739 2886 11745
rect 2830 11551 2860 11739
rect 2915 11730 3115 11755
rect 3196 11745 3200 11805
rect 3144 11739 3200 11745
rect 2915 11710 2985 11730
rect 2890 11670 2985 11710
rect 3045 11710 3115 11730
rect 3045 11670 3140 11710
rect 2890 11620 3140 11670
rect 2890 11580 2985 11620
rect 2915 11560 2985 11580
rect 3045 11580 3140 11620
rect 3045 11560 3115 11580
rect 2830 11545 2886 11551
rect 2830 11485 2834 11545
rect 2915 11535 3115 11560
rect 3170 11551 3200 11739
rect 3144 11545 3200 11551
rect 2886 11485 3144 11505
rect 3196 11485 3200 11545
rect 2830 11475 3200 11485
rect 3230 11805 3600 11815
rect 3230 11745 3234 11805
rect 3286 11785 3544 11805
rect 3230 11739 3286 11745
rect 3230 11551 3260 11739
rect 3315 11730 3515 11755
rect 3596 11745 3600 11805
rect 3544 11739 3600 11745
rect 3315 11710 3385 11730
rect 3290 11670 3385 11710
rect 3445 11710 3515 11730
rect 3445 11670 3540 11710
rect 3290 11620 3540 11670
rect 3290 11580 3385 11620
rect 3315 11560 3385 11580
rect 3445 11580 3540 11620
rect 3445 11560 3515 11580
rect 3230 11545 3286 11551
rect 3230 11485 3234 11545
rect 3315 11535 3515 11560
rect 3570 11551 3600 11739
rect 3544 11545 3600 11551
rect 3286 11485 3544 11505
rect 3596 11485 3600 11545
rect 3230 11475 3600 11485
rect 3630 11805 4000 11815
rect 3630 11745 3634 11805
rect 3686 11785 3944 11805
rect 3630 11739 3686 11745
rect 3630 11551 3660 11739
rect 3715 11730 3915 11755
rect 3996 11745 4000 11805
rect 3944 11739 4000 11745
rect 3715 11710 3785 11730
rect 3690 11670 3785 11710
rect 3845 11710 3915 11730
rect 3845 11670 3940 11710
rect 3690 11620 3940 11670
rect 3690 11580 3785 11620
rect 3715 11560 3785 11580
rect 3845 11580 3940 11620
rect 3845 11560 3915 11580
rect 3630 11545 3686 11551
rect 3630 11485 3634 11545
rect 3715 11535 3915 11560
rect 3970 11551 4000 11739
rect 3944 11545 4000 11551
rect 3686 11485 3944 11505
rect 3996 11485 4000 11545
rect 3630 11475 4000 11485
rect 4030 11805 4400 11815
rect 4030 11745 4034 11805
rect 4086 11785 4344 11805
rect 4030 11739 4086 11745
rect 4030 11551 4060 11739
rect 4115 11730 4315 11755
rect 4396 11745 4400 11805
rect 4344 11739 4400 11745
rect 4115 11710 4185 11730
rect 4090 11670 4185 11710
rect 4245 11710 4315 11730
rect 4245 11670 4340 11710
rect 4090 11620 4340 11670
rect 4090 11580 4185 11620
rect 4115 11560 4185 11580
rect 4245 11580 4340 11620
rect 4245 11560 4315 11580
rect 4030 11545 4086 11551
rect 4030 11485 4034 11545
rect 4115 11535 4315 11560
rect 4370 11551 4400 11739
rect 4344 11545 4400 11551
rect 4086 11485 4344 11505
rect 4396 11485 4400 11545
rect 4030 11475 4400 11485
rect 4430 11805 4800 11815
rect 4430 11745 4434 11805
rect 4486 11785 4744 11805
rect 4430 11739 4486 11745
rect 4430 11551 4460 11739
rect 4515 11730 4715 11755
rect 4796 11745 4800 11805
rect 4744 11739 4800 11745
rect 4515 11710 4585 11730
rect 4490 11670 4585 11710
rect 4645 11710 4715 11730
rect 4645 11670 4740 11710
rect 4490 11620 4740 11670
rect 4490 11580 4585 11620
rect 4515 11560 4585 11580
rect 4645 11580 4740 11620
rect 4645 11560 4715 11580
rect 4430 11545 4486 11551
rect 4430 11485 4434 11545
rect 4515 11535 4715 11560
rect 4770 11551 4800 11739
rect 4744 11545 4800 11551
rect 4486 11485 4744 11505
rect 4796 11485 4800 11545
rect 4430 11475 4800 11485
rect 4830 11805 5200 11815
rect 4830 11745 4834 11805
rect 4886 11785 5144 11805
rect 4830 11739 4886 11745
rect 4830 11551 4860 11739
rect 4915 11730 5115 11755
rect 5196 11745 5200 11805
rect 5144 11739 5200 11745
rect 4915 11710 4985 11730
rect 4890 11670 4985 11710
rect 5045 11710 5115 11730
rect 5045 11670 5140 11710
rect 4890 11620 5140 11670
rect 4890 11580 4985 11620
rect 4915 11560 4985 11580
rect 5045 11580 5140 11620
rect 5045 11560 5115 11580
rect 4830 11545 4886 11551
rect 4830 11485 4834 11545
rect 4915 11535 5115 11560
rect 5170 11551 5200 11739
rect 5144 11545 5200 11551
rect 4886 11485 5144 11505
rect 5196 11485 5200 11545
rect 4830 11475 5200 11485
rect 5230 11805 5600 11815
rect 5230 11745 5234 11805
rect 5286 11785 5544 11805
rect 5230 11739 5286 11745
rect 5230 11551 5260 11739
rect 5315 11730 5515 11755
rect 5596 11745 5600 11805
rect 5544 11739 5600 11745
rect 5315 11710 5385 11730
rect 5290 11670 5385 11710
rect 5445 11710 5515 11730
rect 5445 11670 5540 11710
rect 5290 11620 5540 11670
rect 5290 11580 5385 11620
rect 5315 11560 5385 11580
rect 5445 11580 5540 11620
rect 5445 11560 5515 11580
rect 5230 11545 5286 11551
rect 5230 11485 5234 11545
rect 5315 11535 5515 11560
rect 5570 11551 5600 11739
rect 5544 11545 5600 11551
rect 5286 11485 5544 11505
rect 5596 11485 5600 11545
rect 5230 11475 5600 11485
rect 5630 11805 6000 11815
rect 5630 11745 5634 11805
rect 5686 11785 5944 11805
rect 5630 11739 5686 11745
rect 5630 11551 5660 11739
rect 5715 11730 5915 11755
rect 5996 11745 6000 11805
rect 5944 11739 6000 11745
rect 5715 11710 5785 11730
rect 5690 11670 5785 11710
rect 5845 11710 5915 11730
rect 5845 11670 5940 11710
rect 5690 11620 5940 11670
rect 5690 11580 5785 11620
rect 5715 11560 5785 11580
rect 5845 11580 5940 11620
rect 5845 11560 5915 11580
rect 5630 11545 5686 11551
rect 5630 11485 5634 11545
rect 5715 11535 5915 11560
rect 5970 11551 6000 11739
rect 5944 11545 6000 11551
rect 5686 11485 5944 11505
rect 5996 11485 6000 11545
rect 5630 11475 6000 11485
rect 6030 11805 6400 11815
rect 6030 11745 6034 11805
rect 6086 11785 6344 11805
rect 6030 11739 6086 11745
rect 6030 11551 6060 11739
rect 6115 11730 6315 11755
rect 6396 11745 6400 11805
rect 6344 11739 6400 11745
rect 6115 11710 6185 11730
rect 6090 11670 6185 11710
rect 6245 11710 6315 11730
rect 6245 11670 6340 11710
rect 6090 11620 6340 11670
rect 6090 11580 6185 11620
rect 6115 11560 6185 11580
rect 6245 11580 6340 11620
rect 6245 11560 6315 11580
rect 6030 11545 6086 11551
rect 6030 11485 6034 11545
rect 6115 11535 6315 11560
rect 6370 11551 6400 11739
rect 6344 11545 6400 11551
rect 6086 11485 6344 11505
rect 6396 11485 6400 11545
rect 6030 11475 6400 11485
rect 6430 11805 6800 11815
rect 6430 11745 6434 11805
rect 6486 11785 6744 11805
rect 6430 11739 6486 11745
rect 6430 11551 6460 11739
rect 6515 11730 6715 11755
rect 6796 11745 6800 11805
rect 6744 11739 6800 11745
rect 6515 11710 6585 11730
rect 6490 11670 6585 11710
rect 6645 11710 6715 11730
rect 6645 11670 6740 11710
rect 6490 11620 6740 11670
rect 6490 11580 6585 11620
rect 6515 11560 6585 11580
rect 6645 11580 6740 11620
rect 6645 11560 6715 11580
rect 6430 11545 6486 11551
rect 6430 11485 6434 11545
rect 6515 11535 6715 11560
rect 6770 11551 6800 11739
rect 6744 11545 6800 11551
rect 6486 11485 6744 11505
rect 6796 11485 6800 11545
rect 6430 11475 6800 11485
rect 6830 11805 7200 11815
rect 6830 11745 6834 11805
rect 6886 11785 7144 11805
rect 6830 11739 6886 11745
rect 6830 11551 6860 11739
rect 6915 11730 7115 11755
rect 7196 11745 7200 11805
rect 7144 11739 7200 11745
rect 6915 11710 6985 11730
rect 6890 11670 6985 11710
rect 7045 11710 7115 11730
rect 7045 11670 7140 11710
rect 6890 11620 7140 11670
rect 6890 11580 6985 11620
rect 6915 11560 6985 11580
rect 7045 11580 7140 11620
rect 7045 11560 7115 11580
rect 6830 11545 6886 11551
rect 6830 11485 6834 11545
rect 6915 11535 7115 11560
rect 7170 11551 7200 11739
rect 7144 11545 7200 11551
rect 6886 11485 7144 11505
rect 7196 11485 7200 11545
rect 6830 11475 7200 11485
rect 7230 11805 7600 11815
rect 7230 11745 7234 11805
rect 7286 11785 7544 11805
rect 7230 11739 7286 11745
rect 7230 11551 7260 11739
rect 7315 11730 7515 11755
rect 7596 11745 7600 11805
rect 7544 11739 7600 11745
rect 7315 11710 7385 11730
rect 7290 11670 7385 11710
rect 7445 11710 7515 11730
rect 7445 11670 7540 11710
rect 7290 11620 7540 11670
rect 7290 11580 7385 11620
rect 7315 11560 7385 11580
rect 7445 11580 7540 11620
rect 7445 11560 7515 11580
rect 7230 11545 7286 11551
rect 7230 11485 7234 11545
rect 7315 11535 7515 11560
rect 7570 11551 7600 11739
rect 7544 11545 7600 11551
rect 7286 11485 7544 11505
rect 7596 11485 7600 11545
rect 7230 11475 7600 11485
rect 7630 11805 8000 11815
rect 7630 11745 7634 11805
rect 7686 11785 7944 11805
rect 7630 11739 7686 11745
rect 7630 11551 7660 11739
rect 7715 11730 7915 11755
rect 7996 11745 8000 11805
rect 7944 11739 8000 11745
rect 7715 11710 7785 11730
rect 7690 11670 7785 11710
rect 7845 11710 7915 11730
rect 7845 11670 7940 11710
rect 7690 11620 7940 11670
rect 7690 11580 7785 11620
rect 7715 11560 7785 11580
rect 7845 11580 7940 11620
rect 7845 11560 7915 11580
rect 7630 11545 7686 11551
rect 7630 11485 7634 11545
rect 7715 11535 7915 11560
rect 7970 11551 8000 11739
rect 7944 11545 8000 11551
rect 7686 11485 7944 11505
rect 7996 11485 8000 11545
rect 7630 11475 8000 11485
rect 8030 11805 8400 11815
rect 8030 11745 8034 11805
rect 8086 11785 8344 11805
rect 8030 11739 8086 11745
rect 8030 11551 8060 11739
rect 8115 11730 8315 11755
rect 8396 11745 8400 11805
rect 8344 11739 8400 11745
rect 8115 11710 8185 11730
rect 8090 11670 8185 11710
rect 8245 11710 8315 11730
rect 8245 11670 8340 11710
rect 8090 11620 8340 11670
rect 8090 11580 8185 11620
rect 8115 11560 8185 11580
rect 8245 11580 8340 11620
rect 8245 11560 8315 11580
rect 8030 11545 8086 11551
rect 8030 11485 8034 11545
rect 8115 11535 8315 11560
rect 8370 11551 8400 11739
rect 8344 11545 8400 11551
rect 8086 11485 8344 11505
rect 8396 11485 8400 11545
rect 8030 11475 8400 11485
rect 8430 11805 8800 11815
rect 8430 11745 8434 11805
rect 8486 11785 8744 11805
rect 8430 11739 8486 11745
rect 8430 11551 8460 11739
rect 8515 11730 8715 11755
rect 8796 11745 8800 11805
rect 8744 11739 8800 11745
rect 8515 11710 8585 11730
rect 8490 11670 8585 11710
rect 8645 11710 8715 11730
rect 8645 11670 8740 11710
rect 8490 11620 8740 11670
rect 8490 11580 8585 11620
rect 8515 11560 8585 11580
rect 8645 11580 8740 11620
rect 8645 11560 8715 11580
rect 8430 11545 8486 11551
rect 8430 11485 8434 11545
rect 8515 11535 8715 11560
rect 8770 11551 8800 11739
rect 8744 11545 8800 11551
rect 8486 11485 8744 11505
rect 8796 11485 8800 11545
rect 8430 11475 8800 11485
rect 8830 11805 9200 11815
rect 8830 11745 8834 11805
rect 8886 11785 9144 11805
rect 8830 11739 8886 11745
rect 8830 11551 8860 11739
rect 8915 11730 9115 11755
rect 9196 11745 9200 11805
rect 9144 11739 9200 11745
rect 8915 11710 8985 11730
rect 8890 11670 8985 11710
rect 9045 11710 9115 11730
rect 9045 11670 9140 11710
rect 8890 11620 9140 11670
rect 8890 11580 8985 11620
rect 8915 11560 8985 11580
rect 9045 11580 9140 11620
rect 9045 11560 9115 11580
rect 8830 11545 8886 11551
rect 8830 11485 8834 11545
rect 8915 11535 9115 11560
rect 9170 11551 9200 11739
rect 9144 11545 9200 11551
rect 8886 11485 9144 11505
rect 9196 11485 9200 11545
rect 8830 11475 9200 11485
rect 9230 11805 9600 11815
rect 9230 11745 9234 11805
rect 9286 11785 9544 11805
rect 9230 11739 9286 11745
rect 9230 11551 9260 11739
rect 9315 11730 9515 11755
rect 9596 11745 9600 11805
rect 9544 11739 9600 11745
rect 9315 11710 9385 11730
rect 9290 11670 9385 11710
rect 9445 11710 9515 11730
rect 9445 11670 9540 11710
rect 9290 11620 9540 11670
rect 9290 11580 9385 11620
rect 9315 11560 9385 11580
rect 9445 11580 9540 11620
rect 9445 11560 9515 11580
rect 9230 11545 9286 11551
rect 9230 11485 9234 11545
rect 9315 11535 9515 11560
rect 9570 11551 9600 11739
rect 9544 11545 9600 11551
rect 9286 11485 9544 11505
rect 9596 11485 9600 11545
rect 9230 11475 9600 11485
rect 9630 11805 10000 11815
rect 9630 11745 9634 11805
rect 9686 11785 9944 11805
rect 9630 11739 9686 11745
rect 9630 11551 9660 11739
rect 9715 11730 9915 11755
rect 9996 11745 10000 11805
rect 9944 11739 10000 11745
rect 9715 11710 9785 11730
rect 9690 11670 9785 11710
rect 9845 11710 9915 11730
rect 9845 11670 9940 11710
rect 9690 11620 9940 11670
rect 9690 11580 9785 11620
rect 9715 11560 9785 11580
rect 9845 11580 9940 11620
rect 9845 11560 9915 11580
rect 9630 11545 9686 11551
rect 9630 11485 9634 11545
rect 9715 11535 9915 11560
rect 9970 11551 10000 11739
rect 9944 11545 10000 11551
rect 9686 11485 9944 11505
rect 9996 11485 10000 11545
rect 9630 11475 10000 11485
rect 10030 11805 10400 11815
rect 10030 11745 10034 11805
rect 10086 11785 10344 11805
rect 10030 11739 10086 11745
rect 10030 11551 10060 11739
rect 10115 11730 10315 11755
rect 10396 11745 10400 11805
rect 10344 11739 10400 11745
rect 10115 11710 10185 11730
rect 10090 11670 10185 11710
rect 10245 11710 10315 11730
rect 10245 11670 10340 11710
rect 10090 11620 10340 11670
rect 10090 11580 10185 11620
rect 10115 11560 10185 11580
rect 10245 11580 10340 11620
rect 10245 11560 10315 11580
rect 10030 11545 10086 11551
rect 10030 11485 10034 11545
rect 10115 11535 10315 11560
rect 10370 11551 10400 11739
rect 10344 11545 10400 11551
rect 10086 11485 10344 11505
rect 10396 11485 10400 11545
rect 10030 11475 10400 11485
rect 10430 11805 10800 11815
rect 10430 11745 10434 11805
rect 10486 11785 10744 11805
rect 10430 11739 10486 11745
rect 10430 11551 10460 11739
rect 10515 11730 10715 11755
rect 10796 11745 10800 11805
rect 10744 11739 10800 11745
rect 10515 11710 10585 11730
rect 10490 11670 10585 11710
rect 10645 11710 10715 11730
rect 10645 11670 10740 11710
rect 10490 11620 10740 11670
rect 10490 11580 10585 11620
rect 10515 11560 10585 11580
rect 10645 11580 10740 11620
rect 10645 11560 10715 11580
rect 10430 11545 10486 11551
rect 10430 11485 10434 11545
rect 10515 11535 10715 11560
rect 10770 11551 10800 11739
rect 10744 11545 10800 11551
rect 10486 11485 10744 11505
rect 10796 11485 10800 11545
rect 10430 11475 10800 11485
rect 10830 11805 11200 11815
rect 10830 11745 10834 11805
rect 10886 11785 11144 11805
rect 10830 11739 10886 11745
rect 10830 11551 10860 11739
rect 10915 11730 11115 11755
rect 11196 11745 11200 11805
rect 11144 11739 11200 11745
rect 10915 11710 10985 11730
rect 10890 11670 10985 11710
rect 11045 11710 11115 11730
rect 11045 11670 11140 11710
rect 10890 11620 11140 11670
rect 10890 11580 10985 11620
rect 10915 11560 10985 11580
rect 11045 11580 11140 11620
rect 11045 11560 11115 11580
rect 10830 11545 10886 11551
rect 10830 11485 10834 11545
rect 10915 11535 11115 11560
rect 11170 11551 11200 11739
rect 11144 11545 11200 11551
rect 10886 11485 11144 11505
rect 11196 11485 11200 11545
rect 10830 11475 11200 11485
rect 11230 11805 11600 11815
rect 11230 11745 11234 11805
rect 11286 11785 11544 11805
rect 11230 11739 11286 11745
rect 11230 11551 11260 11739
rect 11315 11730 11515 11755
rect 11596 11745 11600 11805
rect 11544 11739 11600 11745
rect 11315 11710 11385 11730
rect 11290 11670 11385 11710
rect 11445 11710 11515 11730
rect 11445 11670 11540 11710
rect 11290 11620 11540 11670
rect 11290 11580 11385 11620
rect 11315 11560 11385 11580
rect 11445 11580 11540 11620
rect 11445 11560 11515 11580
rect 11230 11545 11286 11551
rect 11230 11485 11234 11545
rect 11315 11535 11515 11560
rect 11570 11551 11600 11739
rect 11544 11545 11600 11551
rect 11286 11485 11544 11505
rect 11596 11485 11600 11545
rect 11230 11475 11600 11485
rect 11630 11805 12000 11815
rect 11630 11745 11634 11805
rect 11686 11785 11944 11805
rect 11630 11739 11686 11745
rect 11630 11551 11660 11739
rect 11715 11730 11915 11755
rect 11996 11745 12000 11805
rect 11944 11739 12000 11745
rect 11715 11710 11785 11730
rect 11690 11670 11785 11710
rect 11845 11710 11915 11730
rect 11845 11670 11940 11710
rect 11690 11620 11940 11670
rect 11690 11580 11785 11620
rect 11715 11560 11785 11580
rect 11845 11580 11940 11620
rect 11845 11560 11915 11580
rect 11630 11545 11686 11551
rect 11630 11485 11634 11545
rect 11715 11535 11915 11560
rect 11970 11551 12000 11739
rect 11944 11545 12000 11551
rect 11686 11485 11944 11505
rect 11996 11485 12000 11545
rect 11630 11475 12000 11485
rect 12030 11805 12400 11815
rect 12030 11745 12034 11805
rect 12086 11785 12344 11805
rect 12030 11739 12086 11745
rect 12030 11551 12060 11739
rect 12115 11730 12315 11755
rect 12396 11745 12400 11805
rect 12344 11739 12400 11745
rect 12115 11710 12185 11730
rect 12090 11670 12185 11710
rect 12245 11710 12315 11730
rect 12245 11670 12340 11710
rect 12090 11620 12340 11670
rect 12090 11580 12185 11620
rect 12115 11560 12185 11580
rect 12245 11580 12340 11620
rect 12245 11560 12315 11580
rect 12030 11545 12086 11551
rect 12030 11485 12034 11545
rect 12115 11535 12315 11560
rect 12370 11551 12400 11739
rect 12344 11545 12400 11551
rect 12086 11485 12344 11505
rect 12396 11485 12400 11545
rect 12030 11475 12400 11485
rect 12430 11805 12800 11815
rect 12430 11745 12434 11805
rect 12486 11785 12744 11805
rect 12430 11739 12486 11745
rect 12430 11551 12460 11739
rect 12515 11730 12715 11755
rect 12796 11745 12800 11805
rect 12744 11739 12800 11745
rect 12515 11710 12585 11730
rect 12490 11670 12585 11710
rect 12645 11710 12715 11730
rect 12645 11670 12740 11710
rect 12490 11620 12740 11670
rect 12490 11580 12585 11620
rect 12515 11560 12585 11580
rect 12645 11580 12740 11620
rect 12645 11560 12715 11580
rect 12430 11545 12486 11551
rect 12430 11485 12434 11545
rect 12515 11535 12715 11560
rect 12770 11551 12800 11739
rect 12744 11545 12800 11551
rect 12486 11485 12744 11505
rect 12796 11485 12800 11545
rect 12430 11475 12800 11485
rect 12830 11805 13200 11815
rect 12830 11745 12834 11805
rect 12886 11785 13144 11805
rect 12830 11739 12886 11745
rect 12830 11551 12860 11739
rect 12915 11730 13115 11755
rect 13196 11745 13200 11805
rect 13144 11739 13200 11745
rect 12915 11710 12985 11730
rect 12890 11670 12985 11710
rect 13045 11710 13115 11730
rect 13045 11670 13140 11710
rect 12890 11620 13140 11670
rect 12890 11580 12985 11620
rect 12915 11560 12985 11580
rect 13045 11580 13140 11620
rect 13045 11560 13115 11580
rect 12830 11545 12886 11551
rect 12830 11485 12834 11545
rect 12915 11535 13115 11560
rect 13170 11551 13200 11739
rect 13144 11545 13200 11551
rect 12886 11485 13144 11505
rect 13196 11485 13200 11545
rect 12830 11475 13200 11485
rect -370 11435 0 11445
rect -370 11375 -366 11435
rect -314 11415 -56 11435
rect -370 11369 -314 11375
rect -370 11181 -340 11369
rect -285 11360 -85 11385
rect -4 11375 0 11435
rect -56 11369 0 11375
rect -285 11340 -215 11360
rect -310 11300 -215 11340
rect -155 11340 -85 11360
rect -155 11300 -60 11340
rect -310 11250 -60 11300
rect -310 11210 -215 11250
rect -285 11190 -215 11210
rect -155 11210 -60 11250
rect -155 11190 -85 11210
rect -370 11175 -314 11181
rect -370 11115 -366 11175
rect -285 11165 -85 11190
rect -30 11181 0 11369
rect -56 11175 0 11181
rect -314 11115 -56 11135
rect -4 11115 0 11175
rect -370 11105 0 11115
rect 30 11435 400 11445
rect 30 11375 34 11435
rect 86 11415 344 11435
rect 30 11369 86 11375
rect 30 11181 60 11369
rect 115 11360 315 11385
rect 396 11375 400 11435
rect 344 11369 400 11375
rect 115 11340 185 11360
rect 90 11300 185 11340
rect 245 11340 315 11360
rect 245 11300 340 11340
rect 90 11250 340 11300
rect 90 11210 185 11250
rect 115 11190 185 11210
rect 245 11210 340 11250
rect 245 11190 315 11210
rect 30 11175 86 11181
rect 30 11115 34 11175
rect 115 11165 315 11190
rect 370 11181 400 11369
rect 344 11175 400 11181
rect 86 11115 344 11135
rect 396 11115 400 11175
rect 30 11105 400 11115
rect 430 11435 800 11445
rect 430 11375 434 11435
rect 486 11415 744 11435
rect 430 11369 486 11375
rect 430 11181 460 11369
rect 515 11360 715 11385
rect 796 11375 800 11435
rect 744 11369 800 11375
rect 515 11340 585 11360
rect 490 11300 585 11340
rect 645 11340 715 11360
rect 645 11300 740 11340
rect 490 11250 740 11300
rect 490 11210 585 11250
rect 515 11190 585 11210
rect 645 11210 740 11250
rect 645 11190 715 11210
rect 430 11175 486 11181
rect 430 11115 434 11175
rect 515 11165 715 11190
rect 770 11181 800 11369
rect 744 11175 800 11181
rect 486 11115 744 11135
rect 796 11115 800 11175
rect 430 11105 800 11115
rect 830 11435 1200 11445
rect 830 11375 834 11435
rect 886 11415 1144 11435
rect 830 11369 886 11375
rect 830 11181 860 11369
rect 915 11360 1115 11385
rect 1196 11375 1200 11435
rect 1144 11369 1200 11375
rect 915 11340 985 11360
rect 890 11300 985 11340
rect 1045 11340 1115 11360
rect 1045 11300 1140 11340
rect 890 11250 1140 11300
rect 890 11210 985 11250
rect 915 11190 985 11210
rect 1045 11210 1140 11250
rect 1045 11190 1115 11210
rect 830 11175 886 11181
rect 830 11115 834 11175
rect 915 11165 1115 11190
rect 1170 11181 1200 11369
rect 1144 11175 1200 11181
rect 886 11115 1144 11135
rect 1196 11115 1200 11175
rect 830 11105 1200 11115
rect 1230 11435 1600 11445
rect 1230 11375 1234 11435
rect 1286 11415 1544 11435
rect 1230 11369 1286 11375
rect 1230 11181 1260 11369
rect 1315 11360 1515 11385
rect 1596 11375 1600 11435
rect 1544 11369 1600 11375
rect 1315 11340 1385 11360
rect 1290 11300 1385 11340
rect 1445 11340 1515 11360
rect 1445 11300 1540 11340
rect 1290 11250 1540 11300
rect 1290 11210 1385 11250
rect 1315 11190 1385 11210
rect 1445 11210 1540 11250
rect 1445 11190 1515 11210
rect 1230 11175 1286 11181
rect 1230 11115 1234 11175
rect 1315 11165 1515 11190
rect 1570 11181 1600 11369
rect 1544 11175 1600 11181
rect 1286 11115 1544 11135
rect 1596 11115 1600 11175
rect 1230 11105 1600 11115
rect 1630 11435 2000 11445
rect 1630 11375 1634 11435
rect 1686 11415 1944 11435
rect 1630 11369 1686 11375
rect 1630 11181 1660 11369
rect 1715 11360 1915 11385
rect 1996 11375 2000 11435
rect 1944 11369 2000 11375
rect 1715 11340 1785 11360
rect 1690 11300 1785 11340
rect 1845 11340 1915 11360
rect 1845 11300 1940 11340
rect 1690 11250 1940 11300
rect 1690 11210 1785 11250
rect 1715 11190 1785 11210
rect 1845 11210 1940 11250
rect 1845 11190 1915 11210
rect 1630 11175 1686 11181
rect 1630 11115 1634 11175
rect 1715 11165 1915 11190
rect 1970 11181 2000 11369
rect 1944 11175 2000 11181
rect 1686 11115 1944 11135
rect 1996 11115 2000 11175
rect 1630 11105 2000 11115
rect 2030 11435 2400 11445
rect 2030 11375 2034 11435
rect 2086 11415 2344 11435
rect 2030 11369 2086 11375
rect 2030 11181 2060 11369
rect 2115 11360 2315 11385
rect 2396 11375 2400 11435
rect 2344 11369 2400 11375
rect 2115 11340 2185 11360
rect 2090 11300 2185 11340
rect 2245 11340 2315 11360
rect 2245 11300 2340 11340
rect 2090 11250 2340 11300
rect 2090 11210 2185 11250
rect 2115 11190 2185 11210
rect 2245 11210 2340 11250
rect 2245 11190 2315 11210
rect 2030 11175 2086 11181
rect 2030 11115 2034 11175
rect 2115 11165 2315 11190
rect 2370 11181 2400 11369
rect 2344 11175 2400 11181
rect 2086 11115 2344 11135
rect 2396 11115 2400 11175
rect 2030 11105 2400 11115
rect 2430 11435 2800 11445
rect 2430 11375 2434 11435
rect 2486 11415 2744 11435
rect 2430 11369 2486 11375
rect 2430 11181 2460 11369
rect 2515 11360 2715 11385
rect 2796 11375 2800 11435
rect 2744 11369 2800 11375
rect 2515 11340 2585 11360
rect 2490 11300 2585 11340
rect 2645 11340 2715 11360
rect 2645 11300 2740 11340
rect 2490 11250 2740 11300
rect 2490 11210 2585 11250
rect 2515 11190 2585 11210
rect 2645 11210 2740 11250
rect 2645 11190 2715 11210
rect 2430 11175 2486 11181
rect 2430 11115 2434 11175
rect 2515 11165 2715 11190
rect 2770 11181 2800 11369
rect 2744 11175 2800 11181
rect 2486 11115 2744 11135
rect 2796 11115 2800 11175
rect 2430 11105 2800 11115
rect 2830 11435 3200 11445
rect 2830 11375 2834 11435
rect 2886 11415 3144 11435
rect 2830 11369 2886 11375
rect 2830 11181 2860 11369
rect 2915 11360 3115 11385
rect 3196 11375 3200 11435
rect 3144 11369 3200 11375
rect 2915 11340 2985 11360
rect 2890 11300 2985 11340
rect 3045 11340 3115 11360
rect 3045 11300 3140 11340
rect 2890 11250 3140 11300
rect 2890 11210 2985 11250
rect 2915 11190 2985 11210
rect 3045 11210 3140 11250
rect 3045 11190 3115 11210
rect 2830 11175 2886 11181
rect 2830 11115 2834 11175
rect 2915 11165 3115 11190
rect 3170 11181 3200 11369
rect 3144 11175 3200 11181
rect 2886 11115 3144 11135
rect 3196 11115 3200 11175
rect 2830 11105 3200 11115
rect 3230 11435 3600 11445
rect 3230 11375 3234 11435
rect 3286 11415 3544 11435
rect 3230 11369 3286 11375
rect 3230 11181 3260 11369
rect 3315 11360 3515 11385
rect 3596 11375 3600 11435
rect 3544 11369 3600 11375
rect 3315 11340 3385 11360
rect 3290 11300 3385 11340
rect 3445 11340 3515 11360
rect 3445 11300 3540 11340
rect 3290 11250 3540 11300
rect 3290 11210 3385 11250
rect 3315 11190 3385 11210
rect 3445 11210 3540 11250
rect 3445 11190 3515 11210
rect 3230 11175 3286 11181
rect 3230 11115 3234 11175
rect 3315 11165 3515 11190
rect 3570 11181 3600 11369
rect 3544 11175 3600 11181
rect 3286 11115 3544 11135
rect 3596 11115 3600 11175
rect 3230 11105 3600 11115
rect 3630 11435 4000 11445
rect 3630 11375 3634 11435
rect 3686 11415 3944 11435
rect 3630 11369 3686 11375
rect 3630 11181 3660 11369
rect 3715 11360 3915 11385
rect 3996 11375 4000 11435
rect 3944 11369 4000 11375
rect 3715 11340 3785 11360
rect 3690 11300 3785 11340
rect 3845 11340 3915 11360
rect 3845 11300 3940 11340
rect 3690 11250 3940 11300
rect 3690 11210 3785 11250
rect 3715 11190 3785 11210
rect 3845 11210 3940 11250
rect 3845 11190 3915 11210
rect 3630 11175 3686 11181
rect 3630 11115 3634 11175
rect 3715 11165 3915 11190
rect 3970 11181 4000 11369
rect 3944 11175 4000 11181
rect 3686 11115 3944 11135
rect 3996 11115 4000 11175
rect 3630 11105 4000 11115
rect 4030 11435 4400 11445
rect 4030 11375 4034 11435
rect 4086 11415 4344 11435
rect 4030 11369 4086 11375
rect 4030 11181 4060 11369
rect 4115 11360 4315 11385
rect 4396 11375 4400 11435
rect 4344 11369 4400 11375
rect 4115 11340 4185 11360
rect 4090 11300 4185 11340
rect 4245 11340 4315 11360
rect 4245 11300 4340 11340
rect 4090 11250 4340 11300
rect 4090 11210 4185 11250
rect 4115 11190 4185 11210
rect 4245 11210 4340 11250
rect 4245 11190 4315 11210
rect 4030 11175 4086 11181
rect 4030 11115 4034 11175
rect 4115 11165 4315 11190
rect 4370 11181 4400 11369
rect 4344 11175 4400 11181
rect 4086 11115 4344 11135
rect 4396 11115 4400 11175
rect 4030 11105 4400 11115
rect 4430 11435 4800 11445
rect 4430 11375 4434 11435
rect 4486 11415 4744 11435
rect 4430 11369 4486 11375
rect 4430 11181 4460 11369
rect 4515 11360 4715 11385
rect 4796 11375 4800 11435
rect 4744 11369 4800 11375
rect 4515 11340 4585 11360
rect 4490 11300 4585 11340
rect 4645 11340 4715 11360
rect 4645 11300 4740 11340
rect 4490 11250 4740 11300
rect 4490 11210 4585 11250
rect 4515 11190 4585 11210
rect 4645 11210 4740 11250
rect 4645 11190 4715 11210
rect 4430 11175 4486 11181
rect 4430 11115 4434 11175
rect 4515 11165 4715 11190
rect 4770 11181 4800 11369
rect 4744 11175 4800 11181
rect 4486 11115 4744 11135
rect 4796 11115 4800 11175
rect 4430 11105 4800 11115
rect 4830 11435 5200 11445
rect 4830 11375 4834 11435
rect 4886 11415 5144 11435
rect 4830 11369 4886 11375
rect 4830 11181 4860 11369
rect 4915 11360 5115 11385
rect 5196 11375 5200 11435
rect 5144 11369 5200 11375
rect 4915 11340 4985 11360
rect 4890 11300 4985 11340
rect 5045 11340 5115 11360
rect 5045 11300 5140 11340
rect 4890 11250 5140 11300
rect 4890 11210 4985 11250
rect 4915 11190 4985 11210
rect 5045 11210 5140 11250
rect 5045 11190 5115 11210
rect 4830 11175 4886 11181
rect 4830 11115 4834 11175
rect 4915 11165 5115 11190
rect 5170 11181 5200 11369
rect 5144 11175 5200 11181
rect 4886 11115 5144 11135
rect 5196 11115 5200 11175
rect 4830 11105 5200 11115
rect 5230 11435 5600 11445
rect 5230 11375 5234 11435
rect 5286 11415 5544 11435
rect 5230 11369 5286 11375
rect 5230 11181 5260 11369
rect 5315 11360 5515 11385
rect 5596 11375 5600 11435
rect 5544 11369 5600 11375
rect 5315 11340 5385 11360
rect 5290 11300 5385 11340
rect 5445 11340 5515 11360
rect 5445 11300 5540 11340
rect 5290 11250 5540 11300
rect 5290 11210 5385 11250
rect 5315 11190 5385 11210
rect 5445 11210 5540 11250
rect 5445 11190 5515 11210
rect 5230 11175 5286 11181
rect 5230 11115 5234 11175
rect 5315 11165 5515 11190
rect 5570 11181 5600 11369
rect 5544 11175 5600 11181
rect 5286 11115 5544 11135
rect 5596 11115 5600 11175
rect 5230 11105 5600 11115
rect 5630 11435 6000 11445
rect 5630 11375 5634 11435
rect 5686 11415 5944 11435
rect 5630 11369 5686 11375
rect 5630 11181 5660 11369
rect 5715 11360 5915 11385
rect 5996 11375 6000 11435
rect 5944 11369 6000 11375
rect 5715 11340 5785 11360
rect 5690 11300 5785 11340
rect 5845 11340 5915 11360
rect 5845 11300 5940 11340
rect 5690 11250 5940 11300
rect 5690 11210 5785 11250
rect 5715 11190 5785 11210
rect 5845 11210 5940 11250
rect 5845 11190 5915 11210
rect 5630 11175 5686 11181
rect 5630 11115 5634 11175
rect 5715 11165 5915 11190
rect 5970 11181 6000 11369
rect 5944 11175 6000 11181
rect 5686 11115 5944 11135
rect 5996 11115 6000 11175
rect 5630 11105 6000 11115
rect 6030 11435 6400 11445
rect 6030 11375 6034 11435
rect 6086 11415 6344 11435
rect 6030 11369 6086 11375
rect 6030 11181 6060 11369
rect 6115 11360 6315 11385
rect 6396 11375 6400 11435
rect 6344 11369 6400 11375
rect 6115 11340 6185 11360
rect 6090 11300 6185 11340
rect 6245 11340 6315 11360
rect 6245 11300 6340 11340
rect 6090 11250 6340 11300
rect 6090 11210 6185 11250
rect 6115 11190 6185 11210
rect 6245 11210 6340 11250
rect 6245 11190 6315 11210
rect 6030 11175 6086 11181
rect 6030 11115 6034 11175
rect 6115 11165 6315 11190
rect 6370 11181 6400 11369
rect 6344 11175 6400 11181
rect 6086 11115 6344 11135
rect 6396 11115 6400 11175
rect 6030 11105 6400 11115
rect 6430 11435 6800 11445
rect 6430 11375 6434 11435
rect 6486 11415 6744 11435
rect 6430 11369 6486 11375
rect 6430 11181 6460 11369
rect 6515 11360 6715 11385
rect 6796 11375 6800 11435
rect 6744 11369 6800 11375
rect 6515 11340 6585 11360
rect 6490 11300 6585 11340
rect 6645 11340 6715 11360
rect 6645 11300 6740 11340
rect 6490 11250 6740 11300
rect 6490 11210 6585 11250
rect 6515 11190 6585 11210
rect 6645 11210 6740 11250
rect 6645 11190 6715 11210
rect 6430 11175 6486 11181
rect 6430 11115 6434 11175
rect 6515 11165 6715 11190
rect 6770 11181 6800 11369
rect 6744 11175 6800 11181
rect 6486 11115 6744 11135
rect 6796 11115 6800 11175
rect 6430 11105 6800 11115
rect 6830 11435 7200 11445
rect 6830 11375 6834 11435
rect 6886 11415 7144 11435
rect 6830 11369 6886 11375
rect 6830 11181 6860 11369
rect 6915 11360 7115 11385
rect 7196 11375 7200 11435
rect 7144 11369 7200 11375
rect 6915 11340 6985 11360
rect 6890 11300 6985 11340
rect 7045 11340 7115 11360
rect 7045 11300 7140 11340
rect 6890 11250 7140 11300
rect 6890 11210 6985 11250
rect 6915 11190 6985 11210
rect 7045 11210 7140 11250
rect 7045 11190 7115 11210
rect 6830 11175 6886 11181
rect 6830 11115 6834 11175
rect 6915 11165 7115 11190
rect 7170 11181 7200 11369
rect 7144 11175 7200 11181
rect 6886 11115 7144 11135
rect 7196 11115 7200 11175
rect 6830 11105 7200 11115
rect 7230 11435 7600 11445
rect 7230 11375 7234 11435
rect 7286 11415 7544 11435
rect 7230 11369 7286 11375
rect 7230 11181 7260 11369
rect 7315 11360 7515 11385
rect 7596 11375 7600 11435
rect 7544 11369 7600 11375
rect 7315 11340 7385 11360
rect 7290 11300 7385 11340
rect 7445 11340 7515 11360
rect 7445 11300 7540 11340
rect 7290 11250 7540 11300
rect 7290 11210 7385 11250
rect 7315 11190 7385 11210
rect 7445 11210 7540 11250
rect 7445 11190 7515 11210
rect 7230 11175 7286 11181
rect 7230 11115 7234 11175
rect 7315 11165 7515 11190
rect 7570 11181 7600 11369
rect 7544 11175 7600 11181
rect 7286 11115 7544 11135
rect 7596 11115 7600 11175
rect 7230 11105 7600 11115
rect 7630 11435 8000 11445
rect 7630 11375 7634 11435
rect 7686 11415 7944 11435
rect 7630 11369 7686 11375
rect 7630 11181 7660 11369
rect 7715 11360 7915 11385
rect 7996 11375 8000 11435
rect 7944 11369 8000 11375
rect 7715 11340 7785 11360
rect 7690 11300 7785 11340
rect 7845 11340 7915 11360
rect 7845 11300 7940 11340
rect 7690 11250 7940 11300
rect 7690 11210 7785 11250
rect 7715 11190 7785 11210
rect 7845 11210 7940 11250
rect 7845 11190 7915 11210
rect 7630 11175 7686 11181
rect 7630 11115 7634 11175
rect 7715 11165 7915 11190
rect 7970 11181 8000 11369
rect 7944 11175 8000 11181
rect 7686 11115 7944 11135
rect 7996 11115 8000 11175
rect 7630 11105 8000 11115
rect 8030 11435 8400 11445
rect 8030 11375 8034 11435
rect 8086 11415 8344 11435
rect 8030 11369 8086 11375
rect 8030 11181 8060 11369
rect 8115 11360 8315 11385
rect 8396 11375 8400 11435
rect 8344 11369 8400 11375
rect 8115 11340 8185 11360
rect 8090 11300 8185 11340
rect 8245 11340 8315 11360
rect 8245 11300 8340 11340
rect 8090 11250 8340 11300
rect 8090 11210 8185 11250
rect 8115 11190 8185 11210
rect 8245 11210 8340 11250
rect 8245 11190 8315 11210
rect 8030 11175 8086 11181
rect 8030 11115 8034 11175
rect 8115 11165 8315 11190
rect 8370 11181 8400 11369
rect 8344 11175 8400 11181
rect 8086 11115 8344 11135
rect 8396 11115 8400 11175
rect 8030 11105 8400 11115
rect 8430 11435 8800 11445
rect 8430 11375 8434 11435
rect 8486 11415 8744 11435
rect 8430 11369 8486 11375
rect 8430 11181 8460 11369
rect 8515 11360 8715 11385
rect 8796 11375 8800 11435
rect 8744 11369 8800 11375
rect 8515 11340 8585 11360
rect 8490 11300 8585 11340
rect 8645 11340 8715 11360
rect 8645 11300 8740 11340
rect 8490 11250 8740 11300
rect 8490 11210 8585 11250
rect 8515 11190 8585 11210
rect 8645 11210 8740 11250
rect 8645 11190 8715 11210
rect 8430 11175 8486 11181
rect 8430 11115 8434 11175
rect 8515 11165 8715 11190
rect 8770 11181 8800 11369
rect 8744 11175 8800 11181
rect 8486 11115 8744 11135
rect 8796 11115 8800 11175
rect 8430 11105 8800 11115
rect 8830 11435 9200 11445
rect 8830 11375 8834 11435
rect 8886 11415 9144 11435
rect 8830 11369 8886 11375
rect 8830 11181 8860 11369
rect 8915 11360 9115 11385
rect 9196 11375 9200 11435
rect 9144 11369 9200 11375
rect 8915 11340 8985 11360
rect 8890 11300 8985 11340
rect 9045 11340 9115 11360
rect 9045 11300 9140 11340
rect 8890 11250 9140 11300
rect 8890 11210 8985 11250
rect 8915 11190 8985 11210
rect 9045 11210 9140 11250
rect 9045 11190 9115 11210
rect 8830 11175 8886 11181
rect 8830 11115 8834 11175
rect 8915 11165 9115 11190
rect 9170 11181 9200 11369
rect 9144 11175 9200 11181
rect 8886 11115 9144 11135
rect 9196 11115 9200 11175
rect 8830 11105 9200 11115
rect 9230 11435 9600 11445
rect 9230 11375 9234 11435
rect 9286 11415 9544 11435
rect 9230 11369 9286 11375
rect 9230 11181 9260 11369
rect 9315 11360 9515 11385
rect 9596 11375 9600 11435
rect 9544 11369 9600 11375
rect 9315 11340 9385 11360
rect 9290 11300 9385 11340
rect 9445 11340 9515 11360
rect 9445 11300 9540 11340
rect 9290 11250 9540 11300
rect 9290 11210 9385 11250
rect 9315 11190 9385 11210
rect 9445 11210 9540 11250
rect 9445 11190 9515 11210
rect 9230 11175 9286 11181
rect 9230 11115 9234 11175
rect 9315 11165 9515 11190
rect 9570 11181 9600 11369
rect 9544 11175 9600 11181
rect 9286 11115 9544 11135
rect 9596 11115 9600 11175
rect 9230 11105 9600 11115
rect 9630 11435 10000 11445
rect 9630 11375 9634 11435
rect 9686 11415 9944 11435
rect 9630 11369 9686 11375
rect 9630 11181 9660 11369
rect 9715 11360 9915 11385
rect 9996 11375 10000 11435
rect 9944 11369 10000 11375
rect 9715 11340 9785 11360
rect 9690 11300 9785 11340
rect 9845 11340 9915 11360
rect 9845 11300 9940 11340
rect 9690 11250 9940 11300
rect 9690 11210 9785 11250
rect 9715 11190 9785 11210
rect 9845 11210 9940 11250
rect 9845 11190 9915 11210
rect 9630 11175 9686 11181
rect 9630 11115 9634 11175
rect 9715 11165 9915 11190
rect 9970 11181 10000 11369
rect 9944 11175 10000 11181
rect 9686 11115 9944 11135
rect 9996 11115 10000 11175
rect 9630 11105 10000 11115
rect 10030 11435 10400 11445
rect 10030 11375 10034 11435
rect 10086 11415 10344 11435
rect 10030 11369 10086 11375
rect 10030 11181 10060 11369
rect 10115 11360 10315 11385
rect 10396 11375 10400 11435
rect 10344 11369 10400 11375
rect 10115 11340 10185 11360
rect 10090 11300 10185 11340
rect 10245 11340 10315 11360
rect 10245 11300 10340 11340
rect 10090 11250 10340 11300
rect 10090 11210 10185 11250
rect 10115 11190 10185 11210
rect 10245 11210 10340 11250
rect 10245 11190 10315 11210
rect 10030 11175 10086 11181
rect 10030 11115 10034 11175
rect 10115 11165 10315 11190
rect 10370 11181 10400 11369
rect 10344 11175 10400 11181
rect 10086 11115 10344 11135
rect 10396 11115 10400 11175
rect 10030 11105 10400 11115
rect 10430 11435 10800 11445
rect 10430 11375 10434 11435
rect 10486 11415 10744 11435
rect 10430 11369 10486 11375
rect 10430 11181 10460 11369
rect 10515 11360 10715 11385
rect 10796 11375 10800 11435
rect 10744 11369 10800 11375
rect 10515 11340 10585 11360
rect 10490 11300 10585 11340
rect 10645 11340 10715 11360
rect 10645 11300 10740 11340
rect 10490 11250 10740 11300
rect 10490 11210 10585 11250
rect 10515 11190 10585 11210
rect 10645 11210 10740 11250
rect 10645 11190 10715 11210
rect 10430 11175 10486 11181
rect 10430 11115 10434 11175
rect 10515 11165 10715 11190
rect 10770 11181 10800 11369
rect 10744 11175 10800 11181
rect 10486 11115 10744 11135
rect 10796 11115 10800 11175
rect 10430 11105 10800 11115
rect 10830 11435 11200 11445
rect 10830 11375 10834 11435
rect 10886 11415 11144 11435
rect 10830 11369 10886 11375
rect 10830 11181 10860 11369
rect 10915 11360 11115 11385
rect 11196 11375 11200 11435
rect 11144 11369 11200 11375
rect 10915 11340 10985 11360
rect 10890 11300 10985 11340
rect 11045 11340 11115 11360
rect 11045 11300 11140 11340
rect 10890 11250 11140 11300
rect 10890 11210 10985 11250
rect 10915 11190 10985 11210
rect 11045 11210 11140 11250
rect 11045 11190 11115 11210
rect 10830 11175 10886 11181
rect 10830 11115 10834 11175
rect 10915 11165 11115 11190
rect 11170 11181 11200 11369
rect 11144 11175 11200 11181
rect 10886 11115 11144 11135
rect 11196 11115 11200 11175
rect 10830 11105 11200 11115
rect 11230 11435 11600 11445
rect 11230 11375 11234 11435
rect 11286 11415 11544 11435
rect 11230 11369 11286 11375
rect 11230 11181 11260 11369
rect 11315 11360 11515 11385
rect 11596 11375 11600 11435
rect 11544 11369 11600 11375
rect 11315 11340 11385 11360
rect 11290 11300 11385 11340
rect 11445 11340 11515 11360
rect 11445 11300 11540 11340
rect 11290 11250 11540 11300
rect 11290 11210 11385 11250
rect 11315 11190 11385 11210
rect 11445 11210 11540 11250
rect 11445 11190 11515 11210
rect 11230 11175 11286 11181
rect 11230 11115 11234 11175
rect 11315 11165 11515 11190
rect 11570 11181 11600 11369
rect 11544 11175 11600 11181
rect 11286 11115 11544 11135
rect 11596 11115 11600 11175
rect 11230 11105 11600 11115
rect 11630 11435 12000 11445
rect 11630 11375 11634 11435
rect 11686 11415 11944 11435
rect 11630 11369 11686 11375
rect 11630 11181 11660 11369
rect 11715 11360 11915 11385
rect 11996 11375 12000 11435
rect 11944 11369 12000 11375
rect 11715 11340 11785 11360
rect 11690 11300 11785 11340
rect 11845 11340 11915 11360
rect 11845 11300 11940 11340
rect 11690 11250 11940 11300
rect 11690 11210 11785 11250
rect 11715 11190 11785 11210
rect 11845 11210 11940 11250
rect 11845 11190 11915 11210
rect 11630 11175 11686 11181
rect 11630 11115 11634 11175
rect 11715 11165 11915 11190
rect 11970 11181 12000 11369
rect 11944 11175 12000 11181
rect 11686 11115 11944 11135
rect 11996 11115 12000 11175
rect 11630 11105 12000 11115
rect 12030 11435 12400 11445
rect 12030 11375 12034 11435
rect 12086 11415 12344 11435
rect 12030 11369 12086 11375
rect 12030 11181 12060 11369
rect 12115 11360 12315 11385
rect 12396 11375 12400 11435
rect 12344 11369 12400 11375
rect 12115 11340 12185 11360
rect 12090 11300 12185 11340
rect 12245 11340 12315 11360
rect 12245 11300 12340 11340
rect 12090 11250 12340 11300
rect 12090 11210 12185 11250
rect 12115 11190 12185 11210
rect 12245 11210 12340 11250
rect 12245 11190 12315 11210
rect 12030 11175 12086 11181
rect 12030 11115 12034 11175
rect 12115 11165 12315 11190
rect 12370 11181 12400 11369
rect 12344 11175 12400 11181
rect 12086 11115 12344 11135
rect 12396 11115 12400 11175
rect 12030 11105 12400 11115
rect 12430 11435 12800 11445
rect 12430 11375 12434 11435
rect 12486 11415 12744 11435
rect 12430 11369 12486 11375
rect 12430 11181 12460 11369
rect 12515 11360 12715 11385
rect 12796 11375 12800 11435
rect 12744 11369 12800 11375
rect 12515 11340 12585 11360
rect 12490 11300 12585 11340
rect 12645 11340 12715 11360
rect 12645 11300 12740 11340
rect 12490 11250 12740 11300
rect 12490 11210 12585 11250
rect 12515 11190 12585 11210
rect 12645 11210 12740 11250
rect 12645 11190 12715 11210
rect 12430 11175 12486 11181
rect 12430 11115 12434 11175
rect 12515 11165 12715 11190
rect 12770 11181 12800 11369
rect 12744 11175 12800 11181
rect 12486 11115 12744 11135
rect 12796 11115 12800 11175
rect 12430 11105 12800 11115
rect 12830 11435 13200 11445
rect 12830 11375 12834 11435
rect 12886 11415 13144 11435
rect 12830 11369 12886 11375
rect 12830 11181 12860 11369
rect 12915 11360 13115 11385
rect 13196 11375 13200 11435
rect 13144 11369 13200 11375
rect 12915 11340 12985 11360
rect 12890 11300 12985 11340
rect 13045 11340 13115 11360
rect 13045 11300 13140 11340
rect 12890 11250 13140 11300
rect 12890 11210 12985 11250
rect 12915 11190 12985 11210
rect 13045 11210 13140 11250
rect 13045 11190 13115 11210
rect 12830 11175 12886 11181
rect 12830 11115 12834 11175
rect 12915 11165 13115 11190
rect 13170 11181 13200 11369
rect 13144 11175 13200 11181
rect 12886 11115 13144 11135
rect 13196 11115 13200 11175
rect 12830 11105 13200 11115
rect -370 11065 0 11075
rect -370 11005 -366 11065
rect -314 11045 -56 11065
rect -370 10999 -314 11005
rect -370 10811 -340 10999
rect -285 10990 -85 11015
rect -4 11005 0 11065
rect -56 10999 0 11005
rect -285 10970 -215 10990
rect -310 10930 -215 10970
rect -155 10970 -85 10990
rect -155 10930 -60 10970
rect -310 10880 -60 10930
rect -310 10840 -215 10880
rect -285 10820 -215 10840
rect -155 10840 -60 10880
rect -155 10820 -85 10840
rect -370 10805 -314 10811
rect -370 10745 -366 10805
rect -285 10795 -85 10820
rect -30 10811 0 10999
rect -56 10805 0 10811
rect -314 10745 -56 10765
rect -4 10745 0 10805
rect -370 10735 0 10745
rect 30 11065 400 11075
rect 30 11005 34 11065
rect 86 11045 344 11065
rect 30 10999 86 11005
rect 30 10811 60 10999
rect 115 10990 315 11015
rect 396 11005 400 11065
rect 344 10999 400 11005
rect 115 10970 185 10990
rect 90 10930 185 10970
rect 245 10970 315 10990
rect 245 10930 340 10970
rect 90 10880 340 10930
rect 90 10840 185 10880
rect 115 10820 185 10840
rect 245 10840 340 10880
rect 245 10820 315 10840
rect 30 10805 86 10811
rect 30 10745 34 10805
rect 115 10795 315 10820
rect 370 10811 400 10999
rect 344 10805 400 10811
rect 86 10745 344 10765
rect 396 10745 400 10805
rect 30 10735 400 10745
rect 430 11065 800 11075
rect 430 11005 434 11065
rect 486 11045 744 11065
rect 430 10999 486 11005
rect 430 10811 460 10999
rect 515 10990 715 11015
rect 796 11005 800 11065
rect 744 10999 800 11005
rect 515 10970 585 10990
rect 490 10930 585 10970
rect 645 10970 715 10990
rect 645 10930 740 10970
rect 490 10880 740 10930
rect 490 10840 585 10880
rect 515 10820 585 10840
rect 645 10840 740 10880
rect 645 10820 715 10840
rect 430 10805 486 10811
rect 430 10745 434 10805
rect 515 10795 715 10820
rect 770 10811 800 10999
rect 744 10805 800 10811
rect 486 10745 744 10765
rect 796 10745 800 10805
rect 430 10735 800 10745
rect 830 11065 1200 11075
rect 830 11005 834 11065
rect 886 11045 1144 11065
rect 830 10999 886 11005
rect 830 10811 860 10999
rect 915 10990 1115 11015
rect 1196 11005 1200 11065
rect 1144 10999 1200 11005
rect 915 10970 985 10990
rect 890 10930 985 10970
rect 1045 10970 1115 10990
rect 1045 10930 1140 10970
rect 890 10880 1140 10930
rect 890 10840 985 10880
rect 915 10820 985 10840
rect 1045 10840 1140 10880
rect 1045 10820 1115 10840
rect 830 10805 886 10811
rect 830 10745 834 10805
rect 915 10795 1115 10820
rect 1170 10811 1200 10999
rect 1144 10805 1200 10811
rect 886 10745 1144 10765
rect 1196 10745 1200 10805
rect 830 10735 1200 10745
rect 1230 11065 1600 11075
rect 1230 11005 1234 11065
rect 1286 11045 1544 11065
rect 1230 10999 1286 11005
rect 1230 10811 1260 10999
rect 1315 10990 1515 11015
rect 1596 11005 1600 11065
rect 1544 10999 1600 11005
rect 1315 10970 1385 10990
rect 1290 10930 1385 10970
rect 1445 10970 1515 10990
rect 1445 10930 1540 10970
rect 1290 10880 1540 10930
rect 1290 10840 1385 10880
rect 1315 10820 1385 10840
rect 1445 10840 1540 10880
rect 1445 10820 1515 10840
rect 1230 10805 1286 10811
rect 1230 10745 1234 10805
rect 1315 10795 1515 10820
rect 1570 10811 1600 10999
rect 1544 10805 1600 10811
rect 1286 10745 1544 10765
rect 1596 10745 1600 10805
rect 1230 10735 1600 10745
rect 1630 11065 2000 11075
rect 1630 11005 1634 11065
rect 1686 11045 1944 11065
rect 1630 10999 1686 11005
rect 1630 10811 1660 10999
rect 1715 10990 1915 11015
rect 1996 11005 2000 11065
rect 1944 10999 2000 11005
rect 1715 10970 1785 10990
rect 1690 10930 1785 10970
rect 1845 10970 1915 10990
rect 1845 10930 1940 10970
rect 1690 10880 1940 10930
rect 1690 10840 1785 10880
rect 1715 10820 1785 10840
rect 1845 10840 1940 10880
rect 1845 10820 1915 10840
rect 1630 10805 1686 10811
rect 1630 10745 1634 10805
rect 1715 10795 1915 10820
rect 1970 10811 2000 10999
rect 1944 10805 2000 10811
rect 1686 10745 1944 10765
rect 1996 10745 2000 10805
rect 1630 10735 2000 10745
rect 2030 11065 2400 11075
rect 2030 11005 2034 11065
rect 2086 11045 2344 11065
rect 2030 10999 2086 11005
rect 2030 10811 2060 10999
rect 2115 10990 2315 11015
rect 2396 11005 2400 11065
rect 2344 10999 2400 11005
rect 2115 10970 2185 10990
rect 2090 10930 2185 10970
rect 2245 10970 2315 10990
rect 2245 10930 2340 10970
rect 2090 10880 2340 10930
rect 2090 10840 2185 10880
rect 2115 10820 2185 10840
rect 2245 10840 2340 10880
rect 2245 10820 2315 10840
rect 2030 10805 2086 10811
rect 2030 10745 2034 10805
rect 2115 10795 2315 10820
rect 2370 10811 2400 10999
rect 2344 10805 2400 10811
rect 2086 10745 2344 10765
rect 2396 10745 2400 10805
rect 2030 10735 2400 10745
rect 2430 11065 2800 11075
rect 2430 11005 2434 11065
rect 2486 11045 2744 11065
rect 2430 10999 2486 11005
rect 2430 10811 2460 10999
rect 2515 10990 2715 11015
rect 2796 11005 2800 11065
rect 2744 10999 2800 11005
rect 2515 10970 2585 10990
rect 2490 10930 2585 10970
rect 2645 10970 2715 10990
rect 2645 10930 2740 10970
rect 2490 10880 2740 10930
rect 2490 10840 2585 10880
rect 2515 10820 2585 10840
rect 2645 10840 2740 10880
rect 2645 10820 2715 10840
rect 2430 10805 2486 10811
rect 2430 10745 2434 10805
rect 2515 10795 2715 10820
rect 2770 10811 2800 10999
rect 2744 10805 2800 10811
rect 2486 10745 2744 10765
rect 2796 10745 2800 10805
rect 2430 10735 2800 10745
rect 2830 11065 3200 11075
rect 2830 11005 2834 11065
rect 2886 11045 3144 11065
rect 2830 10999 2886 11005
rect 2830 10811 2860 10999
rect 2915 10990 3115 11015
rect 3196 11005 3200 11065
rect 3144 10999 3200 11005
rect 2915 10970 2985 10990
rect 2890 10930 2985 10970
rect 3045 10970 3115 10990
rect 3045 10930 3140 10970
rect 2890 10880 3140 10930
rect 2890 10840 2985 10880
rect 2915 10820 2985 10840
rect 3045 10840 3140 10880
rect 3045 10820 3115 10840
rect 2830 10805 2886 10811
rect 2830 10745 2834 10805
rect 2915 10795 3115 10820
rect 3170 10811 3200 10999
rect 3144 10805 3200 10811
rect 2886 10745 3144 10765
rect 3196 10745 3200 10805
rect 2830 10735 3200 10745
rect 3230 11065 3600 11075
rect 3230 11005 3234 11065
rect 3286 11045 3544 11065
rect 3230 10999 3286 11005
rect 3230 10811 3260 10999
rect 3315 10990 3515 11015
rect 3596 11005 3600 11065
rect 3544 10999 3600 11005
rect 3315 10970 3385 10990
rect 3290 10930 3385 10970
rect 3445 10970 3515 10990
rect 3445 10930 3540 10970
rect 3290 10880 3540 10930
rect 3290 10840 3385 10880
rect 3315 10820 3385 10840
rect 3445 10840 3540 10880
rect 3445 10820 3515 10840
rect 3230 10805 3286 10811
rect 3230 10745 3234 10805
rect 3315 10795 3515 10820
rect 3570 10811 3600 10999
rect 3544 10805 3600 10811
rect 3286 10745 3544 10765
rect 3596 10745 3600 10805
rect 3230 10735 3600 10745
rect 3630 11065 4000 11075
rect 3630 11005 3634 11065
rect 3686 11045 3944 11065
rect 3630 10999 3686 11005
rect 3630 10811 3660 10999
rect 3715 10990 3915 11015
rect 3996 11005 4000 11065
rect 3944 10999 4000 11005
rect 3715 10970 3785 10990
rect 3690 10930 3785 10970
rect 3845 10970 3915 10990
rect 3845 10930 3940 10970
rect 3690 10880 3940 10930
rect 3690 10840 3785 10880
rect 3715 10820 3785 10840
rect 3845 10840 3940 10880
rect 3845 10820 3915 10840
rect 3630 10805 3686 10811
rect 3630 10745 3634 10805
rect 3715 10795 3915 10820
rect 3970 10811 4000 10999
rect 3944 10805 4000 10811
rect 3686 10745 3944 10765
rect 3996 10745 4000 10805
rect 3630 10735 4000 10745
rect 4030 11065 4400 11075
rect 4030 11005 4034 11065
rect 4086 11045 4344 11065
rect 4030 10999 4086 11005
rect 4030 10811 4060 10999
rect 4115 10990 4315 11015
rect 4396 11005 4400 11065
rect 4344 10999 4400 11005
rect 4115 10970 4185 10990
rect 4090 10930 4185 10970
rect 4245 10970 4315 10990
rect 4245 10930 4340 10970
rect 4090 10880 4340 10930
rect 4090 10840 4185 10880
rect 4115 10820 4185 10840
rect 4245 10840 4340 10880
rect 4245 10820 4315 10840
rect 4030 10805 4086 10811
rect 4030 10745 4034 10805
rect 4115 10795 4315 10820
rect 4370 10811 4400 10999
rect 4344 10805 4400 10811
rect 4086 10745 4344 10765
rect 4396 10745 4400 10805
rect 4030 10735 4400 10745
rect 4430 11065 4800 11075
rect 4430 11005 4434 11065
rect 4486 11045 4744 11065
rect 4430 10999 4486 11005
rect 4430 10811 4460 10999
rect 4515 10990 4715 11015
rect 4796 11005 4800 11065
rect 4744 10999 4800 11005
rect 4515 10970 4585 10990
rect 4490 10930 4585 10970
rect 4645 10970 4715 10990
rect 4645 10930 4740 10970
rect 4490 10880 4740 10930
rect 4490 10840 4585 10880
rect 4515 10820 4585 10840
rect 4645 10840 4740 10880
rect 4645 10820 4715 10840
rect 4430 10805 4486 10811
rect 4430 10745 4434 10805
rect 4515 10795 4715 10820
rect 4770 10811 4800 10999
rect 4744 10805 4800 10811
rect 4486 10745 4744 10765
rect 4796 10745 4800 10805
rect 4430 10735 4800 10745
rect 4830 11065 5200 11075
rect 4830 11005 4834 11065
rect 4886 11045 5144 11065
rect 4830 10999 4886 11005
rect 4830 10811 4860 10999
rect 4915 10990 5115 11015
rect 5196 11005 5200 11065
rect 5144 10999 5200 11005
rect 4915 10970 4985 10990
rect 4890 10930 4985 10970
rect 5045 10970 5115 10990
rect 5045 10930 5140 10970
rect 4890 10880 5140 10930
rect 4890 10840 4985 10880
rect 4915 10820 4985 10840
rect 5045 10840 5140 10880
rect 5045 10820 5115 10840
rect 4830 10805 4886 10811
rect 4830 10745 4834 10805
rect 4915 10795 5115 10820
rect 5170 10811 5200 10999
rect 5144 10805 5200 10811
rect 4886 10745 5144 10765
rect 5196 10745 5200 10805
rect 4830 10735 5200 10745
rect 5230 11065 5600 11075
rect 5230 11005 5234 11065
rect 5286 11045 5544 11065
rect 5230 10999 5286 11005
rect 5230 10811 5260 10999
rect 5315 10990 5515 11015
rect 5596 11005 5600 11065
rect 5544 10999 5600 11005
rect 5315 10970 5385 10990
rect 5290 10930 5385 10970
rect 5445 10970 5515 10990
rect 5445 10930 5540 10970
rect 5290 10880 5540 10930
rect 5290 10840 5385 10880
rect 5315 10820 5385 10840
rect 5445 10840 5540 10880
rect 5445 10820 5515 10840
rect 5230 10805 5286 10811
rect 5230 10745 5234 10805
rect 5315 10795 5515 10820
rect 5570 10811 5600 10999
rect 5544 10805 5600 10811
rect 5286 10745 5544 10765
rect 5596 10745 5600 10805
rect 5230 10735 5600 10745
rect 5630 11065 6000 11075
rect 5630 11005 5634 11065
rect 5686 11045 5944 11065
rect 5630 10999 5686 11005
rect 5630 10811 5660 10999
rect 5715 10990 5915 11015
rect 5996 11005 6000 11065
rect 5944 10999 6000 11005
rect 5715 10970 5785 10990
rect 5690 10930 5785 10970
rect 5845 10970 5915 10990
rect 5845 10930 5940 10970
rect 5690 10880 5940 10930
rect 5690 10840 5785 10880
rect 5715 10820 5785 10840
rect 5845 10840 5940 10880
rect 5845 10820 5915 10840
rect 5630 10805 5686 10811
rect 5630 10745 5634 10805
rect 5715 10795 5915 10820
rect 5970 10811 6000 10999
rect 5944 10805 6000 10811
rect 5686 10745 5944 10765
rect 5996 10745 6000 10805
rect 5630 10735 6000 10745
rect 6030 11065 6400 11075
rect 6030 11005 6034 11065
rect 6086 11045 6344 11065
rect 6030 10999 6086 11005
rect 6030 10811 6060 10999
rect 6115 10990 6315 11015
rect 6396 11005 6400 11065
rect 6344 10999 6400 11005
rect 6115 10970 6185 10990
rect 6090 10930 6185 10970
rect 6245 10970 6315 10990
rect 6245 10930 6340 10970
rect 6090 10880 6340 10930
rect 6090 10840 6185 10880
rect 6115 10820 6185 10840
rect 6245 10840 6340 10880
rect 6245 10820 6315 10840
rect 6030 10805 6086 10811
rect 6030 10745 6034 10805
rect 6115 10795 6315 10820
rect 6370 10811 6400 10999
rect 6344 10805 6400 10811
rect 6086 10745 6344 10765
rect 6396 10745 6400 10805
rect 6030 10735 6400 10745
rect 6430 11065 6800 11075
rect 6430 11005 6434 11065
rect 6486 11045 6744 11065
rect 6430 10999 6486 11005
rect 6430 10811 6460 10999
rect 6515 10990 6715 11015
rect 6796 11005 6800 11065
rect 6744 10999 6800 11005
rect 6515 10970 6585 10990
rect 6490 10930 6585 10970
rect 6645 10970 6715 10990
rect 6645 10930 6740 10970
rect 6490 10880 6740 10930
rect 6490 10840 6585 10880
rect 6515 10820 6585 10840
rect 6645 10840 6740 10880
rect 6645 10820 6715 10840
rect 6430 10805 6486 10811
rect 6430 10745 6434 10805
rect 6515 10795 6715 10820
rect 6770 10811 6800 10999
rect 6744 10805 6800 10811
rect 6486 10745 6744 10765
rect 6796 10745 6800 10805
rect 6430 10735 6800 10745
rect 6830 11065 7200 11075
rect 6830 11005 6834 11065
rect 6886 11045 7144 11065
rect 6830 10999 6886 11005
rect 6830 10811 6860 10999
rect 6915 10990 7115 11015
rect 7196 11005 7200 11065
rect 7144 10999 7200 11005
rect 6915 10970 6985 10990
rect 6890 10930 6985 10970
rect 7045 10970 7115 10990
rect 7045 10930 7140 10970
rect 6890 10880 7140 10930
rect 6890 10840 6985 10880
rect 6915 10820 6985 10840
rect 7045 10840 7140 10880
rect 7045 10820 7115 10840
rect 6830 10805 6886 10811
rect 6830 10745 6834 10805
rect 6915 10795 7115 10820
rect 7170 10811 7200 10999
rect 7144 10805 7200 10811
rect 6886 10745 7144 10765
rect 7196 10745 7200 10805
rect 6830 10735 7200 10745
rect 7230 11065 7600 11075
rect 7230 11005 7234 11065
rect 7286 11045 7544 11065
rect 7230 10999 7286 11005
rect 7230 10811 7260 10999
rect 7315 10990 7515 11015
rect 7596 11005 7600 11065
rect 7544 10999 7600 11005
rect 7315 10970 7385 10990
rect 7290 10930 7385 10970
rect 7445 10970 7515 10990
rect 7445 10930 7540 10970
rect 7290 10880 7540 10930
rect 7290 10840 7385 10880
rect 7315 10820 7385 10840
rect 7445 10840 7540 10880
rect 7445 10820 7515 10840
rect 7230 10805 7286 10811
rect 7230 10745 7234 10805
rect 7315 10795 7515 10820
rect 7570 10811 7600 10999
rect 7544 10805 7600 10811
rect 7286 10745 7544 10765
rect 7596 10745 7600 10805
rect 7230 10735 7600 10745
rect 7630 11065 8000 11075
rect 7630 11005 7634 11065
rect 7686 11045 7944 11065
rect 7630 10999 7686 11005
rect 7630 10811 7660 10999
rect 7715 10990 7915 11015
rect 7996 11005 8000 11065
rect 7944 10999 8000 11005
rect 7715 10970 7785 10990
rect 7690 10930 7785 10970
rect 7845 10970 7915 10990
rect 7845 10930 7940 10970
rect 7690 10880 7940 10930
rect 7690 10840 7785 10880
rect 7715 10820 7785 10840
rect 7845 10840 7940 10880
rect 7845 10820 7915 10840
rect 7630 10805 7686 10811
rect 7630 10745 7634 10805
rect 7715 10795 7915 10820
rect 7970 10811 8000 10999
rect 7944 10805 8000 10811
rect 7686 10745 7944 10765
rect 7996 10745 8000 10805
rect 7630 10735 8000 10745
rect 8030 11065 8400 11075
rect 8030 11005 8034 11065
rect 8086 11045 8344 11065
rect 8030 10999 8086 11005
rect 8030 10811 8060 10999
rect 8115 10990 8315 11015
rect 8396 11005 8400 11065
rect 8344 10999 8400 11005
rect 8115 10970 8185 10990
rect 8090 10930 8185 10970
rect 8245 10970 8315 10990
rect 8245 10930 8340 10970
rect 8090 10880 8340 10930
rect 8090 10840 8185 10880
rect 8115 10820 8185 10840
rect 8245 10840 8340 10880
rect 8245 10820 8315 10840
rect 8030 10805 8086 10811
rect 8030 10745 8034 10805
rect 8115 10795 8315 10820
rect 8370 10811 8400 10999
rect 8344 10805 8400 10811
rect 8086 10745 8344 10765
rect 8396 10745 8400 10805
rect 8030 10735 8400 10745
rect 8430 11065 8800 11075
rect 8430 11005 8434 11065
rect 8486 11045 8744 11065
rect 8430 10999 8486 11005
rect 8430 10811 8460 10999
rect 8515 10990 8715 11015
rect 8796 11005 8800 11065
rect 8744 10999 8800 11005
rect 8515 10970 8585 10990
rect 8490 10930 8585 10970
rect 8645 10970 8715 10990
rect 8645 10930 8740 10970
rect 8490 10880 8740 10930
rect 8490 10840 8585 10880
rect 8515 10820 8585 10840
rect 8645 10840 8740 10880
rect 8645 10820 8715 10840
rect 8430 10805 8486 10811
rect 8430 10745 8434 10805
rect 8515 10795 8715 10820
rect 8770 10811 8800 10999
rect 8744 10805 8800 10811
rect 8486 10745 8744 10765
rect 8796 10745 8800 10805
rect 8430 10735 8800 10745
rect 8830 11065 9200 11075
rect 8830 11005 8834 11065
rect 8886 11045 9144 11065
rect 8830 10999 8886 11005
rect 8830 10811 8860 10999
rect 8915 10990 9115 11015
rect 9196 11005 9200 11065
rect 9144 10999 9200 11005
rect 8915 10970 8985 10990
rect 8890 10930 8985 10970
rect 9045 10970 9115 10990
rect 9045 10930 9140 10970
rect 8890 10880 9140 10930
rect 8890 10840 8985 10880
rect 8915 10820 8985 10840
rect 9045 10840 9140 10880
rect 9045 10820 9115 10840
rect 8830 10805 8886 10811
rect 8830 10745 8834 10805
rect 8915 10795 9115 10820
rect 9170 10811 9200 10999
rect 9144 10805 9200 10811
rect 8886 10745 9144 10765
rect 9196 10745 9200 10805
rect 8830 10735 9200 10745
rect 9230 11065 9600 11075
rect 9230 11005 9234 11065
rect 9286 11045 9544 11065
rect 9230 10999 9286 11005
rect 9230 10811 9260 10999
rect 9315 10990 9515 11015
rect 9596 11005 9600 11065
rect 9544 10999 9600 11005
rect 9315 10970 9385 10990
rect 9290 10930 9385 10970
rect 9445 10970 9515 10990
rect 9445 10930 9540 10970
rect 9290 10880 9540 10930
rect 9290 10840 9385 10880
rect 9315 10820 9385 10840
rect 9445 10840 9540 10880
rect 9445 10820 9515 10840
rect 9230 10805 9286 10811
rect 9230 10745 9234 10805
rect 9315 10795 9515 10820
rect 9570 10811 9600 10999
rect 9544 10805 9600 10811
rect 9286 10745 9544 10765
rect 9596 10745 9600 10805
rect 9230 10735 9600 10745
rect 9630 11065 10000 11075
rect 9630 11005 9634 11065
rect 9686 11045 9944 11065
rect 9630 10999 9686 11005
rect 9630 10811 9660 10999
rect 9715 10990 9915 11015
rect 9996 11005 10000 11065
rect 9944 10999 10000 11005
rect 9715 10970 9785 10990
rect 9690 10930 9785 10970
rect 9845 10970 9915 10990
rect 9845 10930 9940 10970
rect 9690 10880 9940 10930
rect 9690 10840 9785 10880
rect 9715 10820 9785 10840
rect 9845 10840 9940 10880
rect 9845 10820 9915 10840
rect 9630 10805 9686 10811
rect 9630 10745 9634 10805
rect 9715 10795 9915 10820
rect 9970 10811 10000 10999
rect 9944 10805 10000 10811
rect 9686 10745 9944 10765
rect 9996 10745 10000 10805
rect 9630 10735 10000 10745
rect 10030 11065 10400 11075
rect 10030 11005 10034 11065
rect 10086 11045 10344 11065
rect 10030 10999 10086 11005
rect 10030 10811 10060 10999
rect 10115 10990 10315 11015
rect 10396 11005 10400 11065
rect 10344 10999 10400 11005
rect 10115 10970 10185 10990
rect 10090 10930 10185 10970
rect 10245 10970 10315 10990
rect 10245 10930 10340 10970
rect 10090 10880 10340 10930
rect 10090 10840 10185 10880
rect 10115 10820 10185 10840
rect 10245 10840 10340 10880
rect 10245 10820 10315 10840
rect 10030 10805 10086 10811
rect 10030 10745 10034 10805
rect 10115 10795 10315 10820
rect 10370 10811 10400 10999
rect 10344 10805 10400 10811
rect 10086 10745 10344 10765
rect 10396 10745 10400 10805
rect 10030 10735 10400 10745
rect 10430 11065 10800 11075
rect 10430 11005 10434 11065
rect 10486 11045 10744 11065
rect 10430 10999 10486 11005
rect 10430 10811 10460 10999
rect 10515 10990 10715 11015
rect 10796 11005 10800 11065
rect 10744 10999 10800 11005
rect 10515 10970 10585 10990
rect 10490 10930 10585 10970
rect 10645 10970 10715 10990
rect 10645 10930 10740 10970
rect 10490 10880 10740 10930
rect 10490 10840 10585 10880
rect 10515 10820 10585 10840
rect 10645 10840 10740 10880
rect 10645 10820 10715 10840
rect 10430 10805 10486 10811
rect 10430 10745 10434 10805
rect 10515 10795 10715 10820
rect 10770 10811 10800 10999
rect 10744 10805 10800 10811
rect 10486 10745 10744 10765
rect 10796 10745 10800 10805
rect 10430 10735 10800 10745
rect 10830 11065 11200 11075
rect 10830 11005 10834 11065
rect 10886 11045 11144 11065
rect 10830 10999 10886 11005
rect 10830 10811 10860 10999
rect 10915 10990 11115 11015
rect 11196 11005 11200 11065
rect 11144 10999 11200 11005
rect 10915 10970 10985 10990
rect 10890 10930 10985 10970
rect 11045 10970 11115 10990
rect 11045 10930 11140 10970
rect 10890 10880 11140 10930
rect 10890 10840 10985 10880
rect 10915 10820 10985 10840
rect 11045 10840 11140 10880
rect 11045 10820 11115 10840
rect 10830 10805 10886 10811
rect 10830 10745 10834 10805
rect 10915 10795 11115 10820
rect 11170 10811 11200 10999
rect 11144 10805 11200 10811
rect 10886 10745 11144 10765
rect 11196 10745 11200 10805
rect 10830 10735 11200 10745
rect 11230 11065 11600 11075
rect 11230 11005 11234 11065
rect 11286 11045 11544 11065
rect 11230 10999 11286 11005
rect 11230 10811 11260 10999
rect 11315 10990 11515 11015
rect 11596 11005 11600 11065
rect 11544 10999 11600 11005
rect 11315 10970 11385 10990
rect 11290 10930 11385 10970
rect 11445 10970 11515 10990
rect 11445 10930 11540 10970
rect 11290 10880 11540 10930
rect 11290 10840 11385 10880
rect 11315 10820 11385 10840
rect 11445 10840 11540 10880
rect 11445 10820 11515 10840
rect 11230 10805 11286 10811
rect 11230 10745 11234 10805
rect 11315 10795 11515 10820
rect 11570 10811 11600 10999
rect 11544 10805 11600 10811
rect 11286 10745 11544 10765
rect 11596 10745 11600 10805
rect 11230 10735 11600 10745
rect 11630 11065 12000 11075
rect 11630 11005 11634 11065
rect 11686 11045 11944 11065
rect 11630 10999 11686 11005
rect 11630 10811 11660 10999
rect 11715 10990 11915 11015
rect 11996 11005 12000 11065
rect 11944 10999 12000 11005
rect 11715 10970 11785 10990
rect 11690 10930 11785 10970
rect 11845 10970 11915 10990
rect 11845 10930 11940 10970
rect 11690 10880 11940 10930
rect 11690 10840 11785 10880
rect 11715 10820 11785 10840
rect 11845 10840 11940 10880
rect 11845 10820 11915 10840
rect 11630 10805 11686 10811
rect 11630 10745 11634 10805
rect 11715 10795 11915 10820
rect 11970 10811 12000 10999
rect 11944 10805 12000 10811
rect 11686 10745 11944 10765
rect 11996 10745 12000 10805
rect 11630 10735 12000 10745
rect 12030 11065 12400 11075
rect 12030 11005 12034 11065
rect 12086 11045 12344 11065
rect 12030 10999 12086 11005
rect 12030 10811 12060 10999
rect 12115 10990 12315 11015
rect 12396 11005 12400 11065
rect 12344 10999 12400 11005
rect 12115 10970 12185 10990
rect 12090 10930 12185 10970
rect 12245 10970 12315 10990
rect 12245 10930 12340 10970
rect 12090 10880 12340 10930
rect 12090 10840 12185 10880
rect 12115 10820 12185 10840
rect 12245 10840 12340 10880
rect 12245 10820 12315 10840
rect 12030 10805 12086 10811
rect 12030 10745 12034 10805
rect 12115 10795 12315 10820
rect 12370 10811 12400 10999
rect 12344 10805 12400 10811
rect 12086 10745 12344 10765
rect 12396 10745 12400 10805
rect 12030 10735 12400 10745
rect 12430 11065 12800 11075
rect 12430 11005 12434 11065
rect 12486 11045 12744 11065
rect 12430 10999 12486 11005
rect 12430 10811 12460 10999
rect 12515 10990 12715 11015
rect 12796 11005 12800 11065
rect 12744 10999 12800 11005
rect 12515 10970 12585 10990
rect 12490 10930 12585 10970
rect 12645 10970 12715 10990
rect 12645 10930 12740 10970
rect 12490 10880 12740 10930
rect 12490 10840 12585 10880
rect 12515 10820 12585 10840
rect 12645 10840 12740 10880
rect 12645 10820 12715 10840
rect 12430 10805 12486 10811
rect 12430 10745 12434 10805
rect 12515 10795 12715 10820
rect 12770 10811 12800 10999
rect 12744 10805 12800 10811
rect 12486 10745 12744 10765
rect 12796 10745 12800 10805
rect 12430 10735 12800 10745
rect 12830 11065 13200 11075
rect 12830 11005 12834 11065
rect 12886 11045 13144 11065
rect 12830 10999 12886 11005
rect 12830 10811 12860 10999
rect 12915 10990 13115 11015
rect 13196 11005 13200 11065
rect 13144 10999 13200 11005
rect 12915 10970 12985 10990
rect 12890 10930 12985 10970
rect 13045 10970 13115 10990
rect 13045 10930 13140 10970
rect 12890 10880 13140 10930
rect 12890 10840 12985 10880
rect 12915 10820 12985 10840
rect 13045 10840 13140 10880
rect 13045 10820 13115 10840
rect 12830 10805 12886 10811
rect 12830 10745 12834 10805
rect 12915 10795 13115 10820
rect 13170 10811 13200 10999
rect 13144 10805 13200 10811
rect 12886 10745 13144 10765
rect 13196 10745 13200 10805
rect 12830 10735 13200 10745
rect -370 10695 0 10705
rect -370 10635 -366 10695
rect -314 10675 -56 10695
rect -370 10629 -314 10635
rect -370 10441 -340 10629
rect -285 10620 -85 10645
rect -4 10635 0 10695
rect -56 10629 0 10635
rect -285 10600 -215 10620
rect -310 10560 -215 10600
rect -155 10600 -85 10620
rect -155 10560 -60 10600
rect -310 10510 -60 10560
rect -310 10470 -215 10510
rect -285 10450 -215 10470
rect -155 10470 -60 10510
rect -155 10450 -85 10470
rect -370 10435 -314 10441
rect -370 10375 -366 10435
rect -285 10425 -85 10450
rect -30 10441 0 10629
rect -56 10435 0 10441
rect -314 10375 -56 10395
rect -4 10375 0 10435
rect -370 10365 0 10375
rect 30 10695 400 10705
rect 30 10635 34 10695
rect 86 10675 344 10695
rect 30 10629 86 10635
rect 30 10441 60 10629
rect 115 10620 315 10645
rect 396 10635 400 10695
rect 344 10629 400 10635
rect 115 10600 185 10620
rect 90 10560 185 10600
rect 245 10600 315 10620
rect 245 10560 340 10600
rect 90 10510 340 10560
rect 90 10470 185 10510
rect 115 10450 185 10470
rect 245 10470 340 10510
rect 245 10450 315 10470
rect 30 10435 86 10441
rect 30 10375 34 10435
rect 115 10425 315 10450
rect 370 10441 400 10629
rect 344 10435 400 10441
rect 86 10375 344 10395
rect 396 10375 400 10435
rect 30 10365 400 10375
rect 430 10695 800 10705
rect 430 10635 434 10695
rect 486 10675 744 10695
rect 430 10629 486 10635
rect 430 10441 460 10629
rect 515 10620 715 10645
rect 796 10635 800 10695
rect 744 10629 800 10635
rect 515 10600 585 10620
rect 490 10560 585 10600
rect 645 10600 715 10620
rect 645 10560 740 10600
rect 490 10510 740 10560
rect 490 10470 585 10510
rect 515 10450 585 10470
rect 645 10470 740 10510
rect 645 10450 715 10470
rect 430 10435 486 10441
rect 430 10375 434 10435
rect 515 10425 715 10450
rect 770 10441 800 10629
rect 744 10435 800 10441
rect 486 10375 744 10395
rect 796 10375 800 10435
rect 430 10365 800 10375
rect 830 10695 1200 10705
rect 830 10635 834 10695
rect 886 10675 1144 10695
rect 830 10629 886 10635
rect 830 10441 860 10629
rect 915 10620 1115 10645
rect 1196 10635 1200 10695
rect 1144 10629 1200 10635
rect 915 10600 985 10620
rect 890 10560 985 10600
rect 1045 10600 1115 10620
rect 1045 10560 1140 10600
rect 890 10510 1140 10560
rect 890 10470 985 10510
rect 915 10450 985 10470
rect 1045 10470 1140 10510
rect 1045 10450 1115 10470
rect 830 10435 886 10441
rect 830 10375 834 10435
rect 915 10425 1115 10450
rect 1170 10441 1200 10629
rect 1144 10435 1200 10441
rect 886 10375 1144 10395
rect 1196 10375 1200 10435
rect 830 10365 1200 10375
rect 1230 10695 1600 10705
rect 1230 10635 1234 10695
rect 1286 10675 1544 10695
rect 1230 10629 1286 10635
rect 1230 10441 1260 10629
rect 1315 10620 1515 10645
rect 1596 10635 1600 10695
rect 1544 10629 1600 10635
rect 1315 10600 1385 10620
rect 1290 10560 1385 10600
rect 1445 10600 1515 10620
rect 1445 10560 1540 10600
rect 1290 10510 1540 10560
rect 1290 10470 1385 10510
rect 1315 10450 1385 10470
rect 1445 10470 1540 10510
rect 1445 10450 1515 10470
rect 1230 10435 1286 10441
rect 1230 10375 1234 10435
rect 1315 10425 1515 10450
rect 1570 10441 1600 10629
rect 1544 10435 1600 10441
rect 1286 10375 1544 10395
rect 1596 10375 1600 10435
rect 1230 10365 1600 10375
rect 1630 10695 2000 10705
rect 1630 10635 1634 10695
rect 1686 10675 1944 10695
rect 1630 10629 1686 10635
rect 1630 10441 1660 10629
rect 1715 10620 1915 10645
rect 1996 10635 2000 10695
rect 1944 10629 2000 10635
rect 1715 10600 1785 10620
rect 1690 10560 1785 10600
rect 1845 10600 1915 10620
rect 1845 10560 1940 10600
rect 1690 10510 1940 10560
rect 1690 10470 1785 10510
rect 1715 10450 1785 10470
rect 1845 10470 1940 10510
rect 1845 10450 1915 10470
rect 1630 10435 1686 10441
rect 1630 10375 1634 10435
rect 1715 10425 1915 10450
rect 1970 10441 2000 10629
rect 1944 10435 2000 10441
rect 1686 10375 1944 10395
rect 1996 10375 2000 10435
rect 1630 10365 2000 10375
rect 2030 10695 2400 10705
rect 2030 10635 2034 10695
rect 2086 10675 2344 10695
rect 2030 10629 2086 10635
rect 2030 10441 2060 10629
rect 2115 10620 2315 10645
rect 2396 10635 2400 10695
rect 2344 10629 2400 10635
rect 2115 10600 2185 10620
rect 2090 10560 2185 10600
rect 2245 10600 2315 10620
rect 2245 10560 2340 10600
rect 2090 10510 2340 10560
rect 2090 10470 2185 10510
rect 2115 10450 2185 10470
rect 2245 10470 2340 10510
rect 2245 10450 2315 10470
rect 2030 10435 2086 10441
rect 2030 10375 2034 10435
rect 2115 10425 2315 10450
rect 2370 10441 2400 10629
rect 2344 10435 2400 10441
rect 2086 10375 2344 10395
rect 2396 10375 2400 10435
rect 2030 10365 2400 10375
rect 2430 10695 2800 10705
rect 2430 10635 2434 10695
rect 2486 10675 2744 10695
rect 2430 10629 2486 10635
rect 2430 10441 2460 10629
rect 2515 10620 2715 10645
rect 2796 10635 2800 10695
rect 2744 10629 2800 10635
rect 2515 10600 2585 10620
rect 2490 10560 2585 10600
rect 2645 10600 2715 10620
rect 2645 10560 2740 10600
rect 2490 10510 2740 10560
rect 2490 10470 2585 10510
rect 2515 10450 2585 10470
rect 2645 10470 2740 10510
rect 2645 10450 2715 10470
rect 2430 10435 2486 10441
rect 2430 10375 2434 10435
rect 2515 10425 2715 10450
rect 2770 10441 2800 10629
rect 2744 10435 2800 10441
rect 2486 10375 2744 10395
rect 2796 10375 2800 10435
rect 2430 10365 2800 10375
rect 2830 10695 3200 10705
rect 2830 10635 2834 10695
rect 2886 10675 3144 10695
rect 2830 10629 2886 10635
rect 2830 10441 2860 10629
rect 2915 10620 3115 10645
rect 3196 10635 3200 10695
rect 3144 10629 3200 10635
rect 2915 10600 2985 10620
rect 2890 10560 2985 10600
rect 3045 10600 3115 10620
rect 3045 10560 3140 10600
rect 2890 10510 3140 10560
rect 2890 10470 2985 10510
rect 2915 10450 2985 10470
rect 3045 10470 3140 10510
rect 3045 10450 3115 10470
rect 2830 10435 2886 10441
rect 2830 10375 2834 10435
rect 2915 10425 3115 10450
rect 3170 10441 3200 10629
rect 3144 10435 3200 10441
rect 2886 10375 3144 10395
rect 3196 10375 3200 10435
rect 2830 10365 3200 10375
rect 3230 10695 3600 10705
rect 3230 10635 3234 10695
rect 3286 10675 3544 10695
rect 3230 10629 3286 10635
rect 3230 10441 3260 10629
rect 3315 10620 3515 10645
rect 3596 10635 3600 10695
rect 3544 10629 3600 10635
rect 3315 10600 3385 10620
rect 3290 10560 3385 10600
rect 3445 10600 3515 10620
rect 3445 10560 3540 10600
rect 3290 10510 3540 10560
rect 3290 10470 3385 10510
rect 3315 10450 3385 10470
rect 3445 10470 3540 10510
rect 3445 10450 3515 10470
rect 3230 10435 3286 10441
rect 3230 10375 3234 10435
rect 3315 10425 3515 10450
rect 3570 10441 3600 10629
rect 3544 10435 3600 10441
rect 3286 10375 3544 10395
rect 3596 10375 3600 10435
rect 3230 10365 3600 10375
rect 3630 10695 4000 10705
rect 3630 10635 3634 10695
rect 3686 10675 3944 10695
rect 3630 10629 3686 10635
rect 3630 10441 3660 10629
rect 3715 10620 3915 10645
rect 3996 10635 4000 10695
rect 3944 10629 4000 10635
rect 3715 10600 3785 10620
rect 3690 10560 3785 10600
rect 3845 10600 3915 10620
rect 3845 10560 3940 10600
rect 3690 10510 3940 10560
rect 3690 10470 3785 10510
rect 3715 10450 3785 10470
rect 3845 10470 3940 10510
rect 3845 10450 3915 10470
rect 3630 10435 3686 10441
rect 3630 10375 3634 10435
rect 3715 10425 3915 10450
rect 3970 10441 4000 10629
rect 3944 10435 4000 10441
rect 3686 10375 3944 10395
rect 3996 10375 4000 10435
rect 3630 10365 4000 10375
rect 4030 10695 4400 10705
rect 4030 10635 4034 10695
rect 4086 10675 4344 10695
rect 4030 10629 4086 10635
rect 4030 10441 4060 10629
rect 4115 10620 4315 10645
rect 4396 10635 4400 10695
rect 4344 10629 4400 10635
rect 4115 10600 4185 10620
rect 4090 10560 4185 10600
rect 4245 10600 4315 10620
rect 4245 10560 4340 10600
rect 4090 10510 4340 10560
rect 4090 10470 4185 10510
rect 4115 10450 4185 10470
rect 4245 10470 4340 10510
rect 4245 10450 4315 10470
rect 4030 10435 4086 10441
rect 4030 10375 4034 10435
rect 4115 10425 4315 10450
rect 4370 10441 4400 10629
rect 4344 10435 4400 10441
rect 4086 10375 4344 10395
rect 4396 10375 4400 10435
rect 4030 10365 4400 10375
rect 4430 10695 4800 10705
rect 4430 10635 4434 10695
rect 4486 10675 4744 10695
rect 4430 10629 4486 10635
rect 4430 10441 4460 10629
rect 4515 10620 4715 10645
rect 4796 10635 4800 10695
rect 4744 10629 4800 10635
rect 4515 10600 4585 10620
rect 4490 10560 4585 10600
rect 4645 10600 4715 10620
rect 4645 10560 4740 10600
rect 4490 10510 4740 10560
rect 4490 10470 4585 10510
rect 4515 10450 4585 10470
rect 4645 10470 4740 10510
rect 4645 10450 4715 10470
rect 4430 10435 4486 10441
rect 4430 10375 4434 10435
rect 4515 10425 4715 10450
rect 4770 10441 4800 10629
rect 4744 10435 4800 10441
rect 4486 10375 4744 10395
rect 4796 10375 4800 10435
rect 4430 10365 4800 10375
rect 4830 10695 5200 10705
rect 4830 10635 4834 10695
rect 4886 10675 5144 10695
rect 4830 10629 4886 10635
rect 4830 10441 4860 10629
rect 4915 10620 5115 10645
rect 5196 10635 5200 10695
rect 5144 10629 5200 10635
rect 4915 10600 4985 10620
rect 4890 10560 4985 10600
rect 5045 10600 5115 10620
rect 5045 10560 5140 10600
rect 4890 10510 5140 10560
rect 4890 10470 4985 10510
rect 4915 10450 4985 10470
rect 5045 10470 5140 10510
rect 5045 10450 5115 10470
rect 4830 10435 4886 10441
rect 4830 10375 4834 10435
rect 4915 10425 5115 10450
rect 5170 10441 5200 10629
rect 5144 10435 5200 10441
rect 4886 10375 5144 10395
rect 5196 10375 5200 10435
rect 4830 10365 5200 10375
rect 5230 10695 5600 10705
rect 5230 10635 5234 10695
rect 5286 10675 5544 10695
rect 5230 10629 5286 10635
rect 5230 10441 5260 10629
rect 5315 10620 5515 10645
rect 5596 10635 5600 10695
rect 5544 10629 5600 10635
rect 5315 10600 5385 10620
rect 5290 10560 5385 10600
rect 5445 10600 5515 10620
rect 5445 10560 5540 10600
rect 5290 10510 5540 10560
rect 5290 10470 5385 10510
rect 5315 10450 5385 10470
rect 5445 10470 5540 10510
rect 5445 10450 5515 10470
rect 5230 10435 5286 10441
rect 5230 10375 5234 10435
rect 5315 10425 5515 10450
rect 5570 10441 5600 10629
rect 5544 10435 5600 10441
rect 5286 10375 5544 10395
rect 5596 10375 5600 10435
rect 5230 10365 5600 10375
rect 5630 10695 6000 10705
rect 5630 10635 5634 10695
rect 5686 10675 5944 10695
rect 5630 10629 5686 10635
rect 5630 10441 5660 10629
rect 5715 10620 5915 10645
rect 5996 10635 6000 10695
rect 5944 10629 6000 10635
rect 5715 10600 5785 10620
rect 5690 10560 5785 10600
rect 5845 10600 5915 10620
rect 5845 10560 5940 10600
rect 5690 10510 5940 10560
rect 5690 10470 5785 10510
rect 5715 10450 5785 10470
rect 5845 10470 5940 10510
rect 5845 10450 5915 10470
rect 5630 10435 5686 10441
rect 5630 10375 5634 10435
rect 5715 10425 5915 10450
rect 5970 10441 6000 10629
rect 5944 10435 6000 10441
rect 5686 10375 5944 10395
rect 5996 10375 6000 10435
rect 5630 10365 6000 10375
rect 6030 10695 6400 10705
rect 6030 10635 6034 10695
rect 6086 10675 6344 10695
rect 6030 10629 6086 10635
rect 6030 10441 6060 10629
rect 6115 10620 6315 10645
rect 6396 10635 6400 10695
rect 6344 10629 6400 10635
rect 6115 10600 6185 10620
rect 6090 10560 6185 10600
rect 6245 10600 6315 10620
rect 6245 10560 6340 10600
rect 6090 10510 6340 10560
rect 6090 10470 6185 10510
rect 6115 10450 6185 10470
rect 6245 10470 6340 10510
rect 6245 10450 6315 10470
rect 6030 10435 6086 10441
rect 6030 10375 6034 10435
rect 6115 10425 6315 10450
rect 6370 10441 6400 10629
rect 6344 10435 6400 10441
rect 6086 10375 6344 10395
rect 6396 10375 6400 10435
rect 6030 10365 6400 10375
rect 6430 10695 6800 10705
rect 6430 10635 6434 10695
rect 6486 10675 6744 10695
rect 6430 10629 6486 10635
rect 6430 10441 6460 10629
rect 6515 10620 6715 10645
rect 6796 10635 6800 10695
rect 6744 10629 6800 10635
rect 6515 10600 6585 10620
rect 6490 10560 6585 10600
rect 6645 10600 6715 10620
rect 6645 10560 6740 10600
rect 6490 10510 6740 10560
rect 6490 10470 6585 10510
rect 6515 10450 6585 10470
rect 6645 10470 6740 10510
rect 6645 10450 6715 10470
rect 6430 10435 6486 10441
rect 6430 10375 6434 10435
rect 6515 10425 6715 10450
rect 6770 10441 6800 10629
rect 6744 10435 6800 10441
rect 6486 10375 6744 10395
rect 6796 10375 6800 10435
rect 6430 10365 6800 10375
rect 6830 10695 7200 10705
rect 6830 10635 6834 10695
rect 6886 10675 7144 10695
rect 6830 10629 6886 10635
rect 6830 10441 6860 10629
rect 6915 10620 7115 10645
rect 7196 10635 7200 10695
rect 7144 10629 7200 10635
rect 6915 10600 6985 10620
rect 6890 10560 6985 10600
rect 7045 10600 7115 10620
rect 7045 10560 7140 10600
rect 6890 10510 7140 10560
rect 6890 10470 6985 10510
rect 6915 10450 6985 10470
rect 7045 10470 7140 10510
rect 7045 10450 7115 10470
rect 6830 10435 6886 10441
rect 6830 10375 6834 10435
rect 6915 10425 7115 10450
rect 7170 10441 7200 10629
rect 7144 10435 7200 10441
rect 6886 10375 7144 10395
rect 7196 10375 7200 10435
rect 6830 10365 7200 10375
rect 7230 10695 7600 10705
rect 7230 10635 7234 10695
rect 7286 10675 7544 10695
rect 7230 10629 7286 10635
rect 7230 10441 7260 10629
rect 7315 10620 7515 10645
rect 7596 10635 7600 10695
rect 7544 10629 7600 10635
rect 7315 10600 7385 10620
rect 7290 10560 7385 10600
rect 7445 10600 7515 10620
rect 7445 10560 7540 10600
rect 7290 10510 7540 10560
rect 7290 10470 7385 10510
rect 7315 10450 7385 10470
rect 7445 10470 7540 10510
rect 7445 10450 7515 10470
rect 7230 10435 7286 10441
rect 7230 10375 7234 10435
rect 7315 10425 7515 10450
rect 7570 10441 7600 10629
rect 7544 10435 7600 10441
rect 7286 10375 7544 10395
rect 7596 10375 7600 10435
rect 7230 10365 7600 10375
rect 7630 10695 8000 10705
rect 7630 10635 7634 10695
rect 7686 10675 7944 10695
rect 7630 10629 7686 10635
rect 7630 10441 7660 10629
rect 7715 10620 7915 10645
rect 7996 10635 8000 10695
rect 7944 10629 8000 10635
rect 7715 10600 7785 10620
rect 7690 10560 7785 10600
rect 7845 10600 7915 10620
rect 7845 10560 7940 10600
rect 7690 10510 7940 10560
rect 7690 10470 7785 10510
rect 7715 10450 7785 10470
rect 7845 10470 7940 10510
rect 7845 10450 7915 10470
rect 7630 10435 7686 10441
rect 7630 10375 7634 10435
rect 7715 10425 7915 10450
rect 7970 10441 8000 10629
rect 7944 10435 8000 10441
rect 7686 10375 7944 10395
rect 7996 10375 8000 10435
rect 7630 10365 8000 10375
rect 8030 10695 8400 10705
rect 8030 10635 8034 10695
rect 8086 10675 8344 10695
rect 8030 10629 8086 10635
rect 8030 10441 8060 10629
rect 8115 10620 8315 10645
rect 8396 10635 8400 10695
rect 8344 10629 8400 10635
rect 8115 10600 8185 10620
rect 8090 10560 8185 10600
rect 8245 10600 8315 10620
rect 8245 10560 8340 10600
rect 8090 10510 8340 10560
rect 8090 10470 8185 10510
rect 8115 10450 8185 10470
rect 8245 10470 8340 10510
rect 8245 10450 8315 10470
rect 8030 10435 8086 10441
rect 8030 10375 8034 10435
rect 8115 10425 8315 10450
rect 8370 10441 8400 10629
rect 8344 10435 8400 10441
rect 8086 10375 8344 10395
rect 8396 10375 8400 10435
rect 8030 10365 8400 10375
rect 8430 10695 8800 10705
rect 8430 10635 8434 10695
rect 8486 10675 8744 10695
rect 8430 10629 8486 10635
rect 8430 10441 8460 10629
rect 8515 10620 8715 10645
rect 8796 10635 8800 10695
rect 8744 10629 8800 10635
rect 8515 10600 8585 10620
rect 8490 10560 8585 10600
rect 8645 10600 8715 10620
rect 8645 10560 8740 10600
rect 8490 10510 8740 10560
rect 8490 10470 8585 10510
rect 8515 10450 8585 10470
rect 8645 10470 8740 10510
rect 8645 10450 8715 10470
rect 8430 10435 8486 10441
rect 8430 10375 8434 10435
rect 8515 10425 8715 10450
rect 8770 10441 8800 10629
rect 8744 10435 8800 10441
rect 8486 10375 8744 10395
rect 8796 10375 8800 10435
rect 8430 10365 8800 10375
rect 8830 10695 9200 10705
rect 8830 10635 8834 10695
rect 8886 10675 9144 10695
rect 8830 10629 8886 10635
rect 8830 10441 8860 10629
rect 8915 10620 9115 10645
rect 9196 10635 9200 10695
rect 9144 10629 9200 10635
rect 8915 10600 8985 10620
rect 8890 10560 8985 10600
rect 9045 10600 9115 10620
rect 9045 10560 9140 10600
rect 8890 10510 9140 10560
rect 8890 10470 8985 10510
rect 8915 10450 8985 10470
rect 9045 10470 9140 10510
rect 9045 10450 9115 10470
rect 8830 10435 8886 10441
rect 8830 10375 8834 10435
rect 8915 10425 9115 10450
rect 9170 10441 9200 10629
rect 9144 10435 9200 10441
rect 8886 10375 9144 10395
rect 9196 10375 9200 10435
rect 8830 10365 9200 10375
rect 9230 10695 9600 10705
rect 9230 10635 9234 10695
rect 9286 10675 9544 10695
rect 9230 10629 9286 10635
rect 9230 10441 9260 10629
rect 9315 10620 9515 10645
rect 9596 10635 9600 10695
rect 9544 10629 9600 10635
rect 9315 10600 9385 10620
rect 9290 10560 9385 10600
rect 9445 10600 9515 10620
rect 9445 10560 9540 10600
rect 9290 10510 9540 10560
rect 9290 10470 9385 10510
rect 9315 10450 9385 10470
rect 9445 10470 9540 10510
rect 9445 10450 9515 10470
rect 9230 10435 9286 10441
rect 9230 10375 9234 10435
rect 9315 10425 9515 10450
rect 9570 10441 9600 10629
rect 9544 10435 9600 10441
rect 9286 10375 9544 10395
rect 9596 10375 9600 10435
rect 9230 10365 9600 10375
rect 9630 10695 10000 10705
rect 9630 10635 9634 10695
rect 9686 10675 9944 10695
rect 9630 10629 9686 10635
rect 9630 10441 9660 10629
rect 9715 10620 9915 10645
rect 9996 10635 10000 10695
rect 9944 10629 10000 10635
rect 9715 10600 9785 10620
rect 9690 10560 9785 10600
rect 9845 10600 9915 10620
rect 9845 10560 9940 10600
rect 9690 10510 9940 10560
rect 9690 10470 9785 10510
rect 9715 10450 9785 10470
rect 9845 10470 9940 10510
rect 9845 10450 9915 10470
rect 9630 10435 9686 10441
rect 9630 10375 9634 10435
rect 9715 10425 9915 10450
rect 9970 10441 10000 10629
rect 9944 10435 10000 10441
rect 9686 10375 9944 10395
rect 9996 10375 10000 10435
rect 9630 10365 10000 10375
rect 10030 10695 10400 10705
rect 10030 10635 10034 10695
rect 10086 10675 10344 10695
rect 10030 10629 10086 10635
rect 10030 10441 10060 10629
rect 10115 10620 10315 10645
rect 10396 10635 10400 10695
rect 10344 10629 10400 10635
rect 10115 10600 10185 10620
rect 10090 10560 10185 10600
rect 10245 10600 10315 10620
rect 10245 10560 10340 10600
rect 10090 10510 10340 10560
rect 10090 10470 10185 10510
rect 10115 10450 10185 10470
rect 10245 10470 10340 10510
rect 10245 10450 10315 10470
rect 10030 10435 10086 10441
rect 10030 10375 10034 10435
rect 10115 10425 10315 10450
rect 10370 10441 10400 10629
rect 10344 10435 10400 10441
rect 10086 10375 10344 10395
rect 10396 10375 10400 10435
rect 10030 10365 10400 10375
rect 10430 10695 10800 10705
rect 10430 10635 10434 10695
rect 10486 10675 10744 10695
rect 10430 10629 10486 10635
rect 10430 10441 10460 10629
rect 10515 10620 10715 10645
rect 10796 10635 10800 10695
rect 10744 10629 10800 10635
rect 10515 10600 10585 10620
rect 10490 10560 10585 10600
rect 10645 10600 10715 10620
rect 10645 10560 10740 10600
rect 10490 10510 10740 10560
rect 10490 10470 10585 10510
rect 10515 10450 10585 10470
rect 10645 10470 10740 10510
rect 10645 10450 10715 10470
rect 10430 10435 10486 10441
rect 10430 10375 10434 10435
rect 10515 10425 10715 10450
rect 10770 10441 10800 10629
rect 10744 10435 10800 10441
rect 10486 10375 10744 10395
rect 10796 10375 10800 10435
rect 10430 10365 10800 10375
rect 10830 10695 11200 10705
rect 10830 10635 10834 10695
rect 10886 10675 11144 10695
rect 10830 10629 10886 10635
rect 10830 10441 10860 10629
rect 10915 10620 11115 10645
rect 11196 10635 11200 10695
rect 11144 10629 11200 10635
rect 10915 10600 10985 10620
rect 10890 10560 10985 10600
rect 11045 10600 11115 10620
rect 11045 10560 11140 10600
rect 10890 10510 11140 10560
rect 10890 10470 10985 10510
rect 10915 10450 10985 10470
rect 11045 10470 11140 10510
rect 11045 10450 11115 10470
rect 10830 10435 10886 10441
rect 10830 10375 10834 10435
rect 10915 10425 11115 10450
rect 11170 10441 11200 10629
rect 11144 10435 11200 10441
rect 10886 10375 11144 10395
rect 11196 10375 11200 10435
rect 10830 10365 11200 10375
rect 11230 10695 11600 10705
rect 11230 10635 11234 10695
rect 11286 10675 11544 10695
rect 11230 10629 11286 10635
rect 11230 10441 11260 10629
rect 11315 10620 11515 10645
rect 11596 10635 11600 10695
rect 11544 10629 11600 10635
rect 11315 10600 11385 10620
rect 11290 10560 11385 10600
rect 11445 10600 11515 10620
rect 11445 10560 11540 10600
rect 11290 10510 11540 10560
rect 11290 10470 11385 10510
rect 11315 10450 11385 10470
rect 11445 10470 11540 10510
rect 11445 10450 11515 10470
rect 11230 10435 11286 10441
rect 11230 10375 11234 10435
rect 11315 10425 11515 10450
rect 11570 10441 11600 10629
rect 11544 10435 11600 10441
rect 11286 10375 11544 10395
rect 11596 10375 11600 10435
rect 11230 10365 11600 10375
rect 11630 10695 12000 10705
rect 11630 10635 11634 10695
rect 11686 10675 11944 10695
rect 11630 10629 11686 10635
rect 11630 10441 11660 10629
rect 11715 10620 11915 10645
rect 11996 10635 12000 10695
rect 11944 10629 12000 10635
rect 11715 10600 11785 10620
rect 11690 10560 11785 10600
rect 11845 10600 11915 10620
rect 11845 10560 11940 10600
rect 11690 10510 11940 10560
rect 11690 10470 11785 10510
rect 11715 10450 11785 10470
rect 11845 10470 11940 10510
rect 11845 10450 11915 10470
rect 11630 10435 11686 10441
rect 11630 10375 11634 10435
rect 11715 10425 11915 10450
rect 11970 10441 12000 10629
rect 11944 10435 12000 10441
rect 11686 10375 11944 10395
rect 11996 10375 12000 10435
rect 11630 10365 12000 10375
rect 12030 10695 12400 10705
rect 12030 10635 12034 10695
rect 12086 10675 12344 10695
rect 12030 10629 12086 10635
rect 12030 10441 12060 10629
rect 12115 10620 12315 10645
rect 12396 10635 12400 10695
rect 12344 10629 12400 10635
rect 12115 10600 12185 10620
rect 12090 10560 12185 10600
rect 12245 10600 12315 10620
rect 12245 10560 12340 10600
rect 12090 10510 12340 10560
rect 12090 10470 12185 10510
rect 12115 10450 12185 10470
rect 12245 10470 12340 10510
rect 12245 10450 12315 10470
rect 12030 10435 12086 10441
rect 12030 10375 12034 10435
rect 12115 10425 12315 10450
rect 12370 10441 12400 10629
rect 12344 10435 12400 10441
rect 12086 10375 12344 10395
rect 12396 10375 12400 10435
rect 12030 10365 12400 10375
rect 12430 10695 12800 10705
rect 12430 10635 12434 10695
rect 12486 10675 12744 10695
rect 12430 10629 12486 10635
rect 12430 10441 12460 10629
rect 12515 10620 12715 10645
rect 12796 10635 12800 10695
rect 12744 10629 12800 10635
rect 12515 10600 12585 10620
rect 12490 10560 12585 10600
rect 12645 10600 12715 10620
rect 12645 10560 12740 10600
rect 12490 10510 12740 10560
rect 12490 10470 12585 10510
rect 12515 10450 12585 10470
rect 12645 10470 12740 10510
rect 12645 10450 12715 10470
rect 12430 10435 12486 10441
rect 12430 10375 12434 10435
rect 12515 10425 12715 10450
rect 12770 10441 12800 10629
rect 12744 10435 12800 10441
rect 12486 10375 12744 10395
rect 12796 10375 12800 10435
rect 12430 10365 12800 10375
rect 12830 10695 13200 10705
rect 12830 10635 12834 10695
rect 12886 10675 13144 10695
rect 12830 10629 12886 10635
rect 12830 10441 12860 10629
rect 12915 10620 13115 10645
rect 13196 10635 13200 10695
rect 13144 10629 13200 10635
rect 12915 10600 12985 10620
rect 12890 10560 12985 10600
rect 13045 10600 13115 10620
rect 13045 10560 13140 10600
rect 12890 10510 13140 10560
rect 12890 10470 12985 10510
rect 12915 10450 12985 10470
rect 13045 10470 13140 10510
rect 13045 10450 13115 10470
rect 12830 10435 12886 10441
rect 12830 10375 12834 10435
rect 12915 10425 13115 10450
rect 13170 10441 13200 10629
rect 13144 10435 13200 10441
rect 12886 10375 13144 10395
rect 13196 10375 13200 10435
rect 12830 10365 13200 10375
rect -370 10325 0 10335
rect -370 10265 -366 10325
rect -314 10305 -56 10325
rect -370 10259 -314 10265
rect -370 10071 -340 10259
rect -285 10250 -85 10275
rect -4 10265 0 10325
rect -56 10259 0 10265
rect -285 10230 -215 10250
rect -310 10190 -215 10230
rect -155 10230 -85 10250
rect -155 10190 -60 10230
rect -310 10140 -60 10190
rect -310 10100 -215 10140
rect -285 10080 -215 10100
rect -155 10100 -60 10140
rect -155 10080 -85 10100
rect -370 10065 -314 10071
rect -370 10005 -366 10065
rect -285 10055 -85 10080
rect -30 10071 0 10259
rect -56 10065 0 10071
rect -314 10005 -56 10025
rect -4 10005 0 10065
rect -370 9995 0 10005
rect 30 10325 400 10335
rect 30 10265 34 10325
rect 86 10305 344 10325
rect 30 10259 86 10265
rect 30 10071 60 10259
rect 115 10250 315 10275
rect 396 10265 400 10325
rect 344 10259 400 10265
rect 115 10230 185 10250
rect 90 10190 185 10230
rect 245 10230 315 10250
rect 245 10190 340 10230
rect 90 10140 340 10190
rect 90 10100 185 10140
rect 115 10080 185 10100
rect 245 10100 340 10140
rect 245 10080 315 10100
rect 30 10065 86 10071
rect 30 10005 34 10065
rect 115 10055 315 10080
rect 370 10071 400 10259
rect 344 10065 400 10071
rect 86 10005 344 10025
rect 396 10005 400 10065
rect 30 9995 400 10005
rect 430 10325 800 10335
rect 430 10265 434 10325
rect 486 10305 744 10325
rect 430 10259 486 10265
rect 430 10071 460 10259
rect 515 10250 715 10275
rect 796 10265 800 10325
rect 744 10259 800 10265
rect 515 10230 585 10250
rect 490 10190 585 10230
rect 645 10230 715 10250
rect 645 10190 740 10230
rect 490 10140 740 10190
rect 490 10100 585 10140
rect 515 10080 585 10100
rect 645 10100 740 10140
rect 645 10080 715 10100
rect 430 10065 486 10071
rect 430 10005 434 10065
rect 515 10055 715 10080
rect 770 10071 800 10259
rect 744 10065 800 10071
rect 486 10005 744 10025
rect 796 10005 800 10065
rect 430 9995 800 10005
rect 830 10325 1200 10335
rect 830 10265 834 10325
rect 886 10305 1144 10325
rect 830 10259 886 10265
rect 830 10071 860 10259
rect 915 10250 1115 10275
rect 1196 10265 1200 10325
rect 1144 10259 1200 10265
rect 915 10230 985 10250
rect 890 10190 985 10230
rect 1045 10230 1115 10250
rect 1045 10190 1140 10230
rect 890 10140 1140 10190
rect 890 10100 985 10140
rect 915 10080 985 10100
rect 1045 10100 1140 10140
rect 1045 10080 1115 10100
rect 830 10065 886 10071
rect 830 10005 834 10065
rect 915 10055 1115 10080
rect 1170 10071 1200 10259
rect 1144 10065 1200 10071
rect 886 10005 1144 10025
rect 1196 10005 1200 10065
rect 830 9995 1200 10005
rect 1230 10325 1600 10335
rect 1230 10265 1234 10325
rect 1286 10305 1544 10325
rect 1230 10259 1286 10265
rect 1230 10071 1260 10259
rect 1315 10250 1515 10275
rect 1596 10265 1600 10325
rect 1544 10259 1600 10265
rect 1315 10230 1385 10250
rect 1290 10190 1385 10230
rect 1445 10230 1515 10250
rect 1445 10190 1540 10230
rect 1290 10140 1540 10190
rect 1290 10100 1385 10140
rect 1315 10080 1385 10100
rect 1445 10100 1540 10140
rect 1445 10080 1515 10100
rect 1230 10065 1286 10071
rect 1230 10005 1234 10065
rect 1315 10055 1515 10080
rect 1570 10071 1600 10259
rect 1544 10065 1600 10071
rect 1286 10005 1544 10025
rect 1596 10005 1600 10065
rect 1230 9995 1600 10005
rect 1630 10325 2000 10335
rect 1630 10265 1634 10325
rect 1686 10305 1944 10325
rect 1630 10259 1686 10265
rect 1630 10071 1660 10259
rect 1715 10250 1915 10275
rect 1996 10265 2000 10325
rect 1944 10259 2000 10265
rect 1715 10230 1785 10250
rect 1690 10190 1785 10230
rect 1845 10230 1915 10250
rect 1845 10190 1940 10230
rect 1690 10140 1940 10190
rect 1690 10100 1785 10140
rect 1715 10080 1785 10100
rect 1845 10100 1940 10140
rect 1845 10080 1915 10100
rect 1630 10065 1686 10071
rect 1630 10005 1634 10065
rect 1715 10055 1915 10080
rect 1970 10071 2000 10259
rect 1944 10065 2000 10071
rect 1686 10005 1944 10025
rect 1996 10005 2000 10065
rect 1630 9995 2000 10005
rect 2030 10325 2400 10335
rect 2030 10265 2034 10325
rect 2086 10305 2344 10325
rect 2030 10259 2086 10265
rect 2030 10071 2060 10259
rect 2115 10250 2315 10275
rect 2396 10265 2400 10325
rect 2344 10259 2400 10265
rect 2115 10230 2185 10250
rect 2090 10190 2185 10230
rect 2245 10230 2315 10250
rect 2245 10190 2340 10230
rect 2090 10140 2340 10190
rect 2090 10100 2185 10140
rect 2115 10080 2185 10100
rect 2245 10100 2340 10140
rect 2245 10080 2315 10100
rect 2030 10065 2086 10071
rect 2030 10005 2034 10065
rect 2115 10055 2315 10080
rect 2370 10071 2400 10259
rect 2344 10065 2400 10071
rect 2086 10005 2344 10025
rect 2396 10005 2400 10065
rect 2030 9995 2400 10005
rect 2430 10325 2800 10335
rect 2430 10265 2434 10325
rect 2486 10305 2744 10325
rect 2430 10259 2486 10265
rect 2430 10071 2460 10259
rect 2515 10250 2715 10275
rect 2796 10265 2800 10325
rect 2744 10259 2800 10265
rect 2515 10230 2585 10250
rect 2490 10190 2585 10230
rect 2645 10230 2715 10250
rect 2645 10190 2740 10230
rect 2490 10140 2740 10190
rect 2490 10100 2585 10140
rect 2515 10080 2585 10100
rect 2645 10100 2740 10140
rect 2645 10080 2715 10100
rect 2430 10065 2486 10071
rect 2430 10005 2434 10065
rect 2515 10055 2715 10080
rect 2770 10071 2800 10259
rect 2744 10065 2800 10071
rect 2486 10005 2744 10025
rect 2796 10005 2800 10065
rect 2430 9995 2800 10005
rect 2830 10325 3200 10335
rect 2830 10265 2834 10325
rect 2886 10305 3144 10325
rect 2830 10259 2886 10265
rect 2830 10071 2860 10259
rect 2915 10250 3115 10275
rect 3196 10265 3200 10325
rect 3144 10259 3200 10265
rect 2915 10230 2985 10250
rect 2890 10190 2985 10230
rect 3045 10230 3115 10250
rect 3045 10190 3140 10230
rect 2890 10140 3140 10190
rect 2890 10100 2985 10140
rect 2915 10080 2985 10100
rect 3045 10100 3140 10140
rect 3045 10080 3115 10100
rect 2830 10065 2886 10071
rect 2830 10005 2834 10065
rect 2915 10055 3115 10080
rect 3170 10071 3200 10259
rect 3144 10065 3200 10071
rect 2886 10005 3144 10025
rect 3196 10005 3200 10065
rect 2830 9995 3200 10005
rect 3230 10325 3600 10335
rect 3230 10265 3234 10325
rect 3286 10305 3544 10325
rect 3230 10259 3286 10265
rect 3230 10071 3260 10259
rect 3315 10250 3515 10275
rect 3596 10265 3600 10325
rect 3544 10259 3600 10265
rect 3315 10230 3385 10250
rect 3290 10190 3385 10230
rect 3445 10230 3515 10250
rect 3445 10190 3540 10230
rect 3290 10140 3540 10190
rect 3290 10100 3385 10140
rect 3315 10080 3385 10100
rect 3445 10100 3540 10140
rect 3445 10080 3515 10100
rect 3230 10065 3286 10071
rect 3230 10005 3234 10065
rect 3315 10055 3515 10080
rect 3570 10071 3600 10259
rect 3544 10065 3600 10071
rect 3286 10005 3544 10025
rect 3596 10005 3600 10065
rect 3230 9995 3600 10005
rect 3630 10325 4000 10335
rect 3630 10265 3634 10325
rect 3686 10305 3944 10325
rect 3630 10259 3686 10265
rect 3630 10071 3660 10259
rect 3715 10250 3915 10275
rect 3996 10265 4000 10325
rect 3944 10259 4000 10265
rect 3715 10230 3785 10250
rect 3690 10190 3785 10230
rect 3845 10230 3915 10250
rect 3845 10190 3940 10230
rect 3690 10140 3940 10190
rect 3690 10100 3785 10140
rect 3715 10080 3785 10100
rect 3845 10100 3940 10140
rect 3845 10080 3915 10100
rect 3630 10065 3686 10071
rect 3630 10005 3634 10065
rect 3715 10055 3915 10080
rect 3970 10071 4000 10259
rect 3944 10065 4000 10071
rect 3686 10005 3944 10025
rect 3996 10005 4000 10065
rect 3630 9995 4000 10005
rect 4030 10325 4400 10335
rect 4030 10265 4034 10325
rect 4086 10305 4344 10325
rect 4030 10259 4086 10265
rect 4030 10071 4060 10259
rect 4115 10250 4315 10275
rect 4396 10265 4400 10325
rect 4344 10259 4400 10265
rect 4115 10230 4185 10250
rect 4090 10190 4185 10230
rect 4245 10230 4315 10250
rect 4245 10190 4340 10230
rect 4090 10140 4340 10190
rect 4090 10100 4185 10140
rect 4115 10080 4185 10100
rect 4245 10100 4340 10140
rect 4245 10080 4315 10100
rect 4030 10065 4086 10071
rect 4030 10005 4034 10065
rect 4115 10055 4315 10080
rect 4370 10071 4400 10259
rect 4344 10065 4400 10071
rect 4086 10005 4344 10025
rect 4396 10005 4400 10065
rect 4030 9995 4400 10005
rect 4430 10325 4800 10335
rect 4430 10265 4434 10325
rect 4486 10305 4744 10325
rect 4430 10259 4486 10265
rect 4430 10071 4460 10259
rect 4515 10250 4715 10275
rect 4796 10265 4800 10325
rect 4744 10259 4800 10265
rect 4515 10230 4585 10250
rect 4490 10190 4585 10230
rect 4645 10230 4715 10250
rect 4645 10190 4740 10230
rect 4490 10140 4740 10190
rect 4490 10100 4585 10140
rect 4515 10080 4585 10100
rect 4645 10100 4740 10140
rect 4645 10080 4715 10100
rect 4430 10065 4486 10071
rect 4430 10005 4434 10065
rect 4515 10055 4715 10080
rect 4770 10071 4800 10259
rect 4744 10065 4800 10071
rect 4486 10005 4744 10025
rect 4796 10005 4800 10065
rect 4430 9995 4800 10005
rect 4830 10325 5200 10335
rect 4830 10265 4834 10325
rect 4886 10305 5144 10325
rect 4830 10259 4886 10265
rect 4830 10071 4860 10259
rect 4915 10250 5115 10275
rect 5196 10265 5200 10325
rect 5144 10259 5200 10265
rect 4915 10230 4985 10250
rect 4890 10190 4985 10230
rect 5045 10230 5115 10250
rect 5045 10190 5140 10230
rect 4890 10140 5140 10190
rect 4890 10100 4985 10140
rect 4915 10080 4985 10100
rect 5045 10100 5140 10140
rect 5045 10080 5115 10100
rect 4830 10065 4886 10071
rect 4830 10005 4834 10065
rect 4915 10055 5115 10080
rect 5170 10071 5200 10259
rect 5144 10065 5200 10071
rect 4886 10005 5144 10025
rect 5196 10005 5200 10065
rect 4830 9995 5200 10005
rect 5230 10325 5600 10335
rect 5230 10265 5234 10325
rect 5286 10305 5544 10325
rect 5230 10259 5286 10265
rect 5230 10071 5260 10259
rect 5315 10250 5515 10275
rect 5596 10265 5600 10325
rect 5544 10259 5600 10265
rect 5315 10230 5385 10250
rect 5290 10190 5385 10230
rect 5445 10230 5515 10250
rect 5445 10190 5540 10230
rect 5290 10140 5540 10190
rect 5290 10100 5385 10140
rect 5315 10080 5385 10100
rect 5445 10100 5540 10140
rect 5445 10080 5515 10100
rect 5230 10065 5286 10071
rect 5230 10005 5234 10065
rect 5315 10055 5515 10080
rect 5570 10071 5600 10259
rect 5544 10065 5600 10071
rect 5286 10005 5544 10025
rect 5596 10005 5600 10065
rect 5230 9995 5600 10005
rect 5630 10325 6000 10335
rect 5630 10265 5634 10325
rect 5686 10305 5944 10325
rect 5630 10259 5686 10265
rect 5630 10071 5660 10259
rect 5715 10250 5915 10275
rect 5996 10265 6000 10325
rect 5944 10259 6000 10265
rect 5715 10230 5785 10250
rect 5690 10190 5785 10230
rect 5845 10230 5915 10250
rect 5845 10190 5940 10230
rect 5690 10140 5940 10190
rect 5690 10100 5785 10140
rect 5715 10080 5785 10100
rect 5845 10100 5940 10140
rect 5845 10080 5915 10100
rect 5630 10065 5686 10071
rect 5630 10005 5634 10065
rect 5715 10055 5915 10080
rect 5970 10071 6000 10259
rect 5944 10065 6000 10071
rect 5686 10005 5944 10025
rect 5996 10005 6000 10065
rect 5630 9995 6000 10005
rect 6030 10325 6400 10335
rect 6030 10265 6034 10325
rect 6086 10305 6344 10325
rect 6030 10259 6086 10265
rect 6030 10071 6060 10259
rect 6115 10250 6315 10275
rect 6396 10265 6400 10325
rect 6344 10259 6400 10265
rect 6115 10230 6185 10250
rect 6090 10190 6185 10230
rect 6245 10230 6315 10250
rect 6245 10190 6340 10230
rect 6090 10140 6340 10190
rect 6090 10100 6185 10140
rect 6115 10080 6185 10100
rect 6245 10100 6340 10140
rect 6245 10080 6315 10100
rect 6030 10065 6086 10071
rect 6030 10005 6034 10065
rect 6115 10055 6315 10080
rect 6370 10071 6400 10259
rect 6344 10065 6400 10071
rect 6086 10005 6344 10025
rect 6396 10005 6400 10065
rect 6030 9995 6400 10005
rect 6430 10325 6800 10335
rect 6430 10265 6434 10325
rect 6486 10305 6744 10325
rect 6430 10259 6486 10265
rect 6430 10071 6460 10259
rect 6515 10250 6715 10275
rect 6796 10265 6800 10325
rect 6744 10259 6800 10265
rect 6515 10230 6585 10250
rect 6490 10190 6585 10230
rect 6645 10230 6715 10250
rect 6645 10190 6740 10230
rect 6490 10140 6740 10190
rect 6490 10100 6585 10140
rect 6515 10080 6585 10100
rect 6645 10100 6740 10140
rect 6645 10080 6715 10100
rect 6430 10065 6486 10071
rect 6430 10005 6434 10065
rect 6515 10055 6715 10080
rect 6770 10071 6800 10259
rect 6744 10065 6800 10071
rect 6486 10005 6744 10025
rect 6796 10005 6800 10065
rect 6430 9995 6800 10005
rect 6830 10325 7200 10335
rect 6830 10265 6834 10325
rect 6886 10305 7144 10325
rect 6830 10259 6886 10265
rect 6830 10071 6860 10259
rect 6915 10250 7115 10275
rect 7196 10265 7200 10325
rect 7144 10259 7200 10265
rect 6915 10230 6985 10250
rect 6890 10190 6985 10230
rect 7045 10230 7115 10250
rect 7045 10190 7140 10230
rect 6890 10140 7140 10190
rect 6890 10100 6985 10140
rect 6915 10080 6985 10100
rect 7045 10100 7140 10140
rect 7045 10080 7115 10100
rect 6830 10065 6886 10071
rect 6830 10005 6834 10065
rect 6915 10055 7115 10080
rect 7170 10071 7200 10259
rect 7144 10065 7200 10071
rect 6886 10005 7144 10025
rect 7196 10005 7200 10065
rect 6830 9995 7200 10005
rect 7230 10325 7600 10335
rect 7230 10265 7234 10325
rect 7286 10305 7544 10325
rect 7230 10259 7286 10265
rect 7230 10071 7260 10259
rect 7315 10250 7515 10275
rect 7596 10265 7600 10325
rect 7544 10259 7600 10265
rect 7315 10230 7385 10250
rect 7290 10190 7385 10230
rect 7445 10230 7515 10250
rect 7445 10190 7540 10230
rect 7290 10140 7540 10190
rect 7290 10100 7385 10140
rect 7315 10080 7385 10100
rect 7445 10100 7540 10140
rect 7445 10080 7515 10100
rect 7230 10065 7286 10071
rect 7230 10005 7234 10065
rect 7315 10055 7515 10080
rect 7570 10071 7600 10259
rect 7544 10065 7600 10071
rect 7286 10005 7544 10025
rect 7596 10005 7600 10065
rect 7230 9995 7600 10005
rect 7630 10325 8000 10335
rect 7630 10265 7634 10325
rect 7686 10305 7944 10325
rect 7630 10259 7686 10265
rect 7630 10071 7660 10259
rect 7715 10250 7915 10275
rect 7996 10265 8000 10325
rect 7944 10259 8000 10265
rect 7715 10230 7785 10250
rect 7690 10190 7785 10230
rect 7845 10230 7915 10250
rect 7845 10190 7940 10230
rect 7690 10140 7940 10190
rect 7690 10100 7785 10140
rect 7715 10080 7785 10100
rect 7845 10100 7940 10140
rect 7845 10080 7915 10100
rect 7630 10065 7686 10071
rect 7630 10005 7634 10065
rect 7715 10055 7915 10080
rect 7970 10071 8000 10259
rect 7944 10065 8000 10071
rect 7686 10005 7944 10025
rect 7996 10005 8000 10065
rect 7630 9995 8000 10005
rect 8030 10325 8400 10335
rect 8030 10265 8034 10325
rect 8086 10305 8344 10325
rect 8030 10259 8086 10265
rect 8030 10071 8060 10259
rect 8115 10250 8315 10275
rect 8396 10265 8400 10325
rect 8344 10259 8400 10265
rect 8115 10230 8185 10250
rect 8090 10190 8185 10230
rect 8245 10230 8315 10250
rect 8245 10190 8340 10230
rect 8090 10140 8340 10190
rect 8090 10100 8185 10140
rect 8115 10080 8185 10100
rect 8245 10100 8340 10140
rect 8245 10080 8315 10100
rect 8030 10065 8086 10071
rect 8030 10005 8034 10065
rect 8115 10055 8315 10080
rect 8370 10071 8400 10259
rect 8344 10065 8400 10071
rect 8086 10005 8344 10025
rect 8396 10005 8400 10065
rect 8030 9995 8400 10005
rect 8430 10325 8800 10335
rect 8430 10265 8434 10325
rect 8486 10305 8744 10325
rect 8430 10259 8486 10265
rect 8430 10071 8460 10259
rect 8515 10250 8715 10275
rect 8796 10265 8800 10325
rect 8744 10259 8800 10265
rect 8515 10230 8585 10250
rect 8490 10190 8585 10230
rect 8645 10230 8715 10250
rect 8645 10190 8740 10230
rect 8490 10140 8740 10190
rect 8490 10100 8585 10140
rect 8515 10080 8585 10100
rect 8645 10100 8740 10140
rect 8645 10080 8715 10100
rect 8430 10065 8486 10071
rect 8430 10005 8434 10065
rect 8515 10055 8715 10080
rect 8770 10071 8800 10259
rect 8744 10065 8800 10071
rect 8486 10005 8744 10025
rect 8796 10005 8800 10065
rect 8430 9995 8800 10005
rect 8830 10325 9200 10335
rect 8830 10265 8834 10325
rect 8886 10305 9144 10325
rect 8830 10259 8886 10265
rect 8830 10071 8860 10259
rect 8915 10250 9115 10275
rect 9196 10265 9200 10325
rect 9144 10259 9200 10265
rect 8915 10230 8985 10250
rect 8890 10190 8985 10230
rect 9045 10230 9115 10250
rect 9045 10190 9140 10230
rect 8890 10140 9140 10190
rect 8890 10100 8985 10140
rect 8915 10080 8985 10100
rect 9045 10100 9140 10140
rect 9045 10080 9115 10100
rect 8830 10065 8886 10071
rect 8830 10005 8834 10065
rect 8915 10055 9115 10080
rect 9170 10071 9200 10259
rect 9144 10065 9200 10071
rect 8886 10005 9144 10025
rect 9196 10005 9200 10065
rect 8830 9995 9200 10005
rect 9230 10325 9600 10335
rect 9230 10265 9234 10325
rect 9286 10305 9544 10325
rect 9230 10259 9286 10265
rect 9230 10071 9260 10259
rect 9315 10250 9515 10275
rect 9596 10265 9600 10325
rect 9544 10259 9600 10265
rect 9315 10230 9385 10250
rect 9290 10190 9385 10230
rect 9445 10230 9515 10250
rect 9445 10190 9540 10230
rect 9290 10140 9540 10190
rect 9290 10100 9385 10140
rect 9315 10080 9385 10100
rect 9445 10100 9540 10140
rect 9445 10080 9515 10100
rect 9230 10065 9286 10071
rect 9230 10005 9234 10065
rect 9315 10055 9515 10080
rect 9570 10071 9600 10259
rect 9544 10065 9600 10071
rect 9286 10005 9544 10025
rect 9596 10005 9600 10065
rect 9230 9995 9600 10005
rect 9630 10325 10000 10335
rect 9630 10265 9634 10325
rect 9686 10305 9944 10325
rect 9630 10259 9686 10265
rect 9630 10071 9660 10259
rect 9715 10250 9915 10275
rect 9996 10265 10000 10325
rect 9944 10259 10000 10265
rect 9715 10230 9785 10250
rect 9690 10190 9785 10230
rect 9845 10230 9915 10250
rect 9845 10190 9940 10230
rect 9690 10140 9940 10190
rect 9690 10100 9785 10140
rect 9715 10080 9785 10100
rect 9845 10100 9940 10140
rect 9845 10080 9915 10100
rect 9630 10065 9686 10071
rect 9630 10005 9634 10065
rect 9715 10055 9915 10080
rect 9970 10071 10000 10259
rect 9944 10065 10000 10071
rect 9686 10005 9944 10025
rect 9996 10005 10000 10065
rect 9630 9995 10000 10005
rect 10030 10325 10400 10335
rect 10030 10265 10034 10325
rect 10086 10305 10344 10325
rect 10030 10259 10086 10265
rect 10030 10071 10060 10259
rect 10115 10250 10315 10275
rect 10396 10265 10400 10325
rect 10344 10259 10400 10265
rect 10115 10230 10185 10250
rect 10090 10190 10185 10230
rect 10245 10230 10315 10250
rect 10245 10190 10340 10230
rect 10090 10140 10340 10190
rect 10090 10100 10185 10140
rect 10115 10080 10185 10100
rect 10245 10100 10340 10140
rect 10245 10080 10315 10100
rect 10030 10065 10086 10071
rect 10030 10005 10034 10065
rect 10115 10055 10315 10080
rect 10370 10071 10400 10259
rect 10344 10065 10400 10071
rect 10086 10005 10344 10025
rect 10396 10005 10400 10065
rect 10030 9995 10400 10005
rect 10430 10325 10800 10335
rect 10430 10265 10434 10325
rect 10486 10305 10744 10325
rect 10430 10259 10486 10265
rect 10430 10071 10460 10259
rect 10515 10250 10715 10275
rect 10796 10265 10800 10325
rect 10744 10259 10800 10265
rect 10515 10230 10585 10250
rect 10490 10190 10585 10230
rect 10645 10230 10715 10250
rect 10645 10190 10740 10230
rect 10490 10140 10740 10190
rect 10490 10100 10585 10140
rect 10515 10080 10585 10100
rect 10645 10100 10740 10140
rect 10645 10080 10715 10100
rect 10430 10065 10486 10071
rect 10430 10005 10434 10065
rect 10515 10055 10715 10080
rect 10770 10071 10800 10259
rect 10744 10065 10800 10071
rect 10486 10005 10744 10025
rect 10796 10005 10800 10065
rect 10430 9995 10800 10005
rect 10830 10325 11200 10335
rect 10830 10265 10834 10325
rect 10886 10305 11144 10325
rect 10830 10259 10886 10265
rect 10830 10071 10860 10259
rect 10915 10250 11115 10275
rect 11196 10265 11200 10325
rect 11144 10259 11200 10265
rect 10915 10230 10985 10250
rect 10890 10190 10985 10230
rect 11045 10230 11115 10250
rect 11045 10190 11140 10230
rect 10890 10140 11140 10190
rect 10890 10100 10985 10140
rect 10915 10080 10985 10100
rect 11045 10100 11140 10140
rect 11045 10080 11115 10100
rect 10830 10065 10886 10071
rect 10830 10005 10834 10065
rect 10915 10055 11115 10080
rect 11170 10071 11200 10259
rect 11144 10065 11200 10071
rect 10886 10005 11144 10025
rect 11196 10005 11200 10065
rect 10830 9995 11200 10005
rect 11230 10325 11600 10335
rect 11230 10265 11234 10325
rect 11286 10305 11544 10325
rect 11230 10259 11286 10265
rect 11230 10071 11260 10259
rect 11315 10250 11515 10275
rect 11596 10265 11600 10325
rect 11544 10259 11600 10265
rect 11315 10230 11385 10250
rect 11290 10190 11385 10230
rect 11445 10230 11515 10250
rect 11445 10190 11540 10230
rect 11290 10140 11540 10190
rect 11290 10100 11385 10140
rect 11315 10080 11385 10100
rect 11445 10100 11540 10140
rect 11445 10080 11515 10100
rect 11230 10065 11286 10071
rect 11230 10005 11234 10065
rect 11315 10055 11515 10080
rect 11570 10071 11600 10259
rect 11544 10065 11600 10071
rect 11286 10005 11544 10025
rect 11596 10005 11600 10065
rect 11230 9995 11600 10005
rect 11630 10325 12000 10335
rect 11630 10265 11634 10325
rect 11686 10305 11944 10325
rect 11630 10259 11686 10265
rect 11630 10071 11660 10259
rect 11715 10250 11915 10275
rect 11996 10265 12000 10325
rect 11944 10259 12000 10265
rect 11715 10230 11785 10250
rect 11690 10190 11785 10230
rect 11845 10230 11915 10250
rect 11845 10190 11940 10230
rect 11690 10140 11940 10190
rect 11690 10100 11785 10140
rect 11715 10080 11785 10100
rect 11845 10100 11940 10140
rect 11845 10080 11915 10100
rect 11630 10065 11686 10071
rect 11630 10005 11634 10065
rect 11715 10055 11915 10080
rect 11970 10071 12000 10259
rect 11944 10065 12000 10071
rect 11686 10005 11944 10025
rect 11996 10005 12000 10065
rect 11630 9995 12000 10005
rect 12030 10325 12400 10335
rect 12030 10265 12034 10325
rect 12086 10305 12344 10325
rect 12030 10259 12086 10265
rect 12030 10071 12060 10259
rect 12115 10250 12315 10275
rect 12396 10265 12400 10325
rect 12344 10259 12400 10265
rect 12115 10230 12185 10250
rect 12090 10190 12185 10230
rect 12245 10230 12315 10250
rect 12245 10190 12340 10230
rect 12090 10140 12340 10190
rect 12090 10100 12185 10140
rect 12115 10080 12185 10100
rect 12245 10100 12340 10140
rect 12245 10080 12315 10100
rect 12030 10065 12086 10071
rect 12030 10005 12034 10065
rect 12115 10055 12315 10080
rect 12370 10071 12400 10259
rect 12344 10065 12400 10071
rect 12086 10005 12344 10025
rect 12396 10005 12400 10065
rect 12030 9995 12400 10005
rect 12430 10325 12800 10335
rect 12430 10265 12434 10325
rect 12486 10305 12744 10325
rect 12430 10259 12486 10265
rect 12430 10071 12460 10259
rect 12515 10250 12715 10275
rect 12796 10265 12800 10325
rect 12744 10259 12800 10265
rect 12515 10230 12585 10250
rect 12490 10190 12585 10230
rect 12645 10230 12715 10250
rect 12645 10190 12740 10230
rect 12490 10140 12740 10190
rect 12490 10100 12585 10140
rect 12515 10080 12585 10100
rect 12645 10100 12740 10140
rect 12645 10080 12715 10100
rect 12430 10065 12486 10071
rect 12430 10005 12434 10065
rect 12515 10055 12715 10080
rect 12770 10071 12800 10259
rect 12744 10065 12800 10071
rect 12486 10005 12744 10025
rect 12796 10005 12800 10065
rect 12430 9995 12800 10005
rect 12830 10325 13200 10335
rect 12830 10265 12834 10325
rect 12886 10305 13144 10325
rect 12830 10259 12886 10265
rect 12830 10071 12860 10259
rect 12915 10250 13115 10275
rect 13196 10265 13200 10325
rect 13144 10259 13200 10265
rect 12915 10230 12985 10250
rect 12890 10190 12985 10230
rect 13045 10230 13115 10250
rect 13045 10190 13140 10230
rect 12890 10140 13140 10190
rect 12890 10100 12985 10140
rect 12915 10080 12985 10100
rect 13045 10100 13140 10140
rect 13045 10080 13115 10100
rect 12830 10065 12886 10071
rect 12830 10005 12834 10065
rect 12915 10055 13115 10080
rect 13170 10071 13200 10259
rect 13144 10065 13200 10071
rect 12886 10005 13144 10025
rect 13196 10005 13200 10065
rect 12830 9995 13200 10005
rect -370 9955 0 9965
rect -370 9895 -366 9955
rect -314 9935 -56 9955
rect -370 9889 -314 9895
rect -370 9701 -340 9889
rect -285 9880 -85 9905
rect -4 9895 0 9955
rect -56 9889 0 9895
rect -285 9860 -215 9880
rect -310 9820 -215 9860
rect -155 9860 -85 9880
rect -155 9820 -60 9860
rect -310 9770 -60 9820
rect -310 9730 -215 9770
rect -285 9710 -215 9730
rect -155 9730 -60 9770
rect -155 9710 -85 9730
rect -370 9695 -314 9701
rect -370 9635 -366 9695
rect -285 9685 -85 9710
rect -30 9701 0 9889
rect -56 9695 0 9701
rect -314 9635 -56 9655
rect -4 9635 0 9695
rect -370 9625 0 9635
rect 30 9955 400 9965
rect 30 9895 34 9955
rect 86 9935 344 9955
rect 30 9889 86 9895
rect 30 9701 60 9889
rect 115 9880 315 9905
rect 396 9895 400 9955
rect 344 9889 400 9895
rect 115 9860 185 9880
rect 90 9820 185 9860
rect 245 9860 315 9880
rect 245 9820 340 9860
rect 90 9770 340 9820
rect 90 9730 185 9770
rect 115 9710 185 9730
rect 245 9730 340 9770
rect 245 9710 315 9730
rect 30 9695 86 9701
rect 30 9635 34 9695
rect 115 9685 315 9710
rect 370 9701 400 9889
rect 344 9695 400 9701
rect 86 9635 344 9655
rect 396 9635 400 9695
rect 30 9625 400 9635
rect 430 9955 800 9965
rect 430 9895 434 9955
rect 486 9935 744 9955
rect 430 9889 486 9895
rect 430 9701 460 9889
rect 515 9880 715 9905
rect 796 9895 800 9955
rect 744 9889 800 9895
rect 515 9860 585 9880
rect 490 9820 585 9860
rect 645 9860 715 9880
rect 645 9820 740 9860
rect 490 9770 740 9820
rect 490 9730 585 9770
rect 515 9710 585 9730
rect 645 9730 740 9770
rect 645 9710 715 9730
rect 430 9695 486 9701
rect 430 9635 434 9695
rect 515 9685 715 9710
rect 770 9701 800 9889
rect 744 9695 800 9701
rect 486 9635 744 9655
rect 796 9635 800 9695
rect 430 9625 800 9635
rect 830 9955 1200 9965
rect 830 9895 834 9955
rect 886 9935 1144 9955
rect 830 9889 886 9895
rect 830 9701 860 9889
rect 915 9880 1115 9905
rect 1196 9895 1200 9955
rect 1144 9889 1200 9895
rect 915 9860 985 9880
rect 890 9820 985 9860
rect 1045 9860 1115 9880
rect 1045 9820 1140 9860
rect 890 9770 1140 9820
rect 890 9730 985 9770
rect 915 9710 985 9730
rect 1045 9730 1140 9770
rect 1045 9710 1115 9730
rect 830 9695 886 9701
rect 830 9635 834 9695
rect 915 9685 1115 9710
rect 1170 9701 1200 9889
rect 1144 9695 1200 9701
rect 886 9635 1144 9655
rect 1196 9635 1200 9695
rect 830 9625 1200 9635
rect 1230 9955 1600 9965
rect 1230 9895 1234 9955
rect 1286 9935 1544 9955
rect 1230 9889 1286 9895
rect 1230 9701 1260 9889
rect 1315 9880 1515 9905
rect 1596 9895 1600 9955
rect 1544 9889 1600 9895
rect 1315 9860 1385 9880
rect 1290 9820 1385 9860
rect 1445 9860 1515 9880
rect 1445 9820 1540 9860
rect 1290 9770 1540 9820
rect 1290 9730 1385 9770
rect 1315 9710 1385 9730
rect 1445 9730 1540 9770
rect 1445 9710 1515 9730
rect 1230 9695 1286 9701
rect 1230 9635 1234 9695
rect 1315 9685 1515 9710
rect 1570 9701 1600 9889
rect 1544 9695 1600 9701
rect 1286 9635 1544 9655
rect 1596 9635 1600 9695
rect 1230 9625 1600 9635
rect 1630 9955 2000 9965
rect 1630 9895 1634 9955
rect 1686 9935 1944 9955
rect 1630 9889 1686 9895
rect 1630 9701 1660 9889
rect 1715 9880 1915 9905
rect 1996 9895 2000 9955
rect 1944 9889 2000 9895
rect 1715 9860 1785 9880
rect 1690 9820 1785 9860
rect 1845 9860 1915 9880
rect 1845 9820 1940 9860
rect 1690 9770 1940 9820
rect 1690 9730 1785 9770
rect 1715 9710 1785 9730
rect 1845 9730 1940 9770
rect 1845 9710 1915 9730
rect 1630 9695 1686 9701
rect 1630 9635 1634 9695
rect 1715 9685 1915 9710
rect 1970 9701 2000 9889
rect 1944 9695 2000 9701
rect 1686 9635 1944 9655
rect 1996 9635 2000 9695
rect 1630 9625 2000 9635
rect 2030 9955 2400 9965
rect 2030 9895 2034 9955
rect 2086 9935 2344 9955
rect 2030 9889 2086 9895
rect 2030 9701 2060 9889
rect 2115 9880 2315 9905
rect 2396 9895 2400 9955
rect 2344 9889 2400 9895
rect 2115 9860 2185 9880
rect 2090 9820 2185 9860
rect 2245 9860 2315 9880
rect 2245 9820 2340 9860
rect 2090 9770 2340 9820
rect 2090 9730 2185 9770
rect 2115 9710 2185 9730
rect 2245 9730 2340 9770
rect 2245 9710 2315 9730
rect 2030 9695 2086 9701
rect 2030 9635 2034 9695
rect 2115 9685 2315 9710
rect 2370 9701 2400 9889
rect 2344 9695 2400 9701
rect 2086 9635 2344 9655
rect 2396 9635 2400 9695
rect 2030 9625 2400 9635
rect 2430 9955 2800 9965
rect 2430 9895 2434 9955
rect 2486 9935 2744 9955
rect 2430 9889 2486 9895
rect 2430 9701 2460 9889
rect 2515 9880 2715 9905
rect 2796 9895 2800 9955
rect 2744 9889 2800 9895
rect 2515 9860 2585 9880
rect 2490 9820 2585 9860
rect 2645 9860 2715 9880
rect 2645 9820 2740 9860
rect 2490 9770 2740 9820
rect 2490 9730 2585 9770
rect 2515 9710 2585 9730
rect 2645 9730 2740 9770
rect 2645 9710 2715 9730
rect 2430 9695 2486 9701
rect 2430 9635 2434 9695
rect 2515 9685 2715 9710
rect 2770 9701 2800 9889
rect 2744 9695 2800 9701
rect 2486 9635 2744 9655
rect 2796 9635 2800 9695
rect 2430 9625 2800 9635
rect 2830 9955 3200 9965
rect 2830 9895 2834 9955
rect 2886 9935 3144 9955
rect 2830 9889 2886 9895
rect 2830 9701 2860 9889
rect 2915 9880 3115 9905
rect 3196 9895 3200 9955
rect 3144 9889 3200 9895
rect 2915 9860 2985 9880
rect 2890 9820 2985 9860
rect 3045 9860 3115 9880
rect 3045 9820 3140 9860
rect 2890 9770 3140 9820
rect 2890 9730 2985 9770
rect 2915 9710 2985 9730
rect 3045 9730 3140 9770
rect 3045 9710 3115 9730
rect 2830 9695 2886 9701
rect 2830 9635 2834 9695
rect 2915 9685 3115 9710
rect 3170 9701 3200 9889
rect 3144 9695 3200 9701
rect 2886 9635 3144 9655
rect 3196 9635 3200 9695
rect 2830 9625 3200 9635
rect 3230 9955 3600 9965
rect 3230 9895 3234 9955
rect 3286 9935 3544 9955
rect 3230 9889 3286 9895
rect 3230 9701 3260 9889
rect 3315 9880 3515 9905
rect 3596 9895 3600 9955
rect 3544 9889 3600 9895
rect 3315 9860 3385 9880
rect 3290 9820 3385 9860
rect 3445 9860 3515 9880
rect 3445 9820 3540 9860
rect 3290 9770 3540 9820
rect 3290 9730 3385 9770
rect 3315 9710 3385 9730
rect 3445 9730 3540 9770
rect 3445 9710 3515 9730
rect 3230 9695 3286 9701
rect 3230 9635 3234 9695
rect 3315 9685 3515 9710
rect 3570 9701 3600 9889
rect 3544 9695 3600 9701
rect 3286 9635 3544 9655
rect 3596 9635 3600 9695
rect 3230 9625 3600 9635
rect 3630 9955 4000 9965
rect 3630 9895 3634 9955
rect 3686 9935 3944 9955
rect 3630 9889 3686 9895
rect 3630 9701 3660 9889
rect 3715 9880 3915 9905
rect 3996 9895 4000 9955
rect 3944 9889 4000 9895
rect 3715 9860 3785 9880
rect 3690 9820 3785 9860
rect 3845 9860 3915 9880
rect 3845 9820 3940 9860
rect 3690 9770 3940 9820
rect 3690 9730 3785 9770
rect 3715 9710 3785 9730
rect 3845 9730 3940 9770
rect 3845 9710 3915 9730
rect 3630 9695 3686 9701
rect 3630 9635 3634 9695
rect 3715 9685 3915 9710
rect 3970 9701 4000 9889
rect 3944 9695 4000 9701
rect 3686 9635 3944 9655
rect 3996 9635 4000 9695
rect 3630 9625 4000 9635
rect 4030 9955 4400 9965
rect 4030 9895 4034 9955
rect 4086 9935 4344 9955
rect 4030 9889 4086 9895
rect 4030 9701 4060 9889
rect 4115 9880 4315 9905
rect 4396 9895 4400 9955
rect 4344 9889 4400 9895
rect 4115 9860 4185 9880
rect 4090 9820 4185 9860
rect 4245 9860 4315 9880
rect 4245 9820 4340 9860
rect 4090 9770 4340 9820
rect 4090 9730 4185 9770
rect 4115 9710 4185 9730
rect 4245 9730 4340 9770
rect 4245 9710 4315 9730
rect 4030 9695 4086 9701
rect 4030 9635 4034 9695
rect 4115 9685 4315 9710
rect 4370 9701 4400 9889
rect 4344 9695 4400 9701
rect 4086 9635 4344 9655
rect 4396 9635 4400 9695
rect 4030 9625 4400 9635
rect 4430 9955 4800 9965
rect 4430 9895 4434 9955
rect 4486 9935 4744 9955
rect 4430 9889 4486 9895
rect 4430 9701 4460 9889
rect 4515 9880 4715 9905
rect 4796 9895 4800 9955
rect 4744 9889 4800 9895
rect 4515 9860 4585 9880
rect 4490 9820 4585 9860
rect 4645 9860 4715 9880
rect 4645 9820 4740 9860
rect 4490 9770 4740 9820
rect 4490 9730 4585 9770
rect 4515 9710 4585 9730
rect 4645 9730 4740 9770
rect 4645 9710 4715 9730
rect 4430 9695 4486 9701
rect 4430 9635 4434 9695
rect 4515 9685 4715 9710
rect 4770 9701 4800 9889
rect 4744 9695 4800 9701
rect 4486 9635 4744 9655
rect 4796 9635 4800 9695
rect 4430 9625 4800 9635
rect 4830 9955 5200 9965
rect 4830 9895 4834 9955
rect 4886 9935 5144 9955
rect 4830 9889 4886 9895
rect 4830 9701 4860 9889
rect 4915 9880 5115 9905
rect 5196 9895 5200 9955
rect 5144 9889 5200 9895
rect 4915 9860 4985 9880
rect 4890 9820 4985 9860
rect 5045 9860 5115 9880
rect 5045 9820 5140 9860
rect 4890 9770 5140 9820
rect 4890 9730 4985 9770
rect 4915 9710 4985 9730
rect 5045 9730 5140 9770
rect 5045 9710 5115 9730
rect 4830 9695 4886 9701
rect 4830 9635 4834 9695
rect 4915 9685 5115 9710
rect 5170 9701 5200 9889
rect 5144 9695 5200 9701
rect 4886 9635 5144 9655
rect 5196 9635 5200 9695
rect 4830 9625 5200 9635
rect 5230 9955 5600 9965
rect 5230 9895 5234 9955
rect 5286 9935 5544 9955
rect 5230 9889 5286 9895
rect 5230 9701 5260 9889
rect 5315 9880 5515 9905
rect 5596 9895 5600 9955
rect 5544 9889 5600 9895
rect 5315 9860 5385 9880
rect 5290 9820 5385 9860
rect 5445 9860 5515 9880
rect 5445 9820 5540 9860
rect 5290 9770 5540 9820
rect 5290 9730 5385 9770
rect 5315 9710 5385 9730
rect 5445 9730 5540 9770
rect 5445 9710 5515 9730
rect 5230 9695 5286 9701
rect 5230 9635 5234 9695
rect 5315 9685 5515 9710
rect 5570 9701 5600 9889
rect 5544 9695 5600 9701
rect 5286 9635 5544 9655
rect 5596 9635 5600 9695
rect 5230 9625 5600 9635
rect 5630 9955 6000 9965
rect 5630 9895 5634 9955
rect 5686 9935 5944 9955
rect 5630 9889 5686 9895
rect 5630 9701 5660 9889
rect 5715 9880 5915 9905
rect 5996 9895 6000 9955
rect 5944 9889 6000 9895
rect 5715 9860 5785 9880
rect 5690 9820 5785 9860
rect 5845 9860 5915 9880
rect 5845 9820 5940 9860
rect 5690 9770 5940 9820
rect 5690 9730 5785 9770
rect 5715 9710 5785 9730
rect 5845 9730 5940 9770
rect 5845 9710 5915 9730
rect 5630 9695 5686 9701
rect 5630 9635 5634 9695
rect 5715 9685 5915 9710
rect 5970 9701 6000 9889
rect 5944 9695 6000 9701
rect 5686 9635 5944 9655
rect 5996 9635 6000 9695
rect 5630 9625 6000 9635
rect 6030 9955 6400 9965
rect 6030 9895 6034 9955
rect 6086 9935 6344 9955
rect 6030 9889 6086 9895
rect 6030 9701 6060 9889
rect 6115 9880 6315 9905
rect 6396 9895 6400 9955
rect 6344 9889 6400 9895
rect 6115 9860 6185 9880
rect 6090 9820 6185 9860
rect 6245 9860 6315 9880
rect 6245 9820 6340 9860
rect 6090 9770 6340 9820
rect 6090 9730 6185 9770
rect 6115 9710 6185 9730
rect 6245 9730 6340 9770
rect 6245 9710 6315 9730
rect 6030 9695 6086 9701
rect 6030 9635 6034 9695
rect 6115 9685 6315 9710
rect 6370 9701 6400 9889
rect 6344 9695 6400 9701
rect 6086 9635 6344 9655
rect 6396 9635 6400 9695
rect 6030 9625 6400 9635
rect 6430 9955 6800 9965
rect 6430 9895 6434 9955
rect 6486 9935 6744 9955
rect 6430 9889 6486 9895
rect 6430 9701 6460 9889
rect 6515 9880 6715 9905
rect 6796 9895 6800 9955
rect 6744 9889 6800 9895
rect 6515 9860 6585 9880
rect 6490 9820 6585 9860
rect 6645 9860 6715 9880
rect 6645 9820 6740 9860
rect 6490 9770 6740 9820
rect 6490 9730 6585 9770
rect 6515 9710 6585 9730
rect 6645 9730 6740 9770
rect 6645 9710 6715 9730
rect 6430 9695 6486 9701
rect 6430 9635 6434 9695
rect 6515 9685 6715 9710
rect 6770 9701 6800 9889
rect 6744 9695 6800 9701
rect 6486 9635 6744 9655
rect 6796 9635 6800 9695
rect 6430 9625 6800 9635
rect 6830 9955 7200 9965
rect 6830 9895 6834 9955
rect 6886 9935 7144 9955
rect 6830 9889 6886 9895
rect 6830 9701 6860 9889
rect 6915 9880 7115 9905
rect 7196 9895 7200 9955
rect 7144 9889 7200 9895
rect 6915 9860 6985 9880
rect 6890 9820 6985 9860
rect 7045 9860 7115 9880
rect 7045 9820 7140 9860
rect 6890 9770 7140 9820
rect 6890 9730 6985 9770
rect 6915 9710 6985 9730
rect 7045 9730 7140 9770
rect 7045 9710 7115 9730
rect 6830 9695 6886 9701
rect 6830 9635 6834 9695
rect 6915 9685 7115 9710
rect 7170 9701 7200 9889
rect 7144 9695 7200 9701
rect 6886 9635 7144 9655
rect 7196 9635 7200 9695
rect 6830 9625 7200 9635
rect 7230 9955 7600 9965
rect 7230 9895 7234 9955
rect 7286 9935 7544 9955
rect 7230 9889 7286 9895
rect 7230 9701 7260 9889
rect 7315 9880 7515 9905
rect 7596 9895 7600 9955
rect 7544 9889 7600 9895
rect 7315 9860 7385 9880
rect 7290 9820 7385 9860
rect 7445 9860 7515 9880
rect 7445 9820 7540 9860
rect 7290 9770 7540 9820
rect 7290 9730 7385 9770
rect 7315 9710 7385 9730
rect 7445 9730 7540 9770
rect 7445 9710 7515 9730
rect 7230 9695 7286 9701
rect 7230 9635 7234 9695
rect 7315 9685 7515 9710
rect 7570 9701 7600 9889
rect 7544 9695 7600 9701
rect 7286 9635 7544 9655
rect 7596 9635 7600 9695
rect 7230 9625 7600 9635
rect 7630 9955 8000 9965
rect 7630 9895 7634 9955
rect 7686 9935 7944 9955
rect 7630 9889 7686 9895
rect 7630 9701 7660 9889
rect 7715 9880 7915 9905
rect 7996 9895 8000 9955
rect 7944 9889 8000 9895
rect 7715 9860 7785 9880
rect 7690 9820 7785 9860
rect 7845 9860 7915 9880
rect 7845 9820 7940 9860
rect 7690 9770 7940 9820
rect 7690 9730 7785 9770
rect 7715 9710 7785 9730
rect 7845 9730 7940 9770
rect 7845 9710 7915 9730
rect 7630 9695 7686 9701
rect 7630 9635 7634 9695
rect 7715 9685 7915 9710
rect 7970 9701 8000 9889
rect 7944 9695 8000 9701
rect 7686 9635 7944 9655
rect 7996 9635 8000 9695
rect 7630 9625 8000 9635
rect 8030 9955 8400 9965
rect 8030 9895 8034 9955
rect 8086 9935 8344 9955
rect 8030 9889 8086 9895
rect 8030 9701 8060 9889
rect 8115 9880 8315 9905
rect 8396 9895 8400 9955
rect 8344 9889 8400 9895
rect 8115 9860 8185 9880
rect 8090 9820 8185 9860
rect 8245 9860 8315 9880
rect 8245 9820 8340 9860
rect 8090 9770 8340 9820
rect 8090 9730 8185 9770
rect 8115 9710 8185 9730
rect 8245 9730 8340 9770
rect 8245 9710 8315 9730
rect 8030 9695 8086 9701
rect 8030 9635 8034 9695
rect 8115 9685 8315 9710
rect 8370 9701 8400 9889
rect 8344 9695 8400 9701
rect 8086 9635 8344 9655
rect 8396 9635 8400 9695
rect 8030 9625 8400 9635
rect 8430 9955 8800 9965
rect 8430 9895 8434 9955
rect 8486 9935 8744 9955
rect 8430 9889 8486 9895
rect 8430 9701 8460 9889
rect 8515 9880 8715 9905
rect 8796 9895 8800 9955
rect 8744 9889 8800 9895
rect 8515 9860 8585 9880
rect 8490 9820 8585 9860
rect 8645 9860 8715 9880
rect 8645 9820 8740 9860
rect 8490 9770 8740 9820
rect 8490 9730 8585 9770
rect 8515 9710 8585 9730
rect 8645 9730 8740 9770
rect 8645 9710 8715 9730
rect 8430 9695 8486 9701
rect 8430 9635 8434 9695
rect 8515 9685 8715 9710
rect 8770 9701 8800 9889
rect 8744 9695 8800 9701
rect 8486 9635 8744 9655
rect 8796 9635 8800 9695
rect 8430 9625 8800 9635
rect 8830 9955 9200 9965
rect 8830 9895 8834 9955
rect 8886 9935 9144 9955
rect 8830 9889 8886 9895
rect 8830 9701 8860 9889
rect 8915 9880 9115 9905
rect 9196 9895 9200 9955
rect 9144 9889 9200 9895
rect 8915 9860 8985 9880
rect 8890 9820 8985 9860
rect 9045 9860 9115 9880
rect 9045 9820 9140 9860
rect 8890 9770 9140 9820
rect 8890 9730 8985 9770
rect 8915 9710 8985 9730
rect 9045 9730 9140 9770
rect 9045 9710 9115 9730
rect 8830 9695 8886 9701
rect 8830 9635 8834 9695
rect 8915 9685 9115 9710
rect 9170 9701 9200 9889
rect 9144 9695 9200 9701
rect 8886 9635 9144 9655
rect 9196 9635 9200 9695
rect 8830 9625 9200 9635
rect 9230 9955 9600 9965
rect 9230 9895 9234 9955
rect 9286 9935 9544 9955
rect 9230 9889 9286 9895
rect 9230 9701 9260 9889
rect 9315 9880 9515 9905
rect 9596 9895 9600 9955
rect 9544 9889 9600 9895
rect 9315 9860 9385 9880
rect 9290 9820 9385 9860
rect 9445 9860 9515 9880
rect 9445 9820 9540 9860
rect 9290 9770 9540 9820
rect 9290 9730 9385 9770
rect 9315 9710 9385 9730
rect 9445 9730 9540 9770
rect 9445 9710 9515 9730
rect 9230 9695 9286 9701
rect 9230 9635 9234 9695
rect 9315 9685 9515 9710
rect 9570 9701 9600 9889
rect 9544 9695 9600 9701
rect 9286 9635 9544 9655
rect 9596 9635 9600 9695
rect 9230 9625 9600 9635
rect 9630 9955 10000 9965
rect 9630 9895 9634 9955
rect 9686 9935 9944 9955
rect 9630 9889 9686 9895
rect 9630 9701 9660 9889
rect 9715 9880 9915 9905
rect 9996 9895 10000 9955
rect 9944 9889 10000 9895
rect 9715 9860 9785 9880
rect 9690 9820 9785 9860
rect 9845 9860 9915 9880
rect 9845 9820 9940 9860
rect 9690 9770 9940 9820
rect 9690 9730 9785 9770
rect 9715 9710 9785 9730
rect 9845 9730 9940 9770
rect 9845 9710 9915 9730
rect 9630 9695 9686 9701
rect 9630 9635 9634 9695
rect 9715 9685 9915 9710
rect 9970 9701 10000 9889
rect 9944 9695 10000 9701
rect 9686 9635 9944 9655
rect 9996 9635 10000 9695
rect 9630 9625 10000 9635
rect 10030 9955 10400 9965
rect 10030 9895 10034 9955
rect 10086 9935 10344 9955
rect 10030 9889 10086 9895
rect 10030 9701 10060 9889
rect 10115 9880 10315 9905
rect 10396 9895 10400 9955
rect 10344 9889 10400 9895
rect 10115 9860 10185 9880
rect 10090 9820 10185 9860
rect 10245 9860 10315 9880
rect 10245 9820 10340 9860
rect 10090 9770 10340 9820
rect 10090 9730 10185 9770
rect 10115 9710 10185 9730
rect 10245 9730 10340 9770
rect 10245 9710 10315 9730
rect 10030 9695 10086 9701
rect 10030 9635 10034 9695
rect 10115 9685 10315 9710
rect 10370 9701 10400 9889
rect 10344 9695 10400 9701
rect 10086 9635 10344 9655
rect 10396 9635 10400 9695
rect 10030 9625 10400 9635
rect 10430 9955 10800 9965
rect 10430 9895 10434 9955
rect 10486 9935 10744 9955
rect 10430 9889 10486 9895
rect 10430 9701 10460 9889
rect 10515 9880 10715 9905
rect 10796 9895 10800 9955
rect 10744 9889 10800 9895
rect 10515 9860 10585 9880
rect 10490 9820 10585 9860
rect 10645 9860 10715 9880
rect 10645 9820 10740 9860
rect 10490 9770 10740 9820
rect 10490 9730 10585 9770
rect 10515 9710 10585 9730
rect 10645 9730 10740 9770
rect 10645 9710 10715 9730
rect 10430 9695 10486 9701
rect 10430 9635 10434 9695
rect 10515 9685 10715 9710
rect 10770 9701 10800 9889
rect 10744 9695 10800 9701
rect 10486 9635 10744 9655
rect 10796 9635 10800 9695
rect 10430 9625 10800 9635
rect 10830 9955 11200 9965
rect 10830 9895 10834 9955
rect 10886 9935 11144 9955
rect 10830 9889 10886 9895
rect 10830 9701 10860 9889
rect 10915 9880 11115 9905
rect 11196 9895 11200 9955
rect 11144 9889 11200 9895
rect 10915 9860 10985 9880
rect 10890 9820 10985 9860
rect 11045 9860 11115 9880
rect 11045 9820 11140 9860
rect 10890 9770 11140 9820
rect 10890 9730 10985 9770
rect 10915 9710 10985 9730
rect 11045 9730 11140 9770
rect 11045 9710 11115 9730
rect 10830 9695 10886 9701
rect 10830 9635 10834 9695
rect 10915 9685 11115 9710
rect 11170 9701 11200 9889
rect 11144 9695 11200 9701
rect 10886 9635 11144 9655
rect 11196 9635 11200 9695
rect 10830 9625 11200 9635
rect 11230 9955 11600 9965
rect 11230 9895 11234 9955
rect 11286 9935 11544 9955
rect 11230 9889 11286 9895
rect 11230 9701 11260 9889
rect 11315 9880 11515 9905
rect 11596 9895 11600 9955
rect 11544 9889 11600 9895
rect 11315 9860 11385 9880
rect 11290 9820 11385 9860
rect 11445 9860 11515 9880
rect 11445 9820 11540 9860
rect 11290 9770 11540 9820
rect 11290 9730 11385 9770
rect 11315 9710 11385 9730
rect 11445 9730 11540 9770
rect 11445 9710 11515 9730
rect 11230 9695 11286 9701
rect 11230 9635 11234 9695
rect 11315 9685 11515 9710
rect 11570 9701 11600 9889
rect 11544 9695 11600 9701
rect 11286 9635 11544 9655
rect 11596 9635 11600 9695
rect 11230 9625 11600 9635
rect 11630 9955 12000 9965
rect 11630 9895 11634 9955
rect 11686 9935 11944 9955
rect 11630 9889 11686 9895
rect 11630 9701 11660 9889
rect 11715 9880 11915 9905
rect 11996 9895 12000 9955
rect 11944 9889 12000 9895
rect 11715 9860 11785 9880
rect 11690 9820 11785 9860
rect 11845 9860 11915 9880
rect 11845 9820 11940 9860
rect 11690 9770 11940 9820
rect 11690 9730 11785 9770
rect 11715 9710 11785 9730
rect 11845 9730 11940 9770
rect 11845 9710 11915 9730
rect 11630 9695 11686 9701
rect 11630 9635 11634 9695
rect 11715 9685 11915 9710
rect 11970 9701 12000 9889
rect 11944 9695 12000 9701
rect 11686 9635 11944 9655
rect 11996 9635 12000 9695
rect 11630 9625 12000 9635
rect 12030 9955 12400 9965
rect 12030 9895 12034 9955
rect 12086 9935 12344 9955
rect 12030 9889 12086 9895
rect 12030 9701 12060 9889
rect 12115 9880 12315 9905
rect 12396 9895 12400 9955
rect 12344 9889 12400 9895
rect 12115 9860 12185 9880
rect 12090 9820 12185 9860
rect 12245 9860 12315 9880
rect 12245 9820 12340 9860
rect 12090 9770 12340 9820
rect 12090 9730 12185 9770
rect 12115 9710 12185 9730
rect 12245 9730 12340 9770
rect 12245 9710 12315 9730
rect 12030 9695 12086 9701
rect 12030 9635 12034 9695
rect 12115 9685 12315 9710
rect 12370 9701 12400 9889
rect 12344 9695 12400 9701
rect 12086 9635 12344 9655
rect 12396 9635 12400 9695
rect 12030 9625 12400 9635
rect 12430 9955 12800 9965
rect 12430 9895 12434 9955
rect 12486 9935 12744 9955
rect 12430 9889 12486 9895
rect 12430 9701 12460 9889
rect 12515 9880 12715 9905
rect 12796 9895 12800 9955
rect 12744 9889 12800 9895
rect 12515 9860 12585 9880
rect 12490 9820 12585 9860
rect 12645 9860 12715 9880
rect 12645 9820 12740 9860
rect 12490 9770 12740 9820
rect 12490 9730 12585 9770
rect 12515 9710 12585 9730
rect 12645 9730 12740 9770
rect 12645 9710 12715 9730
rect 12430 9695 12486 9701
rect 12430 9635 12434 9695
rect 12515 9685 12715 9710
rect 12770 9701 12800 9889
rect 12744 9695 12800 9701
rect 12486 9635 12744 9655
rect 12796 9635 12800 9695
rect 12430 9625 12800 9635
rect 12830 9955 13200 9965
rect 12830 9895 12834 9955
rect 12886 9935 13144 9955
rect 12830 9889 12886 9895
rect 12830 9701 12860 9889
rect 12915 9880 13115 9905
rect 13196 9895 13200 9955
rect 13144 9889 13200 9895
rect 12915 9860 12985 9880
rect 12890 9820 12985 9860
rect 13045 9860 13115 9880
rect 13045 9820 13140 9860
rect 12890 9770 13140 9820
rect 12890 9730 12985 9770
rect 12915 9710 12985 9730
rect 13045 9730 13140 9770
rect 13045 9710 13115 9730
rect 12830 9695 12886 9701
rect 12830 9635 12834 9695
rect 12915 9685 13115 9710
rect 13170 9701 13200 9889
rect 13144 9695 13200 9701
rect 12886 9635 13144 9655
rect 13196 9635 13200 9695
rect 12830 9625 13200 9635
rect -370 9585 0 9595
rect -370 9525 -366 9585
rect -314 9565 -56 9585
rect -370 9519 -314 9525
rect -370 9331 -340 9519
rect -285 9510 -85 9535
rect -4 9525 0 9585
rect -56 9519 0 9525
rect -285 9490 -215 9510
rect -310 9450 -215 9490
rect -155 9490 -85 9510
rect -155 9450 -60 9490
rect -310 9400 -60 9450
rect -310 9360 -215 9400
rect -285 9340 -215 9360
rect -155 9360 -60 9400
rect -155 9340 -85 9360
rect -370 9325 -314 9331
rect -370 9265 -366 9325
rect -285 9315 -85 9340
rect -30 9331 0 9519
rect -56 9325 0 9331
rect -314 9265 -56 9285
rect -4 9265 0 9325
rect -370 9255 0 9265
rect 30 9585 400 9595
rect 30 9525 34 9585
rect 86 9565 344 9585
rect 30 9519 86 9525
rect 30 9331 60 9519
rect 115 9510 315 9535
rect 396 9525 400 9585
rect 344 9519 400 9525
rect 115 9490 185 9510
rect 90 9450 185 9490
rect 245 9490 315 9510
rect 245 9450 340 9490
rect 90 9400 340 9450
rect 90 9360 185 9400
rect 115 9340 185 9360
rect 245 9360 340 9400
rect 245 9340 315 9360
rect 30 9325 86 9331
rect 30 9265 34 9325
rect 115 9315 315 9340
rect 370 9331 400 9519
rect 344 9325 400 9331
rect 86 9265 344 9285
rect 396 9265 400 9325
rect 30 9255 400 9265
rect 430 9585 800 9595
rect 430 9525 434 9585
rect 486 9565 744 9585
rect 430 9519 486 9525
rect 430 9331 460 9519
rect 515 9510 715 9535
rect 796 9525 800 9585
rect 744 9519 800 9525
rect 515 9490 585 9510
rect 490 9450 585 9490
rect 645 9490 715 9510
rect 645 9450 740 9490
rect 490 9400 740 9450
rect 490 9360 585 9400
rect 515 9340 585 9360
rect 645 9360 740 9400
rect 645 9340 715 9360
rect 430 9325 486 9331
rect 430 9265 434 9325
rect 515 9315 715 9340
rect 770 9331 800 9519
rect 744 9325 800 9331
rect 486 9265 744 9285
rect 796 9265 800 9325
rect 430 9255 800 9265
rect 830 9585 1200 9595
rect 830 9525 834 9585
rect 886 9565 1144 9585
rect 830 9519 886 9525
rect 830 9331 860 9519
rect 915 9510 1115 9535
rect 1196 9525 1200 9585
rect 1144 9519 1200 9525
rect 915 9490 985 9510
rect 890 9450 985 9490
rect 1045 9490 1115 9510
rect 1045 9450 1140 9490
rect 890 9400 1140 9450
rect 890 9360 985 9400
rect 915 9340 985 9360
rect 1045 9360 1140 9400
rect 1045 9340 1115 9360
rect 830 9325 886 9331
rect 830 9265 834 9325
rect 915 9315 1115 9340
rect 1170 9331 1200 9519
rect 1144 9325 1200 9331
rect 886 9265 1144 9285
rect 1196 9265 1200 9325
rect 830 9255 1200 9265
rect 1230 9585 1600 9595
rect 1230 9525 1234 9585
rect 1286 9565 1544 9585
rect 1230 9519 1286 9525
rect 1230 9331 1260 9519
rect 1315 9510 1515 9535
rect 1596 9525 1600 9585
rect 1544 9519 1600 9525
rect 1315 9490 1385 9510
rect 1290 9450 1385 9490
rect 1445 9490 1515 9510
rect 1445 9450 1540 9490
rect 1290 9400 1540 9450
rect 1290 9360 1385 9400
rect 1315 9340 1385 9360
rect 1445 9360 1540 9400
rect 1445 9340 1515 9360
rect 1230 9325 1286 9331
rect 1230 9265 1234 9325
rect 1315 9315 1515 9340
rect 1570 9331 1600 9519
rect 1544 9325 1600 9331
rect 1286 9265 1544 9285
rect 1596 9265 1600 9325
rect 1230 9255 1600 9265
rect 1630 9585 2000 9595
rect 1630 9525 1634 9585
rect 1686 9565 1944 9585
rect 1630 9519 1686 9525
rect 1630 9331 1660 9519
rect 1715 9510 1915 9535
rect 1996 9525 2000 9585
rect 1944 9519 2000 9525
rect 1715 9490 1785 9510
rect 1690 9450 1785 9490
rect 1845 9490 1915 9510
rect 1845 9450 1940 9490
rect 1690 9400 1940 9450
rect 1690 9360 1785 9400
rect 1715 9340 1785 9360
rect 1845 9360 1940 9400
rect 1845 9340 1915 9360
rect 1630 9325 1686 9331
rect 1630 9265 1634 9325
rect 1715 9315 1915 9340
rect 1970 9331 2000 9519
rect 1944 9325 2000 9331
rect 1686 9265 1944 9285
rect 1996 9265 2000 9325
rect 1630 9255 2000 9265
rect 2030 9585 2400 9595
rect 2030 9525 2034 9585
rect 2086 9565 2344 9585
rect 2030 9519 2086 9525
rect 2030 9331 2060 9519
rect 2115 9510 2315 9535
rect 2396 9525 2400 9585
rect 2344 9519 2400 9525
rect 2115 9490 2185 9510
rect 2090 9450 2185 9490
rect 2245 9490 2315 9510
rect 2245 9450 2340 9490
rect 2090 9400 2340 9450
rect 2090 9360 2185 9400
rect 2115 9340 2185 9360
rect 2245 9360 2340 9400
rect 2245 9340 2315 9360
rect 2030 9325 2086 9331
rect 2030 9265 2034 9325
rect 2115 9315 2315 9340
rect 2370 9331 2400 9519
rect 2344 9325 2400 9331
rect 2086 9265 2344 9285
rect 2396 9265 2400 9325
rect 2030 9255 2400 9265
rect 2430 9585 2800 9595
rect 2430 9525 2434 9585
rect 2486 9565 2744 9585
rect 2430 9519 2486 9525
rect 2430 9331 2460 9519
rect 2515 9510 2715 9535
rect 2796 9525 2800 9585
rect 2744 9519 2800 9525
rect 2515 9490 2585 9510
rect 2490 9450 2585 9490
rect 2645 9490 2715 9510
rect 2645 9450 2740 9490
rect 2490 9400 2740 9450
rect 2490 9360 2585 9400
rect 2515 9340 2585 9360
rect 2645 9360 2740 9400
rect 2645 9340 2715 9360
rect 2430 9325 2486 9331
rect 2430 9265 2434 9325
rect 2515 9315 2715 9340
rect 2770 9331 2800 9519
rect 2744 9325 2800 9331
rect 2486 9265 2744 9285
rect 2796 9265 2800 9325
rect 2430 9255 2800 9265
rect 2830 9585 3200 9595
rect 2830 9525 2834 9585
rect 2886 9565 3144 9585
rect 2830 9519 2886 9525
rect 2830 9331 2860 9519
rect 2915 9510 3115 9535
rect 3196 9525 3200 9585
rect 3144 9519 3200 9525
rect 2915 9490 2985 9510
rect 2890 9450 2985 9490
rect 3045 9490 3115 9510
rect 3045 9450 3140 9490
rect 2890 9400 3140 9450
rect 2890 9360 2985 9400
rect 2915 9340 2985 9360
rect 3045 9360 3140 9400
rect 3045 9340 3115 9360
rect 2830 9325 2886 9331
rect 2830 9265 2834 9325
rect 2915 9315 3115 9340
rect 3170 9331 3200 9519
rect 3144 9325 3200 9331
rect 2886 9265 3144 9285
rect 3196 9265 3200 9325
rect 2830 9255 3200 9265
rect 3230 9585 3600 9595
rect 3230 9525 3234 9585
rect 3286 9565 3544 9585
rect 3230 9519 3286 9525
rect 3230 9331 3260 9519
rect 3315 9510 3515 9535
rect 3596 9525 3600 9585
rect 3544 9519 3600 9525
rect 3315 9490 3385 9510
rect 3290 9450 3385 9490
rect 3445 9490 3515 9510
rect 3445 9450 3540 9490
rect 3290 9400 3540 9450
rect 3290 9360 3385 9400
rect 3315 9340 3385 9360
rect 3445 9360 3540 9400
rect 3445 9340 3515 9360
rect 3230 9325 3286 9331
rect 3230 9265 3234 9325
rect 3315 9315 3515 9340
rect 3570 9331 3600 9519
rect 3544 9325 3600 9331
rect 3286 9265 3544 9285
rect 3596 9265 3600 9325
rect 3230 9255 3600 9265
rect 3630 9585 4000 9595
rect 3630 9525 3634 9585
rect 3686 9565 3944 9585
rect 3630 9519 3686 9525
rect 3630 9331 3660 9519
rect 3715 9510 3915 9535
rect 3996 9525 4000 9585
rect 3944 9519 4000 9525
rect 3715 9490 3785 9510
rect 3690 9450 3785 9490
rect 3845 9490 3915 9510
rect 3845 9450 3940 9490
rect 3690 9400 3940 9450
rect 3690 9360 3785 9400
rect 3715 9340 3785 9360
rect 3845 9360 3940 9400
rect 3845 9340 3915 9360
rect 3630 9325 3686 9331
rect 3630 9265 3634 9325
rect 3715 9315 3915 9340
rect 3970 9331 4000 9519
rect 3944 9325 4000 9331
rect 3686 9265 3944 9285
rect 3996 9265 4000 9325
rect 3630 9255 4000 9265
rect 4030 9585 4400 9595
rect 4030 9525 4034 9585
rect 4086 9565 4344 9585
rect 4030 9519 4086 9525
rect 4030 9331 4060 9519
rect 4115 9510 4315 9535
rect 4396 9525 4400 9585
rect 4344 9519 4400 9525
rect 4115 9490 4185 9510
rect 4090 9450 4185 9490
rect 4245 9490 4315 9510
rect 4245 9450 4340 9490
rect 4090 9400 4340 9450
rect 4090 9360 4185 9400
rect 4115 9340 4185 9360
rect 4245 9360 4340 9400
rect 4245 9340 4315 9360
rect 4030 9325 4086 9331
rect 4030 9265 4034 9325
rect 4115 9315 4315 9340
rect 4370 9331 4400 9519
rect 4344 9325 4400 9331
rect 4086 9265 4344 9285
rect 4396 9265 4400 9325
rect 4030 9255 4400 9265
rect 4430 9585 4800 9595
rect 4430 9525 4434 9585
rect 4486 9565 4744 9585
rect 4430 9519 4486 9525
rect 4430 9331 4460 9519
rect 4515 9510 4715 9535
rect 4796 9525 4800 9585
rect 4744 9519 4800 9525
rect 4515 9490 4585 9510
rect 4490 9450 4585 9490
rect 4645 9490 4715 9510
rect 4645 9450 4740 9490
rect 4490 9400 4740 9450
rect 4490 9360 4585 9400
rect 4515 9340 4585 9360
rect 4645 9360 4740 9400
rect 4645 9340 4715 9360
rect 4430 9325 4486 9331
rect 4430 9265 4434 9325
rect 4515 9315 4715 9340
rect 4770 9331 4800 9519
rect 4744 9325 4800 9331
rect 4486 9265 4744 9285
rect 4796 9265 4800 9325
rect 4430 9255 4800 9265
rect 4830 9585 5200 9595
rect 4830 9525 4834 9585
rect 4886 9565 5144 9585
rect 4830 9519 4886 9525
rect 4830 9331 4860 9519
rect 4915 9510 5115 9535
rect 5196 9525 5200 9585
rect 5144 9519 5200 9525
rect 4915 9490 4985 9510
rect 4890 9450 4985 9490
rect 5045 9490 5115 9510
rect 5045 9450 5140 9490
rect 4890 9400 5140 9450
rect 4890 9360 4985 9400
rect 4915 9340 4985 9360
rect 5045 9360 5140 9400
rect 5045 9340 5115 9360
rect 4830 9325 4886 9331
rect 4830 9265 4834 9325
rect 4915 9315 5115 9340
rect 5170 9331 5200 9519
rect 5144 9325 5200 9331
rect 4886 9265 5144 9285
rect 5196 9265 5200 9325
rect 4830 9255 5200 9265
rect 5230 9585 5600 9595
rect 5230 9525 5234 9585
rect 5286 9565 5544 9585
rect 5230 9519 5286 9525
rect 5230 9331 5260 9519
rect 5315 9510 5515 9535
rect 5596 9525 5600 9585
rect 5544 9519 5600 9525
rect 5315 9490 5385 9510
rect 5290 9450 5385 9490
rect 5445 9490 5515 9510
rect 5445 9450 5540 9490
rect 5290 9400 5540 9450
rect 5290 9360 5385 9400
rect 5315 9340 5385 9360
rect 5445 9360 5540 9400
rect 5445 9340 5515 9360
rect 5230 9325 5286 9331
rect 5230 9265 5234 9325
rect 5315 9315 5515 9340
rect 5570 9331 5600 9519
rect 5544 9325 5600 9331
rect 5286 9265 5544 9285
rect 5596 9265 5600 9325
rect 5230 9255 5600 9265
rect 5630 9585 6000 9595
rect 5630 9525 5634 9585
rect 5686 9565 5944 9585
rect 5630 9519 5686 9525
rect 5630 9331 5660 9519
rect 5715 9510 5915 9535
rect 5996 9525 6000 9585
rect 5944 9519 6000 9525
rect 5715 9490 5785 9510
rect 5690 9450 5785 9490
rect 5845 9490 5915 9510
rect 5845 9450 5940 9490
rect 5690 9400 5940 9450
rect 5690 9360 5785 9400
rect 5715 9340 5785 9360
rect 5845 9360 5940 9400
rect 5845 9340 5915 9360
rect 5630 9325 5686 9331
rect 5630 9265 5634 9325
rect 5715 9315 5915 9340
rect 5970 9331 6000 9519
rect 5944 9325 6000 9331
rect 5686 9265 5944 9285
rect 5996 9265 6000 9325
rect 5630 9255 6000 9265
rect 6030 9585 6400 9595
rect 6030 9525 6034 9585
rect 6086 9565 6344 9585
rect 6030 9519 6086 9525
rect 6030 9331 6060 9519
rect 6115 9510 6315 9535
rect 6396 9525 6400 9585
rect 6344 9519 6400 9525
rect 6115 9490 6185 9510
rect 6090 9450 6185 9490
rect 6245 9490 6315 9510
rect 6245 9450 6340 9490
rect 6090 9400 6340 9450
rect 6090 9360 6185 9400
rect 6115 9340 6185 9360
rect 6245 9360 6340 9400
rect 6245 9340 6315 9360
rect 6030 9325 6086 9331
rect 6030 9265 6034 9325
rect 6115 9315 6315 9340
rect 6370 9331 6400 9519
rect 6344 9325 6400 9331
rect 6086 9265 6344 9285
rect 6396 9265 6400 9325
rect 6030 9255 6400 9265
rect 6430 9585 6800 9595
rect 6430 9525 6434 9585
rect 6486 9565 6744 9585
rect 6430 9519 6486 9525
rect 6430 9331 6460 9519
rect 6515 9510 6715 9535
rect 6796 9525 6800 9585
rect 6744 9519 6800 9525
rect 6515 9490 6585 9510
rect 6490 9450 6585 9490
rect 6645 9490 6715 9510
rect 6645 9450 6740 9490
rect 6490 9400 6740 9450
rect 6490 9360 6585 9400
rect 6515 9340 6585 9360
rect 6645 9360 6740 9400
rect 6645 9340 6715 9360
rect 6430 9325 6486 9331
rect 6430 9265 6434 9325
rect 6515 9315 6715 9340
rect 6770 9331 6800 9519
rect 6744 9325 6800 9331
rect 6486 9265 6744 9285
rect 6796 9265 6800 9325
rect 6430 9255 6800 9265
rect 6830 9585 7200 9595
rect 6830 9525 6834 9585
rect 6886 9565 7144 9585
rect 6830 9519 6886 9525
rect 6830 9331 6860 9519
rect 6915 9510 7115 9535
rect 7196 9525 7200 9585
rect 7144 9519 7200 9525
rect 6915 9490 6985 9510
rect 6890 9450 6985 9490
rect 7045 9490 7115 9510
rect 7045 9450 7140 9490
rect 6890 9400 7140 9450
rect 6890 9360 6985 9400
rect 6915 9340 6985 9360
rect 7045 9360 7140 9400
rect 7045 9340 7115 9360
rect 6830 9325 6886 9331
rect 6830 9265 6834 9325
rect 6915 9315 7115 9340
rect 7170 9331 7200 9519
rect 7144 9325 7200 9331
rect 6886 9265 7144 9285
rect 7196 9265 7200 9325
rect 6830 9255 7200 9265
rect 7230 9585 7600 9595
rect 7230 9525 7234 9585
rect 7286 9565 7544 9585
rect 7230 9519 7286 9525
rect 7230 9331 7260 9519
rect 7315 9510 7515 9535
rect 7596 9525 7600 9585
rect 7544 9519 7600 9525
rect 7315 9490 7385 9510
rect 7290 9450 7385 9490
rect 7445 9490 7515 9510
rect 7445 9450 7540 9490
rect 7290 9400 7540 9450
rect 7290 9360 7385 9400
rect 7315 9340 7385 9360
rect 7445 9360 7540 9400
rect 7445 9340 7515 9360
rect 7230 9325 7286 9331
rect 7230 9265 7234 9325
rect 7315 9315 7515 9340
rect 7570 9331 7600 9519
rect 7544 9325 7600 9331
rect 7286 9265 7544 9285
rect 7596 9265 7600 9325
rect 7230 9255 7600 9265
rect 7630 9585 8000 9595
rect 7630 9525 7634 9585
rect 7686 9565 7944 9585
rect 7630 9519 7686 9525
rect 7630 9331 7660 9519
rect 7715 9510 7915 9535
rect 7996 9525 8000 9585
rect 7944 9519 8000 9525
rect 7715 9490 7785 9510
rect 7690 9450 7785 9490
rect 7845 9490 7915 9510
rect 7845 9450 7940 9490
rect 7690 9400 7940 9450
rect 7690 9360 7785 9400
rect 7715 9340 7785 9360
rect 7845 9360 7940 9400
rect 7845 9340 7915 9360
rect 7630 9325 7686 9331
rect 7630 9265 7634 9325
rect 7715 9315 7915 9340
rect 7970 9331 8000 9519
rect 7944 9325 8000 9331
rect 7686 9265 7944 9285
rect 7996 9265 8000 9325
rect 7630 9255 8000 9265
rect 8030 9585 8400 9595
rect 8030 9525 8034 9585
rect 8086 9565 8344 9585
rect 8030 9519 8086 9525
rect 8030 9331 8060 9519
rect 8115 9510 8315 9535
rect 8396 9525 8400 9585
rect 8344 9519 8400 9525
rect 8115 9490 8185 9510
rect 8090 9450 8185 9490
rect 8245 9490 8315 9510
rect 8245 9450 8340 9490
rect 8090 9400 8340 9450
rect 8090 9360 8185 9400
rect 8115 9340 8185 9360
rect 8245 9360 8340 9400
rect 8245 9340 8315 9360
rect 8030 9325 8086 9331
rect 8030 9265 8034 9325
rect 8115 9315 8315 9340
rect 8370 9331 8400 9519
rect 8344 9325 8400 9331
rect 8086 9265 8344 9285
rect 8396 9265 8400 9325
rect 8030 9255 8400 9265
rect 8430 9585 8800 9595
rect 8430 9525 8434 9585
rect 8486 9565 8744 9585
rect 8430 9519 8486 9525
rect 8430 9331 8460 9519
rect 8515 9510 8715 9535
rect 8796 9525 8800 9585
rect 8744 9519 8800 9525
rect 8515 9490 8585 9510
rect 8490 9450 8585 9490
rect 8645 9490 8715 9510
rect 8645 9450 8740 9490
rect 8490 9400 8740 9450
rect 8490 9360 8585 9400
rect 8515 9340 8585 9360
rect 8645 9360 8740 9400
rect 8645 9340 8715 9360
rect 8430 9325 8486 9331
rect 8430 9265 8434 9325
rect 8515 9315 8715 9340
rect 8770 9331 8800 9519
rect 8744 9325 8800 9331
rect 8486 9265 8744 9285
rect 8796 9265 8800 9325
rect 8430 9255 8800 9265
rect 8830 9585 9200 9595
rect 8830 9525 8834 9585
rect 8886 9565 9144 9585
rect 8830 9519 8886 9525
rect 8830 9331 8860 9519
rect 8915 9510 9115 9535
rect 9196 9525 9200 9585
rect 9144 9519 9200 9525
rect 8915 9490 8985 9510
rect 8890 9450 8985 9490
rect 9045 9490 9115 9510
rect 9045 9450 9140 9490
rect 8890 9400 9140 9450
rect 8890 9360 8985 9400
rect 8915 9340 8985 9360
rect 9045 9360 9140 9400
rect 9045 9340 9115 9360
rect 8830 9325 8886 9331
rect 8830 9265 8834 9325
rect 8915 9315 9115 9340
rect 9170 9331 9200 9519
rect 9144 9325 9200 9331
rect 8886 9265 9144 9285
rect 9196 9265 9200 9325
rect 8830 9255 9200 9265
rect 9230 9585 9600 9595
rect 9230 9525 9234 9585
rect 9286 9565 9544 9585
rect 9230 9519 9286 9525
rect 9230 9331 9260 9519
rect 9315 9510 9515 9535
rect 9596 9525 9600 9585
rect 9544 9519 9600 9525
rect 9315 9490 9385 9510
rect 9290 9450 9385 9490
rect 9445 9490 9515 9510
rect 9445 9450 9540 9490
rect 9290 9400 9540 9450
rect 9290 9360 9385 9400
rect 9315 9340 9385 9360
rect 9445 9360 9540 9400
rect 9445 9340 9515 9360
rect 9230 9325 9286 9331
rect 9230 9265 9234 9325
rect 9315 9315 9515 9340
rect 9570 9331 9600 9519
rect 9544 9325 9600 9331
rect 9286 9265 9544 9285
rect 9596 9265 9600 9325
rect 9230 9255 9600 9265
rect 9630 9585 10000 9595
rect 9630 9525 9634 9585
rect 9686 9565 9944 9585
rect 9630 9519 9686 9525
rect 9630 9331 9660 9519
rect 9715 9510 9915 9535
rect 9996 9525 10000 9585
rect 9944 9519 10000 9525
rect 9715 9490 9785 9510
rect 9690 9450 9785 9490
rect 9845 9490 9915 9510
rect 9845 9450 9940 9490
rect 9690 9400 9940 9450
rect 9690 9360 9785 9400
rect 9715 9340 9785 9360
rect 9845 9360 9940 9400
rect 9845 9340 9915 9360
rect 9630 9325 9686 9331
rect 9630 9265 9634 9325
rect 9715 9315 9915 9340
rect 9970 9331 10000 9519
rect 9944 9325 10000 9331
rect 9686 9265 9944 9285
rect 9996 9265 10000 9325
rect 9630 9255 10000 9265
rect 10030 9585 10400 9595
rect 10030 9525 10034 9585
rect 10086 9565 10344 9585
rect 10030 9519 10086 9525
rect 10030 9331 10060 9519
rect 10115 9510 10315 9535
rect 10396 9525 10400 9585
rect 10344 9519 10400 9525
rect 10115 9490 10185 9510
rect 10090 9450 10185 9490
rect 10245 9490 10315 9510
rect 10245 9450 10340 9490
rect 10090 9400 10340 9450
rect 10090 9360 10185 9400
rect 10115 9340 10185 9360
rect 10245 9360 10340 9400
rect 10245 9340 10315 9360
rect 10030 9325 10086 9331
rect 10030 9265 10034 9325
rect 10115 9315 10315 9340
rect 10370 9331 10400 9519
rect 10344 9325 10400 9331
rect 10086 9265 10344 9285
rect 10396 9265 10400 9325
rect 10030 9255 10400 9265
rect 10430 9585 10800 9595
rect 10430 9525 10434 9585
rect 10486 9565 10744 9585
rect 10430 9519 10486 9525
rect 10430 9331 10460 9519
rect 10515 9510 10715 9535
rect 10796 9525 10800 9585
rect 10744 9519 10800 9525
rect 10515 9490 10585 9510
rect 10490 9450 10585 9490
rect 10645 9490 10715 9510
rect 10645 9450 10740 9490
rect 10490 9400 10740 9450
rect 10490 9360 10585 9400
rect 10515 9340 10585 9360
rect 10645 9360 10740 9400
rect 10645 9340 10715 9360
rect 10430 9325 10486 9331
rect 10430 9265 10434 9325
rect 10515 9315 10715 9340
rect 10770 9331 10800 9519
rect 10744 9325 10800 9331
rect 10486 9265 10744 9285
rect 10796 9265 10800 9325
rect 10430 9255 10800 9265
rect 10830 9585 11200 9595
rect 10830 9525 10834 9585
rect 10886 9565 11144 9585
rect 10830 9519 10886 9525
rect 10830 9331 10860 9519
rect 10915 9510 11115 9535
rect 11196 9525 11200 9585
rect 11144 9519 11200 9525
rect 10915 9490 10985 9510
rect 10890 9450 10985 9490
rect 11045 9490 11115 9510
rect 11045 9450 11140 9490
rect 10890 9400 11140 9450
rect 10890 9360 10985 9400
rect 10915 9340 10985 9360
rect 11045 9360 11140 9400
rect 11045 9340 11115 9360
rect 10830 9325 10886 9331
rect 10830 9265 10834 9325
rect 10915 9315 11115 9340
rect 11170 9331 11200 9519
rect 11144 9325 11200 9331
rect 10886 9265 11144 9285
rect 11196 9265 11200 9325
rect 10830 9255 11200 9265
rect 11230 9585 11600 9595
rect 11230 9525 11234 9585
rect 11286 9565 11544 9585
rect 11230 9519 11286 9525
rect 11230 9331 11260 9519
rect 11315 9510 11515 9535
rect 11596 9525 11600 9585
rect 11544 9519 11600 9525
rect 11315 9490 11385 9510
rect 11290 9450 11385 9490
rect 11445 9490 11515 9510
rect 11445 9450 11540 9490
rect 11290 9400 11540 9450
rect 11290 9360 11385 9400
rect 11315 9340 11385 9360
rect 11445 9360 11540 9400
rect 11445 9340 11515 9360
rect 11230 9325 11286 9331
rect 11230 9265 11234 9325
rect 11315 9315 11515 9340
rect 11570 9331 11600 9519
rect 11544 9325 11600 9331
rect 11286 9265 11544 9285
rect 11596 9265 11600 9325
rect 11230 9255 11600 9265
rect 11630 9585 12000 9595
rect 11630 9525 11634 9585
rect 11686 9565 11944 9585
rect 11630 9519 11686 9525
rect 11630 9331 11660 9519
rect 11715 9510 11915 9535
rect 11996 9525 12000 9585
rect 11944 9519 12000 9525
rect 11715 9490 11785 9510
rect 11690 9450 11785 9490
rect 11845 9490 11915 9510
rect 11845 9450 11940 9490
rect 11690 9400 11940 9450
rect 11690 9360 11785 9400
rect 11715 9340 11785 9360
rect 11845 9360 11940 9400
rect 11845 9340 11915 9360
rect 11630 9325 11686 9331
rect 11630 9265 11634 9325
rect 11715 9315 11915 9340
rect 11970 9331 12000 9519
rect 11944 9325 12000 9331
rect 11686 9265 11944 9285
rect 11996 9265 12000 9325
rect 11630 9255 12000 9265
rect 12030 9585 12400 9595
rect 12030 9525 12034 9585
rect 12086 9565 12344 9585
rect 12030 9519 12086 9525
rect 12030 9331 12060 9519
rect 12115 9510 12315 9535
rect 12396 9525 12400 9585
rect 12344 9519 12400 9525
rect 12115 9490 12185 9510
rect 12090 9450 12185 9490
rect 12245 9490 12315 9510
rect 12245 9450 12340 9490
rect 12090 9400 12340 9450
rect 12090 9360 12185 9400
rect 12115 9340 12185 9360
rect 12245 9360 12340 9400
rect 12245 9340 12315 9360
rect 12030 9325 12086 9331
rect 12030 9265 12034 9325
rect 12115 9315 12315 9340
rect 12370 9331 12400 9519
rect 12344 9325 12400 9331
rect 12086 9265 12344 9285
rect 12396 9265 12400 9325
rect 12030 9255 12400 9265
rect 12430 9585 12800 9595
rect 12430 9525 12434 9585
rect 12486 9565 12744 9585
rect 12430 9519 12486 9525
rect 12430 9331 12460 9519
rect 12515 9510 12715 9535
rect 12796 9525 12800 9585
rect 12744 9519 12800 9525
rect 12515 9490 12585 9510
rect 12490 9450 12585 9490
rect 12645 9490 12715 9510
rect 12645 9450 12740 9490
rect 12490 9400 12740 9450
rect 12490 9360 12585 9400
rect 12515 9340 12585 9360
rect 12645 9360 12740 9400
rect 12645 9340 12715 9360
rect 12430 9325 12486 9331
rect 12430 9265 12434 9325
rect 12515 9315 12715 9340
rect 12770 9331 12800 9519
rect 12744 9325 12800 9331
rect 12486 9265 12744 9285
rect 12796 9265 12800 9325
rect 12430 9255 12800 9265
rect 12830 9585 13200 9595
rect 12830 9525 12834 9585
rect 12886 9565 13144 9585
rect 12830 9519 12886 9525
rect 12830 9331 12860 9519
rect 12915 9510 13115 9535
rect 13196 9525 13200 9585
rect 13144 9519 13200 9525
rect 12915 9490 12985 9510
rect 12890 9450 12985 9490
rect 13045 9490 13115 9510
rect 13045 9450 13140 9490
rect 12890 9400 13140 9450
rect 12890 9360 12985 9400
rect 12915 9340 12985 9360
rect 13045 9360 13140 9400
rect 13045 9340 13115 9360
rect 12830 9325 12886 9331
rect 12830 9265 12834 9325
rect 12915 9315 13115 9340
rect 13170 9331 13200 9519
rect 13144 9325 13200 9331
rect 12886 9265 13144 9285
rect 13196 9265 13200 9325
rect 12830 9255 13200 9265
rect -370 9215 0 9225
rect -370 9155 -366 9215
rect -314 9195 -56 9215
rect -370 9149 -314 9155
rect -370 8961 -340 9149
rect -285 9140 -85 9165
rect -4 9155 0 9215
rect -56 9149 0 9155
rect -285 9120 -215 9140
rect -310 9080 -215 9120
rect -155 9120 -85 9140
rect -155 9080 -60 9120
rect -310 9030 -60 9080
rect -310 8990 -215 9030
rect -285 8970 -215 8990
rect -155 8990 -60 9030
rect -155 8970 -85 8990
rect -370 8955 -314 8961
rect -370 8895 -366 8955
rect -285 8945 -85 8970
rect -30 8961 0 9149
rect -56 8955 0 8961
rect -314 8895 -56 8915
rect -4 8895 0 8955
rect -370 8885 0 8895
rect 30 9215 400 9225
rect 30 9155 34 9215
rect 86 9195 344 9215
rect 30 9149 86 9155
rect 30 8961 60 9149
rect 115 9140 315 9165
rect 396 9155 400 9215
rect 344 9149 400 9155
rect 115 9120 185 9140
rect 90 9080 185 9120
rect 245 9120 315 9140
rect 245 9080 340 9120
rect 90 9030 340 9080
rect 90 8990 185 9030
rect 115 8970 185 8990
rect 245 8990 340 9030
rect 245 8970 315 8990
rect 30 8955 86 8961
rect 30 8895 34 8955
rect 115 8945 315 8970
rect 370 8961 400 9149
rect 344 8955 400 8961
rect 86 8895 344 8915
rect 396 8895 400 8955
rect 30 8885 400 8895
rect 430 9215 800 9225
rect 430 9155 434 9215
rect 486 9195 744 9215
rect 430 9149 486 9155
rect 430 8961 460 9149
rect 515 9140 715 9165
rect 796 9155 800 9215
rect 744 9149 800 9155
rect 515 9120 585 9140
rect 490 9080 585 9120
rect 645 9120 715 9140
rect 645 9080 740 9120
rect 490 9030 740 9080
rect 490 8990 585 9030
rect 515 8970 585 8990
rect 645 8990 740 9030
rect 645 8970 715 8990
rect 430 8955 486 8961
rect 430 8895 434 8955
rect 515 8945 715 8970
rect 770 8961 800 9149
rect 744 8955 800 8961
rect 486 8895 744 8915
rect 796 8895 800 8955
rect 430 8885 800 8895
rect 830 9215 1200 9225
rect 830 9155 834 9215
rect 886 9195 1144 9215
rect 830 9149 886 9155
rect 830 8961 860 9149
rect 915 9140 1115 9165
rect 1196 9155 1200 9215
rect 1144 9149 1200 9155
rect 915 9120 985 9140
rect 890 9080 985 9120
rect 1045 9120 1115 9140
rect 1045 9080 1140 9120
rect 890 9030 1140 9080
rect 890 8990 985 9030
rect 915 8970 985 8990
rect 1045 8990 1140 9030
rect 1045 8970 1115 8990
rect 830 8955 886 8961
rect 830 8895 834 8955
rect 915 8945 1115 8970
rect 1170 8961 1200 9149
rect 1144 8955 1200 8961
rect 886 8895 1144 8915
rect 1196 8895 1200 8955
rect 830 8885 1200 8895
rect 1230 9215 1600 9225
rect 1230 9155 1234 9215
rect 1286 9195 1544 9215
rect 1230 9149 1286 9155
rect 1230 8961 1260 9149
rect 1315 9140 1515 9165
rect 1596 9155 1600 9215
rect 1544 9149 1600 9155
rect 1315 9120 1385 9140
rect 1290 9080 1385 9120
rect 1445 9120 1515 9140
rect 1445 9080 1540 9120
rect 1290 9030 1540 9080
rect 1290 8990 1385 9030
rect 1315 8970 1385 8990
rect 1445 8990 1540 9030
rect 1445 8970 1515 8990
rect 1230 8955 1286 8961
rect 1230 8895 1234 8955
rect 1315 8945 1515 8970
rect 1570 8961 1600 9149
rect 1544 8955 1600 8961
rect 1286 8895 1544 8915
rect 1596 8895 1600 8955
rect 1230 8885 1600 8895
rect 1630 9215 2000 9225
rect 1630 9155 1634 9215
rect 1686 9195 1944 9215
rect 1630 9149 1686 9155
rect 1630 8961 1660 9149
rect 1715 9140 1915 9165
rect 1996 9155 2000 9215
rect 1944 9149 2000 9155
rect 1715 9120 1785 9140
rect 1690 9080 1785 9120
rect 1845 9120 1915 9140
rect 1845 9080 1940 9120
rect 1690 9030 1940 9080
rect 1690 8990 1785 9030
rect 1715 8970 1785 8990
rect 1845 8990 1940 9030
rect 1845 8970 1915 8990
rect 1630 8955 1686 8961
rect 1630 8895 1634 8955
rect 1715 8945 1915 8970
rect 1970 8961 2000 9149
rect 1944 8955 2000 8961
rect 1686 8895 1944 8915
rect 1996 8895 2000 8955
rect 1630 8885 2000 8895
rect 2030 9215 2400 9225
rect 2030 9155 2034 9215
rect 2086 9195 2344 9215
rect 2030 9149 2086 9155
rect 2030 8961 2060 9149
rect 2115 9140 2315 9165
rect 2396 9155 2400 9215
rect 2344 9149 2400 9155
rect 2115 9120 2185 9140
rect 2090 9080 2185 9120
rect 2245 9120 2315 9140
rect 2245 9080 2340 9120
rect 2090 9030 2340 9080
rect 2090 8990 2185 9030
rect 2115 8970 2185 8990
rect 2245 8990 2340 9030
rect 2245 8970 2315 8990
rect 2030 8955 2086 8961
rect 2030 8895 2034 8955
rect 2115 8945 2315 8970
rect 2370 8961 2400 9149
rect 2344 8955 2400 8961
rect 2086 8895 2344 8915
rect 2396 8895 2400 8955
rect 2030 8885 2400 8895
rect 2430 9215 2800 9225
rect 2430 9155 2434 9215
rect 2486 9195 2744 9215
rect 2430 9149 2486 9155
rect 2430 8961 2460 9149
rect 2515 9140 2715 9165
rect 2796 9155 2800 9215
rect 2744 9149 2800 9155
rect 2515 9120 2585 9140
rect 2490 9080 2585 9120
rect 2645 9120 2715 9140
rect 2645 9080 2740 9120
rect 2490 9030 2740 9080
rect 2490 8990 2585 9030
rect 2515 8970 2585 8990
rect 2645 8990 2740 9030
rect 2645 8970 2715 8990
rect 2430 8955 2486 8961
rect 2430 8895 2434 8955
rect 2515 8945 2715 8970
rect 2770 8961 2800 9149
rect 2744 8955 2800 8961
rect 2486 8895 2744 8915
rect 2796 8895 2800 8955
rect 2430 8885 2800 8895
rect 2830 9215 3200 9225
rect 2830 9155 2834 9215
rect 2886 9195 3144 9215
rect 2830 9149 2886 9155
rect 2830 8961 2860 9149
rect 2915 9140 3115 9165
rect 3196 9155 3200 9215
rect 3144 9149 3200 9155
rect 2915 9120 2985 9140
rect 2890 9080 2985 9120
rect 3045 9120 3115 9140
rect 3045 9080 3140 9120
rect 2890 9030 3140 9080
rect 2890 8990 2985 9030
rect 2915 8970 2985 8990
rect 3045 8990 3140 9030
rect 3045 8970 3115 8990
rect 2830 8955 2886 8961
rect 2830 8895 2834 8955
rect 2915 8945 3115 8970
rect 3170 8961 3200 9149
rect 3144 8955 3200 8961
rect 2886 8895 3144 8915
rect 3196 8895 3200 8955
rect 2830 8885 3200 8895
rect 3230 9215 3600 9225
rect 3230 9155 3234 9215
rect 3286 9195 3544 9215
rect 3230 9149 3286 9155
rect 3230 8961 3260 9149
rect 3315 9140 3515 9165
rect 3596 9155 3600 9215
rect 3544 9149 3600 9155
rect 3315 9120 3385 9140
rect 3290 9080 3385 9120
rect 3445 9120 3515 9140
rect 3445 9080 3540 9120
rect 3290 9030 3540 9080
rect 3290 8990 3385 9030
rect 3315 8970 3385 8990
rect 3445 8990 3540 9030
rect 3445 8970 3515 8990
rect 3230 8955 3286 8961
rect 3230 8895 3234 8955
rect 3315 8945 3515 8970
rect 3570 8961 3600 9149
rect 3544 8955 3600 8961
rect 3286 8895 3544 8915
rect 3596 8895 3600 8955
rect 3230 8885 3600 8895
rect 3630 9215 4000 9225
rect 3630 9155 3634 9215
rect 3686 9195 3944 9215
rect 3630 9149 3686 9155
rect 3630 8961 3660 9149
rect 3715 9140 3915 9165
rect 3996 9155 4000 9215
rect 3944 9149 4000 9155
rect 3715 9120 3785 9140
rect 3690 9080 3785 9120
rect 3845 9120 3915 9140
rect 3845 9080 3940 9120
rect 3690 9030 3940 9080
rect 3690 8990 3785 9030
rect 3715 8970 3785 8990
rect 3845 8990 3940 9030
rect 3845 8970 3915 8990
rect 3630 8955 3686 8961
rect 3630 8895 3634 8955
rect 3715 8945 3915 8970
rect 3970 8961 4000 9149
rect 3944 8955 4000 8961
rect 3686 8895 3944 8915
rect 3996 8895 4000 8955
rect 3630 8885 4000 8895
rect 4030 9215 4400 9225
rect 4030 9155 4034 9215
rect 4086 9195 4344 9215
rect 4030 9149 4086 9155
rect 4030 8961 4060 9149
rect 4115 9140 4315 9165
rect 4396 9155 4400 9215
rect 4344 9149 4400 9155
rect 4115 9120 4185 9140
rect 4090 9080 4185 9120
rect 4245 9120 4315 9140
rect 4245 9080 4340 9120
rect 4090 9030 4340 9080
rect 4090 8990 4185 9030
rect 4115 8970 4185 8990
rect 4245 8990 4340 9030
rect 4245 8970 4315 8990
rect 4030 8955 4086 8961
rect 4030 8895 4034 8955
rect 4115 8945 4315 8970
rect 4370 8961 4400 9149
rect 4344 8955 4400 8961
rect 4086 8895 4344 8915
rect 4396 8895 4400 8955
rect 4030 8885 4400 8895
rect 4430 9215 4800 9225
rect 4430 9155 4434 9215
rect 4486 9195 4744 9215
rect 4430 9149 4486 9155
rect 4430 8961 4460 9149
rect 4515 9140 4715 9165
rect 4796 9155 4800 9215
rect 4744 9149 4800 9155
rect 4515 9120 4585 9140
rect 4490 9080 4585 9120
rect 4645 9120 4715 9140
rect 4645 9080 4740 9120
rect 4490 9030 4740 9080
rect 4490 8990 4585 9030
rect 4515 8970 4585 8990
rect 4645 8990 4740 9030
rect 4645 8970 4715 8990
rect 4430 8955 4486 8961
rect 4430 8895 4434 8955
rect 4515 8945 4715 8970
rect 4770 8961 4800 9149
rect 4744 8955 4800 8961
rect 4486 8895 4744 8915
rect 4796 8895 4800 8955
rect 4430 8885 4800 8895
rect 4830 9215 5200 9225
rect 4830 9155 4834 9215
rect 4886 9195 5144 9215
rect 4830 9149 4886 9155
rect 4830 8961 4860 9149
rect 4915 9140 5115 9165
rect 5196 9155 5200 9215
rect 5144 9149 5200 9155
rect 4915 9120 4985 9140
rect 4890 9080 4985 9120
rect 5045 9120 5115 9140
rect 5045 9080 5140 9120
rect 4890 9030 5140 9080
rect 4890 8990 4985 9030
rect 4915 8970 4985 8990
rect 5045 8990 5140 9030
rect 5045 8970 5115 8990
rect 4830 8955 4886 8961
rect 4830 8895 4834 8955
rect 4915 8945 5115 8970
rect 5170 8961 5200 9149
rect 5144 8955 5200 8961
rect 4886 8895 5144 8915
rect 5196 8895 5200 8955
rect 4830 8885 5200 8895
rect 5230 9215 5600 9225
rect 5230 9155 5234 9215
rect 5286 9195 5544 9215
rect 5230 9149 5286 9155
rect 5230 8961 5260 9149
rect 5315 9140 5515 9165
rect 5596 9155 5600 9215
rect 5544 9149 5600 9155
rect 5315 9120 5385 9140
rect 5290 9080 5385 9120
rect 5445 9120 5515 9140
rect 5445 9080 5540 9120
rect 5290 9030 5540 9080
rect 5290 8990 5385 9030
rect 5315 8970 5385 8990
rect 5445 8990 5540 9030
rect 5445 8970 5515 8990
rect 5230 8955 5286 8961
rect 5230 8895 5234 8955
rect 5315 8945 5515 8970
rect 5570 8961 5600 9149
rect 5544 8955 5600 8961
rect 5286 8895 5544 8915
rect 5596 8895 5600 8955
rect 5230 8885 5600 8895
rect 5630 9215 6000 9225
rect 5630 9155 5634 9215
rect 5686 9195 5944 9215
rect 5630 9149 5686 9155
rect 5630 8961 5660 9149
rect 5715 9140 5915 9165
rect 5996 9155 6000 9215
rect 5944 9149 6000 9155
rect 5715 9120 5785 9140
rect 5690 9080 5785 9120
rect 5845 9120 5915 9140
rect 5845 9080 5940 9120
rect 5690 9030 5940 9080
rect 5690 8990 5785 9030
rect 5715 8970 5785 8990
rect 5845 8990 5940 9030
rect 5845 8970 5915 8990
rect 5630 8955 5686 8961
rect 5630 8895 5634 8955
rect 5715 8945 5915 8970
rect 5970 8961 6000 9149
rect 5944 8955 6000 8961
rect 5686 8895 5944 8915
rect 5996 8895 6000 8955
rect 5630 8885 6000 8895
rect 6030 9215 6400 9225
rect 6030 9155 6034 9215
rect 6086 9195 6344 9215
rect 6030 9149 6086 9155
rect 6030 8961 6060 9149
rect 6115 9140 6315 9165
rect 6396 9155 6400 9215
rect 6344 9149 6400 9155
rect 6115 9120 6185 9140
rect 6090 9080 6185 9120
rect 6245 9120 6315 9140
rect 6245 9080 6340 9120
rect 6090 9030 6340 9080
rect 6090 8990 6185 9030
rect 6115 8970 6185 8990
rect 6245 8990 6340 9030
rect 6245 8970 6315 8990
rect 6030 8955 6086 8961
rect 6030 8895 6034 8955
rect 6115 8945 6315 8970
rect 6370 8961 6400 9149
rect 6344 8955 6400 8961
rect 6086 8895 6344 8915
rect 6396 8895 6400 8955
rect 6030 8885 6400 8895
rect 6430 9215 6800 9225
rect 6430 9155 6434 9215
rect 6486 9195 6744 9215
rect 6430 9149 6486 9155
rect 6430 8961 6460 9149
rect 6515 9140 6715 9165
rect 6796 9155 6800 9215
rect 6744 9149 6800 9155
rect 6515 9120 6585 9140
rect 6490 9080 6585 9120
rect 6645 9120 6715 9140
rect 6645 9080 6740 9120
rect 6490 9030 6740 9080
rect 6490 8990 6585 9030
rect 6515 8970 6585 8990
rect 6645 8990 6740 9030
rect 6645 8970 6715 8990
rect 6430 8955 6486 8961
rect 6430 8895 6434 8955
rect 6515 8945 6715 8970
rect 6770 8961 6800 9149
rect 6744 8955 6800 8961
rect 6486 8895 6744 8915
rect 6796 8895 6800 8955
rect 6430 8885 6800 8895
rect 6830 9215 7200 9225
rect 6830 9155 6834 9215
rect 6886 9195 7144 9215
rect 6830 9149 6886 9155
rect 6830 8961 6860 9149
rect 6915 9140 7115 9165
rect 7196 9155 7200 9215
rect 7144 9149 7200 9155
rect 6915 9120 6985 9140
rect 6890 9080 6985 9120
rect 7045 9120 7115 9140
rect 7045 9080 7140 9120
rect 6890 9030 7140 9080
rect 6890 8990 6985 9030
rect 6915 8970 6985 8990
rect 7045 8990 7140 9030
rect 7045 8970 7115 8990
rect 6830 8955 6886 8961
rect 6830 8895 6834 8955
rect 6915 8945 7115 8970
rect 7170 8961 7200 9149
rect 7144 8955 7200 8961
rect 6886 8895 7144 8915
rect 7196 8895 7200 8955
rect 6830 8885 7200 8895
rect 7230 9215 7600 9225
rect 7230 9155 7234 9215
rect 7286 9195 7544 9215
rect 7230 9149 7286 9155
rect 7230 8961 7260 9149
rect 7315 9140 7515 9165
rect 7596 9155 7600 9215
rect 7544 9149 7600 9155
rect 7315 9120 7385 9140
rect 7290 9080 7385 9120
rect 7445 9120 7515 9140
rect 7445 9080 7540 9120
rect 7290 9030 7540 9080
rect 7290 8990 7385 9030
rect 7315 8970 7385 8990
rect 7445 8990 7540 9030
rect 7445 8970 7515 8990
rect 7230 8955 7286 8961
rect 7230 8895 7234 8955
rect 7315 8945 7515 8970
rect 7570 8961 7600 9149
rect 7544 8955 7600 8961
rect 7286 8895 7544 8915
rect 7596 8895 7600 8955
rect 7230 8885 7600 8895
rect 7630 9215 8000 9225
rect 7630 9155 7634 9215
rect 7686 9195 7944 9215
rect 7630 9149 7686 9155
rect 7630 8961 7660 9149
rect 7715 9140 7915 9165
rect 7996 9155 8000 9215
rect 7944 9149 8000 9155
rect 7715 9120 7785 9140
rect 7690 9080 7785 9120
rect 7845 9120 7915 9140
rect 7845 9080 7940 9120
rect 7690 9030 7940 9080
rect 7690 8990 7785 9030
rect 7715 8970 7785 8990
rect 7845 8990 7940 9030
rect 7845 8970 7915 8990
rect 7630 8955 7686 8961
rect 7630 8895 7634 8955
rect 7715 8945 7915 8970
rect 7970 8961 8000 9149
rect 7944 8955 8000 8961
rect 7686 8895 7944 8915
rect 7996 8895 8000 8955
rect 7630 8885 8000 8895
rect 8030 9215 8400 9225
rect 8030 9155 8034 9215
rect 8086 9195 8344 9215
rect 8030 9149 8086 9155
rect 8030 8961 8060 9149
rect 8115 9140 8315 9165
rect 8396 9155 8400 9215
rect 8344 9149 8400 9155
rect 8115 9120 8185 9140
rect 8090 9080 8185 9120
rect 8245 9120 8315 9140
rect 8245 9080 8340 9120
rect 8090 9030 8340 9080
rect 8090 8990 8185 9030
rect 8115 8970 8185 8990
rect 8245 8990 8340 9030
rect 8245 8970 8315 8990
rect 8030 8955 8086 8961
rect 8030 8895 8034 8955
rect 8115 8945 8315 8970
rect 8370 8961 8400 9149
rect 8344 8955 8400 8961
rect 8086 8895 8344 8915
rect 8396 8895 8400 8955
rect 8030 8885 8400 8895
rect 8430 9215 8800 9225
rect 8430 9155 8434 9215
rect 8486 9195 8744 9215
rect 8430 9149 8486 9155
rect 8430 8961 8460 9149
rect 8515 9140 8715 9165
rect 8796 9155 8800 9215
rect 8744 9149 8800 9155
rect 8515 9120 8585 9140
rect 8490 9080 8585 9120
rect 8645 9120 8715 9140
rect 8645 9080 8740 9120
rect 8490 9030 8740 9080
rect 8490 8990 8585 9030
rect 8515 8970 8585 8990
rect 8645 8990 8740 9030
rect 8645 8970 8715 8990
rect 8430 8955 8486 8961
rect 8430 8895 8434 8955
rect 8515 8945 8715 8970
rect 8770 8961 8800 9149
rect 8744 8955 8800 8961
rect 8486 8895 8744 8915
rect 8796 8895 8800 8955
rect 8430 8885 8800 8895
rect 8830 9215 9200 9225
rect 8830 9155 8834 9215
rect 8886 9195 9144 9215
rect 8830 9149 8886 9155
rect 8830 8961 8860 9149
rect 8915 9140 9115 9165
rect 9196 9155 9200 9215
rect 9144 9149 9200 9155
rect 8915 9120 8985 9140
rect 8890 9080 8985 9120
rect 9045 9120 9115 9140
rect 9045 9080 9140 9120
rect 8890 9030 9140 9080
rect 8890 8990 8985 9030
rect 8915 8970 8985 8990
rect 9045 8990 9140 9030
rect 9045 8970 9115 8990
rect 8830 8955 8886 8961
rect 8830 8895 8834 8955
rect 8915 8945 9115 8970
rect 9170 8961 9200 9149
rect 9144 8955 9200 8961
rect 8886 8895 9144 8915
rect 9196 8895 9200 8955
rect 8830 8885 9200 8895
rect 9230 9215 9600 9225
rect 9230 9155 9234 9215
rect 9286 9195 9544 9215
rect 9230 9149 9286 9155
rect 9230 8961 9260 9149
rect 9315 9140 9515 9165
rect 9596 9155 9600 9215
rect 9544 9149 9600 9155
rect 9315 9120 9385 9140
rect 9290 9080 9385 9120
rect 9445 9120 9515 9140
rect 9445 9080 9540 9120
rect 9290 9030 9540 9080
rect 9290 8990 9385 9030
rect 9315 8970 9385 8990
rect 9445 8990 9540 9030
rect 9445 8970 9515 8990
rect 9230 8955 9286 8961
rect 9230 8895 9234 8955
rect 9315 8945 9515 8970
rect 9570 8961 9600 9149
rect 9544 8955 9600 8961
rect 9286 8895 9544 8915
rect 9596 8895 9600 8955
rect 9230 8885 9600 8895
rect 9630 9215 10000 9225
rect 9630 9155 9634 9215
rect 9686 9195 9944 9215
rect 9630 9149 9686 9155
rect 9630 8961 9660 9149
rect 9715 9140 9915 9165
rect 9996 9155 10000 9215
rect 9944 9149 10000 9155
rect 9715 9120 9785 9140
rect 9690 9080 9785 9120
rect 9845 9120 9915 9140
rect 9845 9080 9940 9120
rect 9690 9030 9940 9080
rect 9690 8990 9785 9030
rect 9715 8970 9785 8990
rect 9845 8990 9940 9030
rect 9845 8970 9915 8990
rect 9630 8955 9686 8961
rect 9630 8895 9634 8955
rect 9715 8945 9915 8970
rect 9970 8961 10000 9149
rect 9944 8955 10000 8961
rect 9686 8895 9944 8915
rect 9996 8895 10000 8955
rect 9630 8885 10000 8895
rect 10030 9215 10400 9225
rect 10030 9155 10034 9215
rect 10086 9195 10344 9215
rect 10030 9149 10086 9155
rect 10030 8961 10060 9149
rect 10115 9140 10315 9165
rect 10396 9155 10400 9215
rect 10344 9149 10400 9155
rect 10115 9120 10185 9140
rect 10090 9080 10185 9120
rect 10245 9120 10315 9140
rect 10245 9080 10340 9120
rect 10090 9030 10340 9080
rect 10090 8990 10185 9030
rect 10115 8970 10185 8990
rect 10245 8990 10340 9030
rect 10245 8970 10315 8990
rect 10030 8955 10086 8961
rect 10030 8895 10034 8955
rect 10115 8945 10315 8970
rect 10370 8961 10400 9149
rect 10344 8955 10400 8961
rect 10086 8895 10344 8915
rect 10396 8895 10400 8955
rect 10030 8885 10400 8895
rect 10430 9215 10800 9225
rect 10430 9155 10434 9215
rect 10486 9195 10744 9215
rect 10430 9149 10486 9155
rect 10430 8961 10460 9149
rect 10515 9140 10715 9165
rect 10796 9155 10800 9215
rect 10744 9149 10800 9155
rect 10515 9120 10585 9140
rect 10490 9080 10585 9120
rect 10645 9120 10715 9140
rect 10645 9080 10740 9120
rect 10490 9030 10740 9080
rect 10490 8990 10585 9030
rect 10515 8970 10585 8990
rect 10645 8990 10740 9030
rect 10645 8970 10715 8990
rect 10430 8955 10486 8961
rect 10430 8895 10434 8955
rect 10515 8945 10715 8970
rect 10770 8961 10800 9149
rect 10744 8955 10800 8961
rect 10486 8895 10744 8915
rect 10796 8895 10800 8955
rect 10430 8885 10800 8895
rect 10830 9215 11200 9225
rect 10830 9155 10834 9215
rect 10886 9195 11144 9215
rect 10830 9149 10886 9155
rect 10830 8961 10860 9149
rect 10915 9140 11115 9165
rect 11196 9155 11200 9215
rect 11144 9149 11200 9155
rect 10915 9120 10985 9140
rect 10890 9080 10985 9120
rect 11045 9120 11115 9140
rect 11045 9080 11140 9120
rect 10890 9030 11140 9080
rect 10890 8990 10985 9030
rect 10915 8970 10985 8990
rect 11045 8990 11140 9030
rect 11045 8970 11115 8990
rect 10830 8955 10886 8961
rect 10830 8895 10834 8955
rect 10915 8945 11115 8970
rect 11170 8961 11200 9149
rect 11144 8955 11200 8961
rect 10886 8895 11144 8915
rect 11196 8895 11200 8955
rect 10830 8885 11200 8895
rect 11230 9215 11600 9225
rect 11230 9155 11234 9215
rect 11286 9195 11544 9215
rect 11230 9149 11286 9155
rect 11230 8961 11260 9149
rect 11315 9140 11515 9165
rect 11596 9155 11600 9215
rect 11544 9149 11600 9155
rect 11315 9120 11385 9140
rect 11290 9080 11385 9120
rect 11445 9120 11515 9140
rect 11445 9080 11540 9120
rect 11290 9030 11540 9080
rect 11290 8990 11385 9030
rect 11315 8970 11385 8990
rect 11445 8990 11540 9030
rect 11445 8970 11515 8990
rect 11230 8955 11286 8961
rect 11230 8895 11234 8955
rect 11315 8945 11515 8970
rect 11570 8961 11600 9149
rect 11544 8955 11600 8961
rect 11286 8895 11544 8915
rect 11596 8895 11600 8955
rect 11230 8885 11600 8895
rect 11630 9215 12000 9225
rect 11630 9155 11634 9215
rect 11686 9195 11944 9215
rect 11630 9149 11686 9155
rect 11630 8961 11660 9149
rect 11715 9140 11915 9165
rect 11996 9155 12000 9215
rect 11944 9149 12000 9155
rect 11715 9120 11785 9140
rect 11690 9080 11785 9120
rect 11845 9120 11915 9140
rect 11845 9080 11940 9120
rect 11690 9030 11940 9080
rect 11690 8990 11785 9030
rect 11715 8970 11785 8990
rect 11845 8990 11940 9030
rect 11845 8970 11915 8990
rect 11630 8955 11686 8961
rect 11630 8895 11634 8955
rect 11715 8945 11915 8970
rect 11970 8961 12000 9149
rect 11944 8955 12000 8961
rect 11686 8895 11944 8915
rect 11996 8895 12000 8955
rect 11630 8885 12000 8895
rect 12030 9215 12400 9225
rect 12030 9155 12034 9215
rect 12086 9195 12344 9215
rect 12030 9149 12086 9155
rect 12030 8961 12060 9149
rect 12115 9140 12315 9165
rect 12396 9155 12400 9215
rect 12344 9149 12400 9155
rect 12115 9120 12185 9140
rect 12090 9080 12185 9120
rect 12245 9120 12315 9140
rect 12245 9080 12340 9120
rect 12090 9030 12340 9080
rect 12090 8990 12185 9030
rect 12115 8970 12185 8990
rect 12245 8990 12340 9030
rect 12245 8970 12315 8990
rect 12030 8955 12086 8961
rect 12030 8895 12034 8955
rect 12115 8945 12315 8970
rect 12370 8961 12400 9149
rect 12344 8955 12400 8961
rect 12086 8895 12344 8915
rect 12396 8895 12400 8955
rect 12030 8885 12400 8895
rect 12430 9215 12800 9225
rect 12430 9155 12434 9215
rect 12486 9195 12744 9215
rect 12430 9149 12486 9155
rect 12430 8961 12460 9149
rect 12515 9140 12715 9165
rect 12796 9155 12800 9215
rect 12744 9149 12800 9155
rect 12515 9120 12585 9140
rect 12490 9080 12585 9120
rect 12645 9120 12715 9140
rect 12645 9080 12740 9120
rect 12490 9030 12740 9080
rect 12490 8990 12585 9030
rect 12515 8970 12585 8990
rect 12645 8990 12740 9030
rect 12645 8970 12715 8990
rect 12430 8955 12486 8961
rect 12430 8895 12434 8955
rect 12515 8945 12715 8970
rect 12770 8961 12800 9149
rect 12744 8955 12800 8961
rect 12486 8895 12744 8915
rect 12796 8895 12800 8955
rect 12430 8885 12800 8895
rect 12830 9215 13200 9225
rect 12830 9155 12834 9215
rect 12886 9195 13144 9215
rect 12830 9149 12886 9155
rect 12830 8961 12860 9149
rect 12915 9140 13115 9165
rect 13196 9155 13200 9215
rect 13144 9149 13200 9155
rect 12915 9120 12985 9140
rect 12890 9080 12985 9120
rect 13045 9120 13115 9140
rect 13045 9080 13140 9120
rect 12890 9030 13140 9080
rect 12890 8990 12985 9030
rect 12915 8970 12985 8990
rect 13045 8990 13140 9030
rect 13045 8970 13115 8990
rect 12830 8955 12886 8961
rect 12830 8895 12834 8955
rect 12915 8945 13115 8970
rect 13170 8961 13200 9149
rect 13144 8955 13200 8961
rect 12886 8895 13144 8915
rect 13196 8895 13200 8955
rect 12830 8885 13200 8895
rect -370 8845 0 8855
rect -370 8785 -366 8845
rect -314 8825 -56 8845
rect -370 8779 -314 8785
rect -370 8591 -340 8779
rect -285 8770 -85 8795
rect -4 8785 0 8845
rect -56 8779 0 8785
rect -285 8750 -215 8770
rect -310 8710 -215 8750
rect -155 8750 -85 8770
rect -155 8710 -60 8750
rect -310 8660 -60 8710
rect -310 8620 -215 8660
rect -285 8600 -215 8620
rect -155 8620 -60 8660
rect -155 8600 -85 8620
rect -370 8585 -314 8591
rect -370 8525 -366 8585
rect -285 8575 -85 8600
rect -30 8591 0 8779
rect -56 8585 0 8591
rect -314 8525 -56 8545
rect -4 8525 0 8585
rect -370 8515 0 8525
rect 30 8845 400 8855
rect 30 8785 34 8845
rect 86 8825 344 8845
rect 30 8779 86 8785
rect 30 8591 60 8779
rect 115 8770 315 8795
rect 396 8785 400 8845
rect 344 8779 400 8785
rect 115 8750 185 8770
rect 90 8710 185 8750
rect 245 8750 315 8770
rect 245 8710 340 8750
rect 90 8660 340 8710
rect 90 8620 185 8660
rect 115 8600 185 8620
rect 245 8620 340 8660
rect 245 8600 315 8620
rect 30 8585 86 8591
rect 30 8525 34 8585
rect 115 8575 315 8600
rect 370 8591 400 8779
rect 344 8585 400 8591
rect 86 8525 344 8545
rect 396 8525 400 8585
rect 30 8515 400 8525
rect 430 8845 800 8855
rect 430 8785 434 8845
rect 486 8825 744 8845
rect 430 8779 486 8785
rect 430 8591 460 8779
rect 515 8770 715 8795
rect 796 8785 800 8845
rect 744 8779 800 8785
rect 515 8750 585 8770
rect 490 8710 585 8750
rect 645 8750 715 8770
rect 645 8710 740 8750
rect 490 8660 740 8710
rect 490 8620 585 8660
rect 515 8600 585 8620
rect 645 8620 740 8660
rect 645 8600 715 8620
rect 430 8585 486 8591
rect 430 8525 434 8585
rect 515 8575 715 8600
rect 770 8591 800 8779
rect 744 8585 800 8591
rect 486 8525 744 8545
rect 796 8525 800 8585
rect 430 8515 800 8525
rect 830 8845 1200 8855
rect 830 8785 834 8845
rect 886 8825 1144 8845
rect 830 8779 886 8785
rect 830 8591 860 8779
rect 915 8770 1115 8795
rect 1196 8785 1200 8845
rect 1144 8779 1200 8785
rect 915 8750 985 8770
rect 890 8710 985 8750
rect 1045 8750 1115 8770
rect 1045 8710 1140 8750
rect 890 8660 1140 8710
rect 890 8620 985 8660
rect 915 8600 985 8620
rect 1045 8620 1140 8660
rect 1045 8600 1115 8620
rect 830 8585 886 8591
rect 830 8525 834 8585
rect 915 8575 1115 8600
rect 1170 8591 1200 8779
rect 1144 8585 1200 8591
rect 886 8525 1144 8545
rect 1196 8525 1200 8585
rect 830 8515 1200 8525
rect 1230 8845 1600 8855
rect 1230 8785 1234 8845
rect 1286 8825 1544 8845
rect 1230 8779 1286 8785
rect 1230 8591 1260 8779
rect 1315 8770 1515 8795
rect 1596 8785 1600 8845
rect 1544 8779 1600 8785
rect 1315 8750 1385 8770
rect 1290 8710 1385 8750
rect 1445 8750 1515 8770
rect 1445 8710 1540 8750
rect 1290 8660 1540 8710
rect 1290 8620 1385 8660
rect 1315 8600 1385 8620
rect 1445 8620 1540 8660
rect 1445 8600 1515 8620
rect 1230 8585 1286 8591
rect 1230 8525 1234 8585
rect 1315 8575 1515 8600
rect 1570 8591 1600 8779
rect 1544 8585 1600 8591
rect 1286 8525 1544 8545
rect 1596 8525 1600 8585
rect 1230 8515 1600 8525
rect 1630 8845 2000 8855
rect 1630 8785 1634 8845
rect 1686 8825 1944 8845
rect 1630 8779 1686 8785
rect 1630 8591 1660 8779
rect 1715 8770 1915 8795
rect 1996 8785 2000 8845
rect 1944 8779 2000 8785
rect 1715 8750 1785 8770
rect 1690 8710 1785 8750
rect 1845 8750 1915 8770
rect 1845 8710 1940 8750
rect 1690 8660 1940 8710
rect 1690 8620 1785 8660
rect 1715 8600 1785 8620
rect 1845 8620 1940 8660
rect 1845 8600 1915 8620
rect 1630 8585 1686 8591
rect 1630 8525 1634 8585
rect 1715 8575 1915 8600
rect 1970 8591 2000 8779
rect 1944 8585 2000 8591
rect 1686 8525 1944 8545
rect 1996 8525 2000 8585
rect 1630 8515 2000 8525
rect 2030 8845 2400 8855
rect 2030 8785 2034 8845
rect 2086 8825 2344 8845
rect 2030 8779 2086 8785
rect 2030 8591 2060 8779
rect 2115 8770 2315 8795
rect 2396 8785 2400 8845
rect 2344 8779 2400 8785
rect 2115 8750 2185 8770
rect 2090 8710 2185 8750
rect 2245 8750 2315 8770
rect 2245 8710 2340 8750
rect 2090 8660 2340 8710
rect 2090 8620 2185 8660
rect 2115 8600 2185 8620
rect 2245 8620 2340 8660
rect 2245 8600 2315 8620
rect 2030 8585 2086 8591
rect 2030 8525 2034 8585
rect 2115 8575 2315 8600
rect 2370 8591 2400 8779
rect 2344 8585 2400 8591
rect 2086 8525 2344 8545
rect 2396 8525 2400 8585
rect 2030 8515 2400 8525
rect 2430 8845 2800 8855
rect 2430 8785 2434 8845
rect 2486 8825 2744 8845
rect 2430 8779 2486 8785
rect 2430 8591 2460 8779
rect 2515 8770 2715 8795
rect 2796 8785 2800 8845
rect 2744 8779 2800 8785
rect 2515 8750 2585 8770
rect 2490 8710 2585 8750
rect 2645 8750 2715 8770
rect 2645 8710 2740 8750
rect 2490 8660 2740 8710
rect 2490 8620 2585 8660
rect 2515 8600 2585 8620
rect 2645 8620 2740 8660
rect 2645 8600 2715 8620
rect 2430 8585 2486 8591
rect 2430 8525 2434 8585
rect 2515 8575 2715 8600
rect 2770 8591 2800 8779
rect 2744 8585 2800 8591
rect 2486 8525 2744 8545
rect 2796 8525 2800 8585
rect 2430 8515 2800 8525
rect 2830 8845 3200 8855
rect 2830 8785 2834 8845
rect 2886 8825 3144 8845
rect 2830 8779 2886 8785
rect 2830 8591 2860 8779
rect 2915 8770 3115 8795
rect 3196 8785 3200 8845
rect 3144 8779 3200 8785
rect 2915 8750 2985 8770
rect 2890 8710 2985 8750
rect 3045 8750 3115 8770
rect 3045 8710 3140 8750
rect 2890 8660 3140 8710
rect 2890 8620 2985 8660
rect 2915 8600 2985 8620
rect 3045 8620 3140 8660
rect 3045 8600 3115 8620
rect 2830 8585 2886 8591
rect 2830 8525 2834 8585
rect 2915 8575 3115 8600
rect 3170 8591 3200 8779
rect 3144 8585 3200 8591
rect 2886 8525 3144 8545
rect 3196 8525 3200 8585
rect 2830 8515 3200 8525
rect 3230 8845 3600 8855
rect 3230 8785 3234 8845
rect 3286 8825 3544 8845
rect 3230 8779 3286 8785
rect 3230 8591 3260 8779
rect 3315 8770 3515 8795
rect 3596 8785 3600 8845
rect 3544 8779 3600 8785
rect 3315 8750 3385 8770
rect 3290 8710 3385 8750
rect 3445 8750 3515 8770
rect 3445 8710 3540 8750
rect 3290 8660 3540 8710
rect 3290 8620 3385 8660
rect 3315 8600 3385 8620
rect 3445 8620 3540 8660
rect 3445 8600 3515 8620
rect 3230 8585 3286 8591
rect 3230 8525 3234 8585
rect 3315 8575 3515 8600
rect 3570 8591 3600 8779
rect 3544 8585 3600 8591
rect 3286 8525 3544 8545
rect 3596 8525 3600 8585
rect 3230 8515 3600 8525
rect 3630 8845 4000 8855
rect 3630 8785 3634 8845
rect 3686 8825 3944 8845
rect 3630 8779 3686 8785
rect 3630 8591 3660 8779
rect 3715 8770 3915 8795
rect 3996 8785 4000 8845
rect 3944 8779 4000 8785
rect 3715 8750 3785 8770
rect 3690 8710 3785 8750
rect 3845 8750 3915 8770
rect 3845 8710 3940 8750
rect 3690 8660 3940 8710
rect 3690 8620 3785 8660
rect 3715 8600 3785 8620
rect 3845 8620 3940 8660
rect 3845 8600 3915 8620
rect 3630 8585 3686 8591
rect 3630 8525 3634 8585
rect 3715 8575 3915 8600
rect 3970 8591 4000 8779
rect 3944 8585 4000 8591
rect 3686 8525 3944 8545
rect 3996 8525 4000 8585
rect 3630 8515 4000 8525
rect 4030 8845 4400 8855
rect 4030 8785 4034 8845
rect 4086 8825 4344 8845
rect 4030 8779 4086 8785
rect 4030 8591 4060 8779
rect 4115 8770 4315 8795
rect 4396 8785 4400 8845
rect 4344 8779 4400 8785
rect 4115 8750 4185 8770
rect 4090 8710 4185 8750
rect 4245 8750 4315 8770
rect 4245 8710 4340 8750
rect 4090 8660 4340 8710
rect 4090 8620 4185 8660
rect 4115 8600 4185 8620
rect 4245 8620 4340 8660
rect 4245 8600 4315 8620
rect 4030 8585 4086 8591
rect 4030 8525 4034 8585
rect 4115 8575 4315 8600
rect 4370 8591 4400 8779
rect 4344 8585 4400 8591
rect 4086 8525 4344 8545
rect 4396 8525 4400 8585
rect 4030 8515 4400 8525
rect 4430 8845 4800 8855
rect 4430 8785 4434 8845
rect 4486 8825 4744 8845
rect 4430 8779 4486 8785
rect 4430 8591 4460 8779
rect 4515 8770 4715 8795
rect 4796 8785 4800 8845
rect 4744 8779 4800 8785
rect 4515 8750 4585 8770
rect 4490 8710 4585 8750
rect 4645 8750 4715 8770
rect 4645 8710 4740 8750
rect 4490 8660 4740 8710
rect 4490 8620 4585 8660
rect 4515 8600 4585 8620
rect 4645 8620 4740 8660
rect 4645 8600 4715 8620
rect 4430 8585 4486 8591
rect 4430 8525 4434 8585
rect 4515 8575 4715 8600
rect 4770 8591 4800 8779
rect 4744 8585 4800 8591
rect 4486 8525 4744 8545
rect 4796 8525 4800 8585
rect 4430 8515 4800 8525
rect 4830 8845 5200 8855
rect 4830 8785 4834 8845
rect 4886 8825 5144 8845
rect 4830 8779 4886 8785
rect 4830 8591 4860 8779
rect 4915 8770 5115 8795
rect 5196 8785 5200 8845
rect 5144 8779 5200 8785
rect 4915 8750 4985 8770
rect 4890 8710 4985 8750
rect 5045 8750 5115 8770
rect 5045 8710 5140 8750
rect 4890 8660 5140 8710
rect 4890 8620 4985 8660
rect 4915 8600 4985 8620
rect 5045 8620 5140 8660
rect 5045 8600 5115 8620
rect 4830 8585 4886 8591
rect 4830 8525 4834 8585
rect 4915 8575 5115 8600
rect 5170 8591 5200 8779
rect 5144 8585 5200 8591
rect 4886 8525 5144 8545
rect 5196 8525 5200 8585
rect 4830 8515 5200 8525
rect 5230 8845 5600 8855
rect 5230 8785 5234 8845
rect 5286 8825 5544 8845
rect 5230 8779 5286 8785
rect 5230 8591 5260 8779
rect 5315 8770 5515 8795
rect 5596 8785 5600 8845
rect 5544 8779 5600 8785
rect 5315 8750 5385 8770
rect 5290 8710 5385 8750
rect 5445 8750 5515 8770
rect 5445 8710 5540 8750
rect 5290 8660 5540 8710
rect 5290 8620 5385 8660
rect 5315 8600 5385 8620
rect 5445 8620 5540 8660
rect 5445 8600 5515 8620
rect 5230 8585 5286 8591
rect 5230 8525 5234 8585
rect 5315 8575 5515 8600
rect 5570 8591 5600 8779
rect 5544 8585 5600 8591
rect 5286 8525 5544 8545
rect 5596 8525 5600 8585
rect 5230 8515 5600 8525
rect 5630 8845 6000 8855
rect 5630 8785 5634 8845
rect 5686 8825 5944 8845
rect 5630 8779 5686 8785
rect 5630 8591 5660 8779
rect 5715 8770 5915 8795
rect 5996 8785 6000 8845
rect 5944 8779 6000 8785
rect 5715 8750 5785 8770
rect 5690 8710 5785 8750
rect 5845 8750 5915 8770
rect 5845 8710 5940 8750
rect 5690 8660 5940 8710
rect 5690 8620 5785 8660
rect 5715 8600 5785 8620
rect 5845 8620 5940 8660
rect 5845 8600 5915 8620
rect 5630 8585 5686 8591
rect 5630 8525 5634 8585
rect 5715 8575 5915 8600
rect 5970 8591 6000 8779
rect 5944 8585 6000 8591
rect 5686 8525 5944 8545
rect 5996 8525 6000 8585
rect 5630 8515 6000 8525
rect 6030 8845 6400 8855
rect 6030 8785 6034 8845
rect 6086 8825 6344 8845
rect 6030 8779 6086 8785
rect 6030 8591 6060 8779
rect 6115 8770 6315 8795
rect 6396 8785 6400 8845
rect 6344 8779 6400 8785
rect 6115 8750 6185 8770
rect 6090 8710 6185 8750
rect 6245 8750 6315 8770
rect 6245 8710 6340 8750
rect 6090 8660 6340 8710
rect 6090 8620 6185 8660
rect 6115 8600 6185 8620
rect 6245 8620 6340 8660
rect 6245 8600 6315 8620
rect 6030 8585 6086 8591
rect 6030 8525 6034 8585
rect 6115 8575 6315 8600
rect 6370 8591 6400 8779
rect 6344 8585 6400 8591
rect 6086 8525 6344 8545
rect 6396 8525 6400 8585
rect 6030 8515 6400 8525
rect 6430 8845 6800 8855
rect 6430 8785 6434 8845
rect 6486 8825 6744 8845
rect 6430 8779 6486 8785
rect 6430 8591 6460 8779
rect 6515 8770 6715 8795
rect 6796 8785 6800 8845
rect 6744 8779 6800 8785
rect 6515 8750 6585 8770
rect 6490 8710 6585 8750
rect 6645 8750 6715 8770
rect 6645 8710 6740 8750
rect 6490 8660 6740 8710
rect 6490 8620 6585 8660
rect 6515 8600 6585 8620
rect 6645 8620 6740 8660
rect 6645 8600 6715 8620
rect 6430 8585 6486 8591
rect 6430 8525 6434 8585
rect 6515 8575 6715 8600
rect 6770 8591 6800 8779
rect 6744 8585 6800 8591
rect 6486 8525 6744 8545
rect 6796 8525 6800 8585
rect 6430 8515 6800 8525
rect 6830 8845 7200 8855
rect 6830 8785 6834 8845
rect 6886 8825 7144 8845
rect 6830 8779 6886 8785
rect 6830 8591 6860 8779
rect 6915 8770 7115 8795
rect 7196 8785 7200 8845
rect 7144 8779 7200 8785
rect 6915 8750 6985 8770
rect 6890 8710 6985 8750
rect 7045 8750 7115 8770
rect 7045 8710 7140 8750
rect 6890 8660 7140 8710
rect 6890 8620 6985 8660
rect 6915 8600 6985 8620
rect 7045 8620 7140 8660
rect 7045 8600 7115 8620
rect 6830 8585 6886 8591
rect 6830 8525 6834 8585
rect 6915 8575 7115 8600
rect 7170 8591 7200 8779
rect 7144 8585 7200 8591
rect 6886 8525 7144 8545
rect 7196 8525 7200 8585
rect 6830 8515 7200 8525
rect 7230 8845 7600 8855
rect 7230 8785 7234 8845
rect 7286 8825 7544 8845
rect 7230 8779 7286 8785
rect 7230 8591 7260 8779
rect 7315 8770 7515 8795
rect 7596 8785 7600 8845
rect 7544 8779 7600 8785
rect 7315 8750 7385 8770
rect 7290 8710 7385 8750
rect 7445 8750 7515 8770
rect 7445 8710 7540 8750
rect 7290 8660 7540 8710
rect 7290 8620 7385 8660
rect 7315 8600 7385 8620
rect 7445 8620 7540 8660
rect 7445 8600 7515 8620
rect 7230 8585 7286 8591
rect 7230 8525 7234 8585
rect 7315 8575 7515 8600
rect 7570 8591 7600 8779
rect 7544 8585 7600 8591
rect 7286 8525 7544 8545
rect 7596 8525 7600 8585
rect 7230 8515 7600 8525
rect 7630 8845 8000 8855
rect 7630 8785 7634 8845
rect 7686 8825 7944 8845
rect 7630 8779 7686 8785
rect 7630 8591 7660 8779
rect 7715 8770 7915 8795
rect 7996 8785 8000 8845
rect 7944 8779 8000 8785
rect 7715 8750 7785 8770
rect 7690 8710 7785 8750
rect 7845 8750 7915 8770
rect 7845 8710 7940 8750
rect 7690 8660 7940 8710
rect 7690 8620 7785 8660
rect 7715 8600 7785 8620
rect 7845 8620 7940 8660
rect 7845 8600 7915 8620
rect 7630 8585 7686 8591
rect 7630 8525 7634 8585
rect 7715 8575 7915 8600
rect 7970 8591 8000 8779
rect 7944 8585 8000 8591
rect 7686 8525 7944 8545
rect 7996 8525 8000 8585
rect 7630 8515 8000 8525
rect 8030 8845 8400 8855
rect 8030 8785 8034 8845
rect 8086 8825 8344 8845
rect 8030 8779 8086 8785
rect 8030 8591 8060 8779
rect 8115 8770 8315 8795
rect 8396 8785 8400 8845
rect 8344 8779 8400 8785
rect 8115 8750 8185 8770
rect 8090 8710 8185 8750
rect 8245 8750 8315 8770
rect 8245 8710 8340 8750
rect 8090 8660 8340 8710
rect 8090 8620 8185 8660
rect 8115 8600 8185 8620
rect 8245 8620 8340 8660
rect 8245 8600 8315 8620
rect 8030 8585 8086 8591
rect 8030 8525 8034 8585
rect 8115 8575 8315 8600
rect 8370 8591 8400 8779
rect 8344 8585 8400 8591
rect 8086 8525 8344 8545
rect 8396 8525 8400 8585
rect 8030 8515 8400 8525
rect 8430 8845 8800 8855
rect 8430 8785 8434 8845
rect 8486 8825 8744 8845
rect 8430 8779 8486 8785
rect 8430 8591 8460 8779
rect 8515 8770 8715 8795
rect 8796 8785 8800 8845
rect 8744 8779 8800 8785
rect 8515 8750 8585 8770
rect 8490 8710 8585 8750
rect 8645 8750 8715 8770
rect 8645 8710 8740 8750
rect 8490 8660 8740 8710
rect 8490 8620 8585 8660
rect 8515 8600 8585 8620
rect 8645 8620 8740 8660
rect 8645 8600 8715 8620
rect 8430 8585 8486 8591
rect 8430 8525 8434 8585
rect 8515 8575 8715 8600
rect 8770 8591 8800 8779
rect 8744 8585 8800 8591
rect 8486 8525 8744 8545
rect 8796 8525 8800 8585
rect 8430 8515 8800 8525
rect 8830 8845 9200 8855
rect 8830 8785 8834 8845
rect 8886 8825 9144 8845
rect 8830 8779 8886 8785
rect 8830 8591 8860 8779
rect 8915 8770 9115 8795
rect 9196 8785 9200 8845
rect 9144 8779 9200 8785
rect 8915 8750 8985 8770
rect 8890 8710 8985 8750
rect 9045 8750 9115 8770
rect 9045 8710 9140 8750
rect 8890 8660 9140 8710
rect 8890 8620 8985 8660
rect 8915 8600 8985 8620
rect 9045 8620 9140 8660
rect 9045 8600 9115 8620
rect 8830 8585 8886 8591
rect 8830 8525 8834 8585
rect 8915 8575 9115 8600
rect 9170 8591 9200 8779
rect 9144 8585 9200 8591
rect 8886 8525 9144 8545
rect 9196 8525 9200 8585
rect 8830 8515 9200 8525
rect 9230 8845 9600 8855
rect 9230 8785 9234 8845
rect 9286 8825 9544 8845
rect 9230 8779 9286 8785
rect 9230 8591 9260 8779
rect 9315 8770 9515 8795
rect 9596 8785 9600 8845
rect 9544 8779 9600 8785
rect 9315 8750 9385 8770
rect 9290 8710 9385 8750
rect 9445 8750 9515 8770
rect 9445 8710 9540 8750
rect 9290 8660 9540 8710
rect 9290 8620 9385 8660
rect 9315 8600 9385 8620
rect 9445 8620 9540 8660
rect 9445 8600 9515 8620
rect 9230 8585 9286 8591
rect 9230 8525 9234 8585
rect 9315 8575 9515 8600
rect 9570 8591 9600 8779
rect 9544 8585 9600 8591
rect 9286 8525 9544 8545
rect 9596 8525 9600 8585
rect 9230 8515 9600 8525
rect 9630 8845 10000 8855
rect 9630 8785 9634 8845
rect 9686 8825 9944 8845
rect 9630 8779 9686 8785
rect 9630 8591 9660 8779
rect 9715 8770 9915 8795
rect 9996 8785 10000 8845
rect 9944 8779 10000 8785
rect 9715 8750 9785 8770
rect 9690 8710 9785 8750
rect 9845 8750 9915 8770
rect 9845 8710 9940 8750
rect 9690 8660 9940 8710
rect 9690 8620 9785 8660
rect 9715 8600 9785 8620
rect 9845 8620 9940 8660
rect 9845 8600 9915 8620
rect 9630 8585 9686 8591
rect 9630 8525 9634 8585
rect 9715 8575 9915 8600
rect 9970 8591 10000 8779
rect 9944 8585 10000 8591
rect 9686 8525 9944 8545
rect 9996 8525 10000 8585
rect 9630 8515 10000 8525
rect 10030 8845 10400 8855
rect 10030 8785 10034 8845
rect 10086 8825 10344 8845
rect 10030 8779 10086 8785
rect 10030 8591 10060 8779
rect 10115 8770 10315 8795
rect 10396 8785 10400 8845
rect 10344 8779 10400 8785
rect 10115 8750 10185 8770
rect 10090 8710 10185 8750
rect 10245 8750 10315 8770
rect 10245 8710 10340 8750
rect 10090 8660 10340 8710
rect 10090 8620 10185 8660
rect 10115 8600 10185 8620
rect 10245 8620 10340 8660
rect 10245 8600 10315 8620
rect 10030 8585 10086 8591
rect 10030 8525 10034 8585
rect 10115 8575 10315 8600
rect 10370 8591 10400 8779
rect 10344 8585 10400 8591
rect 10086 8525 10344 8545
rect 10396 8525 10400 8585
rect 10030 8515 10400 8525
rect 10430 8845 10800 8855
rect 10430 8785 10434 8845
rect 10486 8825 10744 8845
rect 10430 8779 10486 8785
rect 10430 8591 10460 8779
rect 10515 8770 10715 8795
rect 10796 8785 10800 8845
rect 10744 8779 10800 8785
rect 10515 8750 10585 8770
rect 10490 8710 10585 8750
rect 10645 8750 10715 8770
rect 10645 8710 10740 8750
rect 10490 8660 10740 8710
rect 10490 8620 10585 8660
rect 10515 8600 10585 8620
rect 10645 8620 10740 8660
rect 10645 8600 10715 8620
rect 10430 8585 10486 8591
rect 10430 8525 10434 8585
rect 10515 8575 10715 8600
rect 10770 8591 10800 8779
rect 10744 8585 10800 8591
rect 10486 8525 10744 8545
rect 10796 8525 10800 8585
rect 10430 8515 10800 8525
rect 10830 8845 11200 8855
rect 10830 8785 10834 8845
rect 10886 8825 11144 8845
rect 10830 8779 10886 8785
rect 10830 8591 10860 8779
rect 10915 8770 11115 8795
rect 11196 8785 11200 8845
rect 11144 8779 11200 8785
rect 10915 8750 10985 8770
rect 10890 8710 10985 8750
rect 11045 8750 11115 8770
rect 11045 8710 11140 8750
rect 10890 8660 11140 8710
rect 10890 8620 10985 8660
rect 10915 8600 10985 8620
rect 11045 8620 11140 8660
rect 11045 8600 11115 8620
rect 10830 8585 10886 8591
rect 10830 8525 10834 8585
rect 10915 8575 11115 8600
rect 11170 8591 11200 8779
rect 11144 8585 11200 8591
rect 10886 8525 11144 8545
rect 11196 8525 11200 8585
rect 10830 8515 11200 8525
rect 11230 8845 11600 8855
rect 11230 8785 11234 8845
rect 11286 8825 11544 8845
rect 11230 8779 11286 8785
rect 11230 8591 11260 8779
rect 11315 8770 11515 8795
rect 11596 8785 11600 8845
rect 11544 8779 11600 8785
rect 11315 8750 11385 8770
rect 11290 8710 11385 8750
rect 11445 8750 11515 8770
rect 11445 8710 11540 8750
rect 11290 8660 11540 8710
rect 11290 8620 11385 8660
rect 11315 8600 11385 8620
rect 11445 8620 11540 8660
rect 11445 8600 11515 8620
rect 11230 8585 11286 8591
rect 11230 8525 11234 8585
rect 11315 8575 11515 8600
rect 11570 8591 11600 8779
rect 11544 8585 11600 8591
rect 11286 8525 11544 8545
rect 11596 8525 11600 8585
rect 11230 8515 11600 8525
rect 11630 8845 12000 8855
rect 11630 8785 11634 8845
rect 11686 8825 11944 8845
rect 11630 8779 11686 8785
rect 11630 8591 11660 8779
rect 11715 8770 11915 8795
rect 11996 8785 12000 8845
rect 11944 8779 12000 8785
rect 11715 8750 11785 8770
rect 11690 8710 11785 8750
rect 11845 8750 11915 8770
rect 11845 8710 11940 8750
rect 11690 8660 11940 8710
rect 11690 8620 11785 8660
rect 11715 8600 11785 8620
rect 11845 8620 11940 8660
rect 11845 8600 11915 8620
rect 11630 8585 11686 8591
rect 11630 8525 11634 8585
rect 11715 8575 11915 8600
rect 11970 8591 12000 8779
rect 11944 8585 12000 8591
rect 11686 8525 11944 8545
rect 11996 8525 12000 8585
rect 11630 8515 12000 8525
rect 12030 8845 12400 8855
rect 12030 8785 12034 8845
rect 12086 8825 12344 8845
rect 12030 8779 12086 8785
rect 12030 8591 12060 8779
rect 12115 8770 12315 8795
rect 12396 8785 12400 8845
rect 12344 8779 12400 8785
rect 12115 8750 12185 8770
rect 12090 8710 12185 8750
rect 12245 8750 12315 8770
rect 12245 8710 12340 8750
rect 12090 8660 12340 8710
rect 12090 8620 12185 8660
rect 12115 8600 12185 8620
rect 12245 8620 12340 8660
rect 12245 8600 12315 8620
rect 12030 8585 12086 8591
rect 12030 8525 12034 8585
rect 12115 8575 12315 8600
rect 12370 8591 12400 8779
rect 12344 8585 12400 8591
rect 12086 8525 12344 8545
rect 12396 8525 12400 8585
rect 12030 8515 12400 8525
rect 12430 8845 12800 8855
rect 12430 8785 12434 8845
rect 12486 8825 12744 8845
rect 12430 8779 12486 8785
rect 12430 8591 12460 8779
rect 12515 8770 12715 8795
rect 12796 8785 12800 8845
rect 12744 8779 12800 8785
rect 12515 8750 12585 8770
rect 12490 8710 12585 8750
rect 12645 8750 12715 8770
rect 12645 8710 12740 8750
rect 12490 8660 12740 8710
rect 12490 8620 12585 8660
rect 12515 8600 12585 8620
rect 12645 8620 12740 8660
rect 12645 8600 12715 8620
rect 12430 8585 12486 8591
rect 12430 8525 12434 8585
rect 12515 8575 12715 8600
rect 12770 8591 12800 8779
rect 12744 8585 12800 8591
rect 12486 8525 12744 8545
rect 12796 8525 12800 8585
rect 12430 8515 12800 8525
rect 12830 8845 13200 8855
rect 12830 8785 12834 8845
rect 12886 8825 13144 8845
rect 12830 8779 12886 8785
rect 12830 8591 12860 8779
rect 12915 8770 13115 8795
rect 13196 8785 13200 8845
rect 13144 8779 13200 8785
rect 12915 8750 12985 8770
rect 12890 8710 12985 8750
rect 13045 8750 13115 8770
rect 13045 8710 13140 8750
rect 12890 8660 13140 8710
rect 12890 8620 12985 8660
rect 12915 8600 12985 8620
rect 13045 8620 13140 8660
rect 13045 8600 13115 8620
rect 12830 8585 12886 8591
rect 12830 8525 12834 8585
rect 12915 8575 13115 8600
rect 13170 8591 13200 8779
rect 13144 8585 13200 8591
rect 12886 8525 13144 8545
rect 13196 8525 13200 8585
rect 12830 8515 13200 8525
rect -370 8475 0 8485
rect -370 8415 -366 8475
rect -314 8455 -56 8475
rect -370 8409 -314 8415
rect -370 8221 -340 8409
rect -285 8400 -85 8425
rect -4 8415 0 8475
rect -56 8409 0 8415
rect -285 8380 -215 8400
rect -310 8340 -215 8380
rect -155 8380 -85 8400
rect -155 8340 -60 8380
rect -310 8290 -60 8340
rect -310 8250 -215 8290
rect -285 8230 -215 8250
rect -155 8250 -60 8290
rect -155 8230 -85 8250
rect -370 8215 -314 8221
rect -370 8155 -366 8215
rect -285 8205 -85 8230
rect -30 8221 0 8409
rect -56 8215 0 8221
rect -314 8155 -56 8175
rect -4 8155 0 8215
rect -370 8145 0 8155
rect 30 8475 400 8485
rect 30 8415 34 8475
rect 86 8455 344 8475
rect 30 8409 86 8415
rect 30 8221 60 8409
rect 115 8400 315 8425
rect 396 8415 400 8475
rect 344 8409 400 8415
rect 115 8380 185 8400
rect 90 8340 185 8380
rect 245 8380 315 8400
rect 245 8340 340 8380
rect 90 8290 340 8340
rect 90 8250 185 8290
rect 115 8230 185 8250
rect 245 8250 340 8290
rect 245 8230 315 8250
rect 30 8215 86 8221
rect 30 8155 34 8215
rect 115 8205 315 8230
rect 370 8221 400 8409
rect 344 8215 400 8221
rect 86 8155 344 8175
rect 396 8155 400 8215
rect 30 8145 400 8155
rect 430 8475 800 8485
rect 430 8415 434 8475
rect 486 8455 744 8475
rect 430 8409 486 8415
rect 430 8221 460 8409
rect 515 8400 715 8425
rect 796 8415 800 8475
rect 744 8409 800 8415
rect 515 8380 585 8400
rect 490 8340 585 8380
rect 645 8380 715 8400
rect 645 8340 740 8380
rect 490 8290 740 8340
rect 490 8250 585 8290
rect 515 8230 585 8250
rect 645 8250 740 8290
rect 645 8230 715 8250
rect 430 8215 486 8221
rect 430 8155 434 8215
rect 515 8205 715 8230
rect 770 8221 800 8409
rect 744 8215 800 8221
rect 486 8155 744 8175
rect 796 8155 800 8215
rect 430 8145 800 8155
rect 830 8475 1200 8485
rect 830 8415 834 8475
rect 886 8455 1144 8475
rect 830 8409 886 8415
rect 830 8221 860 8409
rect 915 8400 1115 8425
rect 1196 8415 1200 8475
rect 1144 8409 1200 8415
rect 915 8380 985 8400
rect 890 8340 985 8380
rect 1045 8380 1115 8400
rect 1045 8340 1140 8380
rect 890 8290 1140 8340
rect 890 8250 985 8290
rect 915 8230 985 8250
rect 1045 8250 1140 8290
rect 1045 8230 1115 8250
rect 830 8215 886 8221
rect 830 8155 834 8215
rect 915 8205 1115 8230
rect 1170 8221 1200 8409
rect 1144 8215 1200 8221
rect 886 8155 1144 8175
rect 1196 8155 1200 8215
rect 830 8145 1200 8155
rect 1230 8475 1600 8485
rect 1230 8415 1234 8475
rect 1286 8455 1544 8475
rect 1230 8409 1286 8415
rect 1230 8221 1260 8409
rect 1315 8400 1515 8425
rect 1596 8415 1600 8475
rect 1544 8409 1600 8415
rect 1315 8380 1385 8400
rect 1290 8340 1385 8380
rect 1445 8380 1515 8400
rect 1445 8340 1540 8380
rect 1290 8290 1540 8340
rect 1290 8250 1385 8290
rect 1315 8230 1385 8250
rect 1445 8250 1540 8290
rect 1445 8230 1515 8250
rect 1230 8215 1286 8221
rect 1230 8155 1234 8215
rect 1315 8205 1515 8230
rect 1570 8221 1600 8409
rect 1544 8215 1600 8221
rect 1286 8155 1544 8175
rect 1596 8155 1600 8215
rect 1230 8145 1600 8155
rect 1630 8475 2000 8485
rect 1630 8415 1634 8475
rect 1686 8455 1944 8475
rect 1630 8409 1686 8415
rect 1630 8221 1660 8409
rect 1715 8400 1915 8425
rect 1996 8415 2000 8475
rect 1944 8409 2000 8415
rect 1715 8380 1785 8400
rect 1690 8340 1785 8380
rect 1845 8380 1915 8400
rect 1845 8340 1940 8380
rect 1690 8290 1940 8340
rect 1690 8250 1785 8290
rect 1715 8230 1785 8250
rect 1845 8250 1940 8290
rect 1845 8230 1915 8250
rect 1630 8215 1686 8221
rect 1630 8155 1634 8215
rect 1715 8205 1915 8230
rect 1970 8221 2000 8409
rect 1944 8215 2000 8221
rect 1686 8155 1944 8175
rect 1996 8155 2000 8215
rect 1630 8145 2000 8155
rect 2030 8475 2400 8485
rect 2030 8415 2034 8475
rect 2086 8455 2344 8475
rect 2030 8409 2086 8415
rect 2030 8221 2060 8409
rect 2115 8400 2315 8425
rect 2396 8415 2400 8475
rect 2344 8409 2400 8415
rect 2115 8380 2185 8400
rect 2090 8340 2185 8380
rect 2245 8380 2315 8400
rect 2245 8340 2340 8380
rect 2090 8290 2340 8340
rect 2090 8250 2185 8290
rect 2115 8230 2185 8250
rect 2245 8250 2340 8290
rect 2245 8230 2315 8250
rect 2030 8215 2086 8221
rect 2030 8155 2034 8215
rect 2115 8205 2315 8230
rect 2370 8221 2400 8409
rect 2344 8215 2400 8221
rect 2086 8155 2344 8175
rect 2396 8155 2400 8215
rect 2030 8145 2400 8155
rect 2430 8475 2800 8485
rect 2430 8415 2434 8475
rect 2486 8455 2744 8475
rect 2430 8409 2486 8415
rect 2430 8221 2460 8409
rect 2515 8400 2715 8425
rect 2796 8415 2800 8475
rect 2744 8409 2800 8415
rect 2515 8380 2585 8400
rect 2490 8340 2585 8380
rect 2645 8380 2715 8400
rect 2645 8340 2740 8380
rect 2490 8290 2740 8340
rect 2490 8250 2585 8290
rect 2515 8230 2585 8250
rect 2645 8250 2740 8290
rect 2645 8230 2715 8250
rect 2430 8215 2486 8221
rect 2430 8155 2434 8215
rect 2515 8205 2715 8230
rect 2770 8221 2800 8409
rect 2744 8215 2800 8221
rect 2486 8155 2744 8175
rect 2796 8155 2800 8215
rect 2430 8145 2800 8155
rect 2830 8475 3200 8485
rect 2830 8415 2834 8475
rect 2886 8455 3144 8475
rect 2830 8409 2886 8415
rect 2830 8221 2860 8409
rect 2915 8400 3115 8425
rect 3196 8415 3200 8475
rect 3144 8409 3200 8415
rect 2915 8380 2985 8400
rect 2890 8340 2985 8380
rect 3045 8380 3115 8400
rect 3045 8340 3140 8380
rect 2890 8290 3140 8340
rect 2890 8250 2985 8290
rect 2915 8230 2985 8250
rect 3045 8250 3140 8290
rect 3045 8230 3115 8250
rect 2830 8215 2886 8221
rect 2830 8155 2834 8215
rect 2915 8205 3115 8230
rect 3170 8221 3200 8409
rect 3144 8215 3200 8221
rect 2886 8155 3144 8175
rect 3196 8155 3200 8215
rect 2830 8145 3200 8155
rect 3230 8475 3600 8485
rect 3230 8415 3234 8475
rect 3286 8455 3544 8475
rect 3230 8409 3286 8415
rect 3230 8221 3260 8409
rect 3315 8400 3515 8425
rect 3596 8415 3600 8475
rect 3544 8409 3600 8415
rect 3315 8380 3385 8400
rect 3290 8340 3385 8380
rect 3445 8380 3515 8400
rect 3445 8340 3540 8380
rect 3290 8290 3540 8340
rect 3290 8250 3385 8290
rect 3315 8230 3385 8250
rect 3445 8250 3540 8290
rect 3445 8230 3515 8250
rect 3230 8215 3286 8221
rect 3230 8155 3234 8215
rect 3315 8205 3515 8230
rect 3570 8221 3600 8409
rect 3544 8215 3600 8221
rect 3286 8155 3544 8175
rect 3596 8155 3600 8215
rect 3230 8145 3600 8155
rect 3630 8475 4000 8485
rect 3630 8415 3634 8475
rect 3686 8455 3944 8475
rect 3630 8409 3686 8415
rect 3630 8221 3660 8409
rect 3715 8400 3915 8425
rect 3996 8415 4000 8475
rect 3944 8409 4000 8415
rect 3715 8380 3785 8400
rect 3690 8340 3785 8380
rect 3845 8380 3915 8400
rect 3845 8340 3940 8380
rect 3690 8290 3940 8340
rect 3690 8250 3785 8290
rect 3715 8230 3785 8250
rect 3845 8250 3940 8290
rect 3845 8230 3915 8250
rect 3630 8215 3686 8221
rect 3630 8155 3634 8215
rect 3715 8205 3915 8230
rect 3970 8221 4000 8409
rect 3944 8215 4000 8221
rect 3686 8155 3944 8175
rect 3996 8155 4000 8215
rect 3630 8145 4000 8155
rect 4030 8475 4400 8485
rect 4030 8415 4034 8475
rect 4086 8455 4344 8475
rect 4030 8409 4086 8415
rect 4030 8221 4060 8409
rect 4115 8400 4315 8425
rect 4396 8415 4400 8475
rect 4344 8409 4400 8415
rect 4115 8380 4185 8400
rect 4090 8340 4185 8380
rect 4245 8380 4315 8400
rect 4245 8340 4340 8380
rect 4090 8290 4340 8340
rect 4090 8250 4185 8290
rect 4115 8230 4185 8250
rect 4245 8250 4340 8290
rect 4245 8230 4315 8250
rect 4030 8215 4086 8221
rect 4030 8155 4034 8215
rect 4115 8205 4315 8230
rect 4370 8221 4400 8409
rect 4344 8215 4400 8221
rect 4086 8155 4344 8175
rect 4396 8155 4400 8215
rect 4030 8145 4400 8155
rect 4430 8475 4800 8485
rect 4430 8415 4434 8475
rect 4486 8455 4744 8475
rect 4430 8409 4486 8415
rect 4430 8221 4460 8409
rect 4515 8400 4715 8425
rect 4796 8415 4800 8475
rect 4744 8409 4800 8415
rect 4515 8380 4585 8400
rect 4490 8340 4585 8380
rect 4645 8380 4715 8400
rect 4645 8340 4740 8380
rect 4490 8290 4740 8340
rect 4490 8250 4585 8290
rect 4515 8230 4585 8250
rect 4645 8250 4740 8290
rect 4645 8230 4715 8250
rect 4430 8215 4486 8221
rect 4430 8155 4434 8215
rect 4515 8205 4715 8230
rect 4770 8221 4800 8409
rect 4744 8215 4800 8221
rect 4486 8155 4744 8175
rect 4796 8155 4800 8215
rect 4430 8145 4800 8155
rect 4830 8475 5200 8485
rect 4830 8415 4834 8475
rect 4886 8455 5144 8475
rect 4830 8409 4886 8415
rect 4830 8221 4860 8409
rect 4915 8400 5115 8425
rect 5196 8415 5200 8475
rect 5144 8409 5200 8415
rect 4915 8380 4985 8400
rect 4890 8340 4985 8380
rect 5045 8380 5115 8400
rect 5045 8340 5140 8380
rect 4890 8290 5140 8340
rect 4890 8250 4985 8290
rect 4915 8230 4985 8250
rect 5045 8250 5140 8290
rect 5045 8230 5115 8250
rect 4830 8215 4886 8221
rect 4830 8155 4834 8215
rect 4915 8205 5115 8230
rect 5170 8221 5200 8409
rect 5144 8215 5200 8221
rect 4886 8155 5144 8175
rect 5196 8155 5200 8215
rect 4830 8145 5200 8155
rect 5230 8475 5600 8485
rect 5230 8415 5234 8475
rect 5286 8455 5544 8475
rect 5230 8409 5286 8415
rect 5230 8221 5260 8409
rect 5315 8400 5515 8425
rect 5596 8415 5600 8475
rect 5544 8409 5600 8415
rect 5315 8380 5385 8400
rect 5290 8340 5385 8380
rect 5445 8380 5515 8400
rect 5445 8340 5540 8380
rect 5290 8290 5540 8340
rect 5290 8250 5385 8290
rect 5315 8230 5385 8250
rect 5445 8250 5540 8290
rect 5445 8230 5515 8250
rect 5230 8215 5286 8221
rect 5230 8155 5234 8215
rect 5315 8205 5515 8230
rect 5570 8221 5600 8409
rect 5544 8215 5600 8221
rect 5286 8155 5544 8175
rect 5596 8155 5600 8215
rect 5230 8145 5600 8155
rect 5630 8475 6000 8485
rect 5630 8415 5634 8475
rect 5686 8455 5944 8475
rect 5630 8409 5686 8415
rect 5630 8221 5660 8409
rect 5715 8400 5915 8425
rect 5996 8415 6000 8475
rect 5944 8409 6000 8415
rect 5715 8380 5785 8400
rect 5690 8340 5785 8380
rect 5845 8380 5915 8400
rect 5845 8340 5940 8380
rect 5690 8290 5940 8340
rect 5690 8250 5785 8290
rect 5715 8230 5785 8250
rect 5845 8250 5940 8290
rect 5845 8230 5915 8250
rect 5630 8215 5686 8221
rect 5630 8155 5634 8215
rect 5715 8205 5915 8230
rect 5970 8221 6000 8409
rect 5944 8215 6000 8221
rect 5686 8155 5944 8175
rect 5996 8155 6000 8215
rect 5630 8145 6000 8155
rect 6030 8475 6400 8485
rect 6030 8415 6034 8475
rect 6086 8455 6344 8475
rect 6030 8409 6086 8415
rect 6030 8221 6060 8409
rect 6115 8400 6315 8425
rect 6396 8415 6400 8475
rect 6344 8409 6400 8415
rect 6115 8380 6185 8400
rect 6090 8340 6185 8380
rect 6245 8380 6315 8400
rect 6245 8340 6340 8380
rect 6090 8290 6340 8340
rect 6090 8250 6185 8290
rect 6115 8230 6185 8250
rect 6245 8250 6340 8290
rect 6245 8230 6315 8250
rect 6030 8215 6086 8221
rect 6030 8155 6034 8215
rect 6115 8205 6315 8230
rect 6370 8221 6400 8409
rect 6344 8215 6400 8221
rect 6086 8155 6344 8175
rect 6396 8155 6400 8215
rect 6030 8145 6400 8155
rect 6430 8475 6800 8485
rect 6430 8415 6434 8475
rect 6486 8455 6744 8475
rect 6430 8409 6486 8415
rect 6430 8221 6460 8409
rect 6515 8400 6715 8425
rect 6796 8415 6800 8475
rect 6744 8409 6800 8415
rect 6515 8380 6585 8400
rect 6490 8340 6585 8380
rect 6645 8380 6715 8400
rect 6645 8340 6740 8380
rect 6490 8290 6740 8340
rect 6490 8250 6585 8290
rect 6515 8230 6585 8250
rect 6645 8250 6740 8290
rect 6645 8230 6715 8250
rect 6430 8215 6486 8221
rect 6430 8155 6434 8215
rect 6515 8205 6715 8230
rect 6770 8221 6800 8409
rect 6744 8215 6800 8221
rect 6486 8155 6744 8175
rect 6796 8155 6800 8215
rect 6430 8145 6800 8155
rect 6830 8475 7200 8485
rect 6830 8415 6834 8475
rect 6886 8455 7144 8475
rect 6830 8409 6886 8415
rect 6830 8221 6860 8409
rect 6915 8400 7115 8425
rect 7196 8415 7200 8475
rect 7144 8409 7200 8415
rect 6915 8380 6985 8400
rect 6890 8340 6985 8380
rect 7045 8380 7115 8400
rect 7045 8340 7140 8380
rect 6890 8290 7140 8340
rect 6890 8250 6985 8290
rect 6915 8230 6985 8250
rect 7045 8250 7140 8290
rect 7045 8230 7115 8250
rect 6830 8215 6886 8221
rect 6830 8155 6834 8215
rect 6915 8205 7115 8230
rect 7170 8221 7200 8409
rect 7144 8215 7200 8221
rect 6886 8155 7144 8175
rect 7196 8155 7200 8215
rect 6830 8145 7200 8155
rect 7230 8475 7600 8485
rect 7230 8415 7234 8475
rect 7286 8455 7544 8475
rect 7230 8409 7286 8415
rect 7230 8221 7260 8409
rect 7315 8400 7515 8425
rect 7596 8415 7600 8475
rect 7544 8409 7600 8415
rect 7315 8380 7385 8400
rect 7290 8340 7385 8380
rect 7445 8380 7515 8400
rect 7445 8340 7540 8380
rect 7290 8290 7540 8340
rect 7290 8250 7385 8290
rect 7315 8230 7385 8250
rect 7445 8250 7540 8290
rect 7445 8230 7515 8250
rect 7230 8215 7286 8221
rect 7230 8155 7234 8215
rect 7315 8205 7515 8230
rect 7570 8221 7600 8409
rect 7544 8215 7600 8221
rect 7286 8155 7544 8175
rect 7596 8155 7600 8215
rect 7230 8145 7600 8155
rect 7630 8475 8000 8485
rect 7630 8415 7634 8475
rect 7686 8455 7944 8475
rect 7630 8409 7686 8415
rect 7630 8221 7660 8409
rect 7715 8400 7915 8425
rect 7996 8415 8000 8475
rect 7944 8409 8000 8415
rect 7715 8380 7785 8400
rect 7690 8340 7785 8380
rect 7845 8380 7915 8400
rect 7845 8340 7940 8380
rect 7690 8290 7940 8340
rect 7690 8250 7785 8290
rect 7715 8230 7785 8250
rect 7845 8250 7940 8290
rect 7845 8230 7915 8250
rect 7630 8215 7686 8221
rect 7630 8155 7634 8215
rect 7715 8205 7915 8230
rect 7970 8221 8000 8409
rect 7944 8215 8000 8221
rect 7686 8155 7944 8175
rect 7996 8155 8000 8215
rect 7630 8145 8000 8155
rect 8030 8475 8400 8485
rect 8030 8415 8034 8475
rect 8086 8455 8344 8475
rect 8030 8409 8086 8415
rect 8030 8221 8060 8409
rect 8115 8400 8315 8425
rect 8396 8415 8400 8475
rect 8344 8409 8400 8415
rect 8115 8380 8185 8400
rect 8090 8340 8185 8380
rect 8245 8380 8315 8400
rect 8245 8340 8340 8380
rect 8090 8290 8340 8340
rect 8090 8250 8185 8290
rect 8115 8230 8185 8250
rect 8245 8250 8340 8290
rect 8245 8230 8315 8250
rect 8030 8215 8086 8221
rect 8030 8155 8034 8215
rect 8115 8205 8315 8230
rect 8370 8221 8400 8409
rect 8344 8215 8400 8221
rect 8086 8155 8344 8175
rect 8396 8155 8400 8215
rect 8030 8145 8400 8155
rect 8430 8475 8800 8485
rect 8430 8415 8434 8475
rect 8486 8455 8744 8475
rect 8430 8409 8486 8415
rect 8430 8221 8460 8409
rect 8515 8400 8715 8425
rect 8796 8415 8800 8475
rect 8744 8409 8800 8415
rect 8515 8380 8585 8400
rect 8490 8340 8585 8380
rect 8645 8380 8715 8400
rect 8645 8340 8740 8380
rect 8490 8290 8740 8340
rect 8490 8250 8585 8290
rect 8515 8230 8585 8250
rect 8645 8250 8740 8290
rect 8645 8230 8715 8250
rect 8430 8215 8486 8221
rect 8430 8155 8434 8215
rect 8515 8205 8715 8230
rect 8770 8221 8800 8409
rect 8744 8215 8800 8221
rect 8486 8155 8744 8175
rect 8796 8155 8800 8215
rect 8430 8145 8800 8155
rect 8830 8475 9200 8485
rect 8830 8415 8834 8475
rect 8886 8455 9144 8475
rect 8830 8409 8886 8415
rect 8830 8221 8860 8409
rect 8915 8400 9115 8425
rect 9196 8415 9200 8475
rect 9144 8409 9200 8415
rect 8915 8380 8985 8400
rect 8890 8340 8985 8380
rect 9045 8380 9115 8400
rect 9045 8340 9140 8380
rect 8890 8290 9140 8340
rect 8890 8250 8985 8290
rect 8915 8230 8985 8250
rect 9045 8250 9140 8290
rect 9045 8230 9115 8250
rect 8830 8215 8886 8221
rect 8830 8155 8834 8215
rect 8915 8205 9115 8230
rect 9170 8221 9200 8409
rect 9144 8215 9200 8221
rect 8886 8155 9144 8175
rect 9196 8155 9200 8215
rect 8830 8145 9200 8155
rect 9230 8475 9600 8485
rect 9230 8415 9234 8475
rect 9286 8455 9544 8475
rect 9230 8409 9286 8415
rect 9230 8221 9260 8409
rect 9315 8400 9515 8425
rect 9596 8415 9600 8475
rect 9544 8409 9600 8415
rect 9315 8380 9385 8400
rect 9290 8340 9385 8380
rect 9445 8380 9515 8400
rect 9445 8340 9540 8380
rect 9290 8290 9540 8340
rect 9290 8250 9385 8290
rect 9315 8230 9385 8250
rect 9445 8250 9540 8290
rect 9445 8230 9515 8250
rect 9230 8215 9286 8221
rect 9230 8155 9234 8215
rect 9315 8205 9515 8230
rect 9570 8221 9600 8409
rect 9544 8215 9600 8221
rect 9286 8155 9544 8175
rect 9596 8155 9600 8215
rect 9230 8145 9600 8155
rect 9630 8475 10000 8485
rect 9630 8415 9634 8475
rect 9686 8455 9944 8475
rect 9630 8409 9686 8415
rect 9630 8221 9660 8409
rect 9715 8400 9915 8425
rect 9996 8415 10000 8475
rect 9944 8409 10000 8415
rect 9715 8380 9785 8400
rect 9690 8340 9785 8380
rect 9845 8380 9915 8400
rect 9845 8340 9940 8380
rect 9690 8290 9940 8340
rect 9690 8250 9785 8290
rect 9715 8230 9785 8250
rect 9845 8250 9940 8290
rect 9845 8230 9915 8250
rect 9630 8215 9686 8221
rect 9630 8155 9634 8215
rect 9715 8205 9915 8230
rect 9970 8221 10000 8409
rect 9944 8215 10000 8221
rect 9686 8155 9944 8175
rect 9996 8155 10000 8215
rect 9630 8145 10000 8155
rect 10030 8475 10400 8485
rect 10030 8415 10034 8475
rect 10086 8455 10344 8475
rect 10030 8409 10086 8415
rect 10030 8221 10060 8409
rect 10115 8400 10315 8425
rect 10396 8415 10400 8475
rect 10344 8409 10400 8415
rect 10115 8380 10185 8400
rect 10090 8340 10185 8380
rect 10245 8380 10315 8400
rect 10245 8340 10340 8380
rect 10090 8290 10340 8340
rect 10090 8250 10185 8290
rect 10115 8230 10185 8250
rect 10245 8250 10340 8290
rect 10245 8230 10315 8250
rect 10030 8215 10086 8221
rect 10030 8155 10034 8215
rect 10115 8205 10315 8230
rect 10370 8221 10400 8409
rect 10344 8215 10400 8221
rect 10086 8155 10344 8175
rect 10396 8155 10400 8215
rect 10030 8145 10400 8155
rect 10430 8475 10800 8485
rect 10430 8415 10434 8475
rect 10486 8455 10744 8475
rect 10430 8409 10486 8415
rect 10430 8221 10460 8409
rect 10515 8400 10715 8425
rect 10796 8415 10800 8475
rect 10744 8409 10800 8415
rect 10515 8380 10585 8400
rect 10490 8340 10585 8380
rect 10645 8380 10715 8400
rect 10645 8340 10740 8380
rect 10490 8290 10740 8340
rect 10490 8250 10585 8290
rect 10515 8230 10585 8250
rect 10645 8250 10740 8290
rect 10645 8230 10715 8250
rect 10430 8215 10486 8221
rect 10430 8155 10434 8215
rect 10515 8205 10715 8230
rect 10770 8221 10800 8409
rect 10744 8215 10800 8221
rect 10486 8155 10744 8175
rect 10796 8155 10800 8215
rect 10430 8145 10800 8155
rect 10830 8475 11200 8485
rect 10830 8415 10834 8475
rect 10886 8455 11144 8475
rect 10830 8409 10886 8415
rect 10830 8221 10860 8409
rect 10915 8400 11115 8425
rect 11196 8415 11200 8475
rect 11144 8409 11200 8415
rect 10915 8380 10985 8400
rect 10890 8340 10985 8380
rect 11045 8380 11115 8400
rect 11045 8340 11140 8380
rect 10890 8290 11140 8340
rect 10890 8250 10985 8290
rect 10915 8230 10985 8250
rect 11045 8250 11140 8290
rect 11045 8230 11115 8250
rect 10830 8215 10886 8221
rect 10830 8155 10834 8215
rect 10915 8205 11115 8230
rect 11170 8221 11200 8409
rect 11144 8215 11200 8221
rect 10886 8155 11144 8175
rect 11196 8155 11200 8215
rect 10830 8145 11200 8155
rect 11230 8475 11600 8485
rect 11230 8415 11234 8475
rect 11286 8455 11544 8475
rect 11230 8409 11286 8415
rect 11230 8221 11260 8409
rect 11315 8400 11515 8425
rect 11596 8415 11600 8475
rect 11544 8409 11600 8415
rect 11315 8380 11385 8400
rect 11290 8340 11385 8380
rect 11445 8380 11515 8400
rect 11445 8340 11540 8380
rect 11290 8290 11540 8340
rect 11290 8250 11385 8290
rect 11315 8230 11385 8250
rect 11445 8250 11540 8290
rect 11445 8230 11515 8250
rect 11230 8215 11286 8221
rect 11230 8155 11234 8215
rect 11315 8205 11515 8230
rect 11570 8221 11600 8409
rect 11544 8215 11600 8221
rect 11286 8155 11544 8175
rect 11596 8155 11600 8215
rect 11230 8145 11600 8155
rect 11630 8475 12000 8485
rect 11630 8415 11634 8475
rect 11686 8455 11944 8475
rect 11630 8409 11686 8415
rect 11630 8221 11660 8409
rect 11715 8400 11915 8425
rect 11996 8415 12000 8475
rect 11944 8409 12000 8415
rect 11715 8380 11785 8400
rect 11690 8340 11785 8380
rect 11845 8380 11915 8400
rect 11845 8340 11940 8380
rect 11690 8290 11940 8340
rect 11690 8250 11785 8290
rect 11715 8230 11785 8250
rect 11845 8250 11940 8290
rect 11845 8230 11915 8250
rect 11630 8215 11686 8221
rect 11630 8155 11634 8215
rect 11715 8205 11915 8230
rect 11970 8221 12000 8409
rect 11944 8215 12000 8221
rect 11686 8155 11944 8175
rect 11996 8155 12000 8215
rect 11630 8145 12000 8155
rect 12030 8475 12400 8485
rect 12030 8415 12034 8475
rect 12086 8455 12344 8475
rect 12030 8409 12086 8415
rect 12030 8221 12060 8409
rect 12115 8400 12315 8425
rect 12396 8415 12400 8475
rect 12344 8409 12400 8415
rect 12115 8380 12185 8400
rect 12090 8340 12185 8380
rect 12245 8380 12315 8400
rect 12245 8340 12340 8380
rect 12090 8290 12340 8340
rect 12090 8250 12185 8290
rect 12115 8230 12185 8250
rect 12245 8250 12340 8290
rect 12245 8230 12315 8250
rect 12030 8215 12086 8221
rect 12030 8155 12034 8215
rect 12115 8205 12315 8230
rect 12370 8221 12400 8409
rect 12344 8215 12400 8221
rect 12086 8155 12344 8175
rect 12396 8155 12400 8215
rect 12030 8145 12400 8155
rect 12430 8475 12800 8485
rect 12430 8415 12434 8475
rect 12486 8455 12744 8475
rect 12430 8409 12486 8415
rect 12430 8221 12460 8409
rect 12515 8400 12715 8425
rect 12796 8415 12800 8475
rect 12744 8409 12800 8415
rect 12515 8380 12585 8400
rect 12490 8340 12585 8380
rect 12645 8380 12715 8400
rect 12645 8340 12740 8380
rect 12490 8290 12740 8340
rect 12490 8250 12585 8290
rect 12515 8230 12585 8250
rect 12645 8250 12740 8290
rect 12645 8230 12715 8250
rect 12430 8215 12486 8221
rect 12430 8155 12434 8215
rect 12515 8205 12715 8230
rect 12770 8221 12800 8409
rect 12744 8215 12800 8221
rect 12486 8155 12744 8175
rect 12796 8155 12800 8215
rect 12430 8145 12800 8155
rect 12830 8475 13200 8485
rect 12830 8415 12834 8475
rect 12886 8455 13144 8475
rect 12830 8409 12886 8415
rect 12830 8221 12860 8409
rect 12915 8400 13115 8425
rect 13196 8415 13200 8475
rect 13144 8409 13200 8415
rect 12915 8380 12985 8400
rect 12890 8340 12985 8380
rect 13045 8380 13115 8400
rect 13045 8340 13140 8380
rect 12890 8290 13140 8340
rect 12890 8250 12985 8290
rect 12915 8230 12985 8250
rect 13045 8250 13140 8290
rect 13045 8230 13115 8250
rect 12830 8215 12886 8221
rect 12830 8155 12834 8215
rect 12915 8205 13115 8230
rect 13170 8221 13200 8409
rect 13144 8215 13200 8221
rect 12886 8155 13144 8175
rect 13196 8155 13200 8215
rect 12830 8145 13200 8155
rect -370 8105 0 8115
rect -370 8045 -366 8105
rect -314 8085 -56 8105
rect -370 8039 -314 8045
rect -370 7851 -340 8039
rect -285 8030 -85 8055
rect -4 8045 0 8105
rect -56 8039 0 8045
rect -285 8010 -215 8030
rect -310 7970 -215 8010
rect -155 8010 -85 8030
rect -155 7970 -60 8010
rect -310 7920 -60 7970
rect -310 7880 -215 7920
rect -285 7860 -215 7880
rect -155 7880 -60 7920
rect -155 7860 -85 7880
rect -370 7845 -314 7851
rect -370 7785 -366 7845
rect -285 7835 -85 7860
rect -30 7851 0 8039
rect -56 7845 0 7851
rect -314 7785 -56 7805
rect -4 7785 0 7845
rect -370 7775 0 7785
rect 30 8105 400 8115
rect 30 8045 34 8105
rect 86 8085 344 8105
rect 30 8039 86 8045
rect 30 7851 60 8039
rect 115 8030 315 8055
rect 396 8045 400 8105
rect 344 8039 400 8045
rect 115 8010 185 8030
rect 90 7970 185 8010
rect 245 8010 315 8030
rect 245 7970 340 8010
rect 90 7920 340 7970
rect 90 7880 185 7920
rect 115 7860 185 7880
rect 245 7880 340 7920
rect 245 7860 315 7880
rect 30 7845 86 7851
rect 30 7785 34 7845
rect 115 7835 315 7860
rect 370 7851 400 8039
rect 344 7845 400 7851
rect 86 7785 344 7805
rect 396 7785 400 7845
rect 30 7775 400 7785
rect 430 8105 800 8115
rect 430 8045 434 8105
rect 486 8085 744 8105
rect 430 8039 486 8045
rect 430 7851 460 8039
rect 515 8030 715 8055
rect 796 8045 800 8105
rect 744 8039 800 8045
rect 515 8010 585 8030
rect 490 7970 585 8010
rect 645 8010 715 8030
rect 645 7970 740 8010
rect 490 7920 740 7970
rect 490 7880 585 7920
rect 515 7860 585 7880
rect 645 7880 740 7920
rect 645 7860 715 7880
rect 430 7845 486 7851
rect 430 7785 434 7845
rect 515 7835 715 7860
rect 770 7851 800 8039
rect 744 7845 800 7851
rect 486 7785 744 7805
rect 796 7785 800 7845
rect 430 7775 800 7785
rect 830 8105 1200 8115
rect 830 8045 834 8105
rect 886 8085 1144 8105
rect 830 8039 886 8045
rect 830 7851 860 8039
rect 915 8030 1115 8055
rect 1196 8045 1200 8105
rect 1144 8039 1200 8045
rect 915 8010 985 8030
rect 890 7970 985 8010
rect 1045 8010 1115 8030
rect 1045 7970 1140 8010
rect 890 7920 1140 7970
rect 890 7880 985 7920
rect 915 7860 985 7880
rect 1045 7880 1140 7920
rect 1045 7860 1115 7880
rect 830 7845 886 7851
rect 830 7785 834 7845
rect 915 7835 1115 7860
rect 1170 7851 1200 8039
rect 1144 7845 1200 7851
rect 886 7785 1144 7805
rect 1196 7785 1200 7845
rect 830 7775 1200 7785
rect 1230 8105 1600 8115
rect 1230 8045 1234 8105
rect 1286 8085 1544 8105
rect 1230 8039 1286 8045
rect 1230 7851 1260 8039
rect 1315 8030 1515 8055
rect 1596 8045 1600 8105
rect 1544 8039 1600 8045
rect 1315 8010 1385 8030
rect 1290 7970 1385 8010
rect 1445 8010 1515 8030
rect 1445 7970 1540 8010
rect 1290 7920 1540 7970
rect 1290 7880 1385 7920
rect 1315 7860 1385 7880
rect 1445 7880 1540 7920
rect 1445 7860 1515 7880
rect 1230 7845 1286 7851
rect 1230 7785 1234 7845
rect 1315 7835 1515 7860
rect 1570 7851 1600 8039
rect 1544 7845 1600 7851
rect 1286 7785 1544 7805
rect 1596 7785 1600 7845
rect 1230 7775 1600 7785
rect 1630 8105 2000 8115
rect 1630 8045 1634 8105
rect 1686 8085 1944 8105
rect 1630 8039 1686 8045
rect 1630 7851 1660 8039
rect 1715 8030 1915 8055
rect 1996 8045 2000 8105
rect 1944 8039 2000 8045
rect 1715 8010 1785 8030
rect 1690 7970 1785 8010
rect 1845 8010 1915 8030
rect 1845 7970 1940 8010
rect 1690 7920 1940 7970
rect 1690 7880 1785 7920
rect 1715 7860 1785 7880
rect 1845 7880 1940 7920
rect 1845 7860 1915 7880
rect 1630 7845 1686 7851
rect 1630 7785 1634 7845
rect 1715 7835 1915 7860
rect 1970 7851 2000 8039
rect 1944 7845 2000 7851
rect 1686 7785 1944 7805
rect 1996 7785 2000 7845
rect 1630 7775 2000 7785
rect 2030 8105 2400 8115
rect 2030 8045 2034 8105
rect 2086 8085 2344 8105
rect 2030 8039 2086 8045
rect 2030 7851 2060 8039
rect 2115 8030 2315 8055
rect 2396 8045 2400 8105
rect 2344 8039 2400 8045
rect 2115 8010 2185 8030
rect 2090 7970 2185 8010
rect 2245 8010 2315 8030
rect 2245 7970 2340 8010
rect 2090 7920 2340 7970
rect 2090 7880 2185 7920
rect 2115 7860 2185 7880
rect 2245 7880 2340 7920
rect 2245 7860 2315 7880
rect 2030 7845 2086 7851
rect 2030 7785 2034 7845
rect 2115 7835 2315 7860
rect 2370 7851 2400 8039
rect 2344 7845 2400 7851
rect 2086 7785 2344 7805
rect 2396 7785 2400 7845
rect 2030 7775 2400 7785
rect 2430 8105 2800 8115
rect 2430 8045 2434 8105
rect 2486 8085 2744 8105
rect 2430 8039 2486 8045
rect 2430 7851 2460 8039
rect 2515 8030 2715 8055
rect 2796 8045 2800 8105
rect 2744 8039 2800 8045
rect 2515 8010 2585 8030
rect 2490 7970 2585 8010
rect 2645 8010 2715 8030
rect 2645 7970 2740 8010
rect 2490 7920 2740 7970
rect 2490 7880 2585 7920
rect 2515 7860 2585 7880
rect 2645 7880 2740 7920
rect 2645 7860 2715 7880
rect 2430 7845 2486 7851
rect 2430 7785 2434 7845
rect 2515 7835 2715 7860
rect 2770 7851 2800 8039
rect 2744 7845 2800 7851
rect 2486 7785 2744 7805
rect 2796 7785 2800 7845
rect 2430 7775 2800 7785
rect 2830 8105 3200 8115
rect 2830 8045 2834 8105
rect 2886 8085 3144 8105
rect 2830 8039 2886 8045
rect 2830 7851 2860 8039
rect 2915 8030 3115 8055
rect 3196 8045 3200 8105
rect 3144 8039 3200 8045
rect 2915 8010 2985 8030
rect 2890 7970 2985 8010
rect 3045 8010 3115 8030
rect 3045 7970 3140 8010
rect 2890 7920 3140 7970
rect 2890 7880 2985 7920
rect 2915 7860 2985 7880
rect 3045 7880 3140 7920
rect 3045 7860 3115 7880
rect 2830 7845 2886 7851
rect 2830 7785 2834 7845
rect 2915 7835 3115 7860
rect 3170 7851 3200 8039
rect 3144 7845 3200 7851
rect 2886 7785 3144 7805
rect 3196 7785 3200 7845
rect 2830 7775 3200 7785
rect 3230 8105 3600 8115
rect 3230 8045 3234 8105
rect 3286 8085 3544 8105
rect 3230 8039 3286 8045
rect 3230 7851 3260 8039
rect 3315 8030 3515 8055
rect 3596 8045 3600 8105
rect 3544 8039 3600 8045
rect 3315 8010 3385 8030
rect 3290 7970 3385 8010
rect 3445 8010 3515 8030
rect 3445 7970 3540 8010
rect 3290 7920 3540 7970
rect 3290 7880 3385 7920
rect 3315 7860 3385 7880
rect 3445 7880 3540 7920
rect 3445 7860 3515 7880
rect 3230 7845 3286 7851
rect 3230 7785 3234 7845
rect 3315 7835 3515 7860
rect 3570 7851 3600 8039
rect 3544 7845 3600 7851
rect 3286 7785 3544 7805
rect 3596 7785 3600 7845
rect 3230 7775 3600 7785
rect 3630 8105 4000 8115
rect 3630 8045 3634 8105
rect 3686 8085 3944 8105
rect 3630 8039 3686 8045
rect 3630 7851 3660 8039
rect 3715 8030 3915 8055
rect 3996 8045 4000 8105
rect 3944 8039 4000 8045
rect 3715 8010 3785 8030
rect 3690 7970 3785 8010
rect 3845 8010 3915 8030
rect 3845 7970 3940 8010
rect 3690 7920 3940 7970
rect 3690 7880 3785 7920
rect 3715 7860 3785 7880
rect 3845 7880 3940 7920
rect 3845 7860 3915 7880
rect 3630 7845 3686 7851
rect 3630 7785 3634 7845
rect 3715 7835 3915 7860
rect 3970 7851 4000 8039
rect 3944 7845 4000 7851
rect 3686 7785 3944 7805
rect 3996 7785 4000 7845
rect 3630 7775 4000 7785
rect 4030 8105 4400 8115
rect 4030 8045 4034 8105
rect 4086 8085 4344 8105
rect 4030 8039 4086 8045
rect 4030 7851 4060 8039
rect 4115 8030 4315 8055
rect 4396 8045 4400 8105
rect 4344 8039 4400 8045
rect 4115 8010 4185 8030
rect 4090 7970 4185 8010
rect 4245 8010 4315 8030
rect 4245 7970 4340 8010
rect 4090 7920 4340 7970
rect 4090 7880 4185 7920
rect 4115 7860 4185 7880
rect 4245 7880 4340 7920
rect 4245 7860 4315 7880
rect 4030 7845 4086 7851
rect 4030 7785 4034 7845
rect 4115 7835 4315 7860
rect 4370 7851 4400 8039
rect 4344 7845 4400 7851
rect 4086 7785 4344 7805
rect 4396 7785 4400 7845
rect 4030 7775 4400 7785
rect 4430 8105 4800 8115
rect 4430 8045 4434 8105
rect 4486 8085 4744 8105
rect 4430 8039 4486 8045
rect 4430 7851 4460 8039
rect 4515 8030 4715 8055
rect 4796 8045 4800 8105
rect 4744 8039 4800 8045
rect 4515 8010 4585 8030
rect 4490 7970 4585 8010
rect 4645 8010 4715 8030
rect 4645 7970 4740 8010
rect 4490 7920 4740 7970
rect 4490 7880 4585 7920
rect 4515 7860 4585 7880
rect 4645 7880 4740 7920
rect 4645 7860 4715 7880
rect 4430 7845 4486 7851
rect 4430 7785 4434 7845
rect 4515 7835 4715 7860
rect 4770 7851 4800 8039
rect 4744 7845 4800 7851
rect 4486 7785 4744 7805
rect 4796 7785 4800 7845
rect 4430 7775 4800 7785
rect 4830 8105 5200 8115
rect 4830 8045 4834 8105
rect 4886 8085 5144 8105
rect 4830 8039 4886 8045
rect 4830 7851 4860 8039
rect 4915 8030 5115 8055
rect 5196 8045 5200 8105
rect 5144 8039 5200 8045
rect 4915 8010 4985 8030
rect 4890 7970 4985 8010
rect 5045 8010 5115 8030
rect 5045 7970 5140 8010
rect 4890 7920 5140 7970
rect 4890 7880 4985 7920
rect 4915 7860 4985 7880
rect 5045 7880 5140 7920
rect 5045 7860 5115 7880
rect 4830 7845 4886 7851
rect 4830 7785 4834 7845
rect 4915 7835 5115 7860
rect 5170 7851 5200 8039
rect 5144 7845 5200 7851
rect 4886 7785 5144 7805
rect 5196 7785 5200 7845
rect 4830 7775 5200 7785
rect 5230 8105 5600 8115
rect 5230 8045 5234 8105
rect 5286 8085 5544 8105
rect 5230 8039 5286 8045
rect 5230 7851 5260 8039
rect 5315 8030 5515 8055
rect 5596 8045 5600 8105
rect 5544 8039 5600 8045
rect 5315 8010 5385 8030
rect 5290 7970 5385 8010
rect 5445 8010 5515 8030
rect 5445 7970 5540 8010
rect 5290 7920 5540 7970
rect 5290 7880 5385 7920
rect 5315 7860 5385 7880
rect 5445 7880 5540 7920
rect 5445 7860 5515 7880
rect 5230 7845 5286 7851
rect 5230 7785 5234 7845
rect 5315 7835 5515 7860
rect 5570 7851 5600 8039
rect 5544 7845 5600 7851
rect 5286 7785 5544 7805
rect 5596 7785 5600 7845
rect 5230 7775 5600 7785
rect 5630 8105 6000 8115
rect 5630 8045 5634 8105
rect 5686 8085 5944 8105
rect 5630 8039 5686 8045
rect 5630 7851 5660 8039
rect 5715 8030 5915 8055
rect 5996 8045 6000 8105
rect 5944 8039 6000 8045
rect 5715 8010 5785 8030
rect 5690 7970 5785 8010
rect 5845 8010 5915 8030
rect 5845 7970 5940 8010
rect 5690 7920 5940 7970
rect 5690 7880 5785 7920
rect 5715 7860 5785 7880
rect 5845 7880 5940 7920
rect 5845 7860 5915 7880
rect 5630 7845 5686 7851
rect 5630 7785 5634 7845
rect 5715 7835 5915 7860
rect 5970 7851 6000 8039
rect 5944 7845 6000 7851
rect 5686 7785 5944 7805
rect 5996 7785 6000 7845
rect 5630 7775 6000 7785
rect 6030 8105 6400 8115
rect 6030 8045 6034 8105
rect 6086 8085 6344 8105
rect 6030 8039 6086 8045
rect 6030 7851 6060 8039
rect 6115 8030 6315 8055
rect 6396 8045 6400 8105
rect 6344 8039 6400 8045
rect 6115 8010 6185 8030
rect 6090 7970 6185 8010
rect 6245 8010 6315 8030
rect 6245 7970 6340 8010
rect 6090 7920 6340 7970
rect 6090 7880 6185 7920
rect 6115 7860 6185 7880
rect 6245 7880 6340 7920
rect 6245 7860 6315 7880
rect 6030 7845 6086 7851
rect 6030 7785 6034 7845
rect 6115 7835 6315 7860
rect 6370 7851 6400 8039
rect 6344 7845 6400 7851
rect 6086 7785 6344 7805
rect 6396 7785 6400 7845
rect 6030 7775 6400 7785
rect 6430 8105 6800 8115
rect 6430 8045 6434 8105
rect 6486 8085 6744 8105
rect 6430 8039 6486 8045
rect 6430 7851 6460 8039
rect 6515 8030 6715 8055
rect 6796 8045 6800 8105
rect 6744 8039 6800 8045
rect 6515 8010 6585 8030
rect 6490 7970 6585 8010
rect 6645 8010 6715 8030
rect 6645 7970 6740 8010
rect 6490 7920 6740 7970
rect 6490 7880 6585 7920
rect 6515 7860 6585 7880
rect 6645 7880 6740 7920
rect 6645 7860 6715 7880
rect 6430 7845 6486 7851
rect 6430 7785 6434 7845
rect 6515 7835 6715 7860
rect 6770 7851 6800 8039
rect 6744 7845 6800 7851
rect 6486 7785 6744 7805
rect 6796 7785 6800 7845
rect 6430 7775 6800 7785
rect 6830 8105 7200 8115
rect 6830 8045 6834 8105
rect 6886 8085 7144 8105
rect 6830 8039 6886 8045
rect 6830 7851 6860 8039
rect 6915 8030 7115 8055
rect 7196 8045 7200 8105
rect 7144 8039 7200 8045
rect 6915 8010 6985 8030
rect 6890 7970 6985 8010
rect 7045 8010 7115 8030
rect 7045 7970 7140 8010
rect 6890 7920 7140 7970
rect 6890 7880 6985 7920
rect 6915 7860 6985 7880
rect 7045 7880 7140 7920
rect 7045 7860 7115 7880
rect 6830 7845 6886 7851
rect 6830 7785 6834 7845
rect 6915 7835 7115 7860
rect 7170 7851 7200 8039
rect 7144 7845 7200 7851
rect 6886 7785 7144 7805
rect 7196 7785 7200 7845
rect 6830 7775 7200 7785
rect 7230 8105 7600 8115
rect 7230 8045 7234 8105
rect 7286 8085 7544 8105
rect 7230 8039 7286 8045
rect 7230 7851 7260 8039
rect 7315 8030 7515 8055
rect 7596 8045 7600 8105
rect 7544 8039 7600 8045
rect 7315 8010 7385 8030
rect 7290 7970 7385 8010
rect 7445 8010 7515 8030
rect 7445 7970 7540 8010
rect 7290 7920 7540 7970
rect 7290 7880 7385 7920
rect 7315 7860 7385 7880
rect 7445 7880 7540 7920
rect 7445 7860 7515 7880
rect 7230 7845 7286 7851
rect 7230 7785 7234 7845
rect 7315 7835 7515 7860
rect 7570 7851 7600 8039
rect 7544 7845 7600 7851
rect 7286 7785 7544 7805
rect 7596 7785 7600 7845
rect 7230 7775 7600 7785
rect 7630 8105 8000 8115
rect 7630 8045 7634 8105
rect 7686 8085 7944 8105
rect 7630 8039 7686 8045
rect 7630 7851 7660 8039
rect 7715 8030 7915 8055
rect 7996 8045 8000 8105
rect 7944 8039 8000 8045
rect 7715 8010 7785 8030
rect 7690 7970 7785 8010
rect 7845 8010 7915 8030
rect 7845 7970 7940 8010
rect 7690 7920 7940 7970
rect 7690 7880 7785 7920
rect 7715 7860 7785 7880
rect 7845 7880 7940 7920
rect 7845 7860 7915 7880
rect 7630 7845 7686 7851
rect 7630 7785 7634 7845
rect 7715 7835 7915 7860
rect 7970 7851 8000 8039
rect 7944 7845 8000 7851
rect 7686 7785 7944 7805
rect 7996 7785 8000 7845
rect 7630 7775 8000 7785
rect 8030 8105 8400 8115
rect 8030 8045 8034 8105
rect 8086 8085 8344 8105
rect 8030 8039 8086 8045
rect 8030 7851 8060 8039
rect 8115 8030 8315 8055
rect 8396 8045 8400 8105
rect 8344 8039 8400 8045
rect 8115 8010 8185 8030
rect 8090 7970 8185 8010
rect 8245 8010 8315 8030
rect 8245 7970 8340 8010
rect 8090 7920 8340 7970
rect 8090 7880 8185 7920
rect 8115 7860 8185 7880
rect 8245 7880 8340 7920
rect 8245 7860 8315 7880
rect 8030 7845 8086 7851
rect 8030 7785 8034 7845
rect 8115 7835 8315 7860
rect 8370 7851 8400 8039
rect 8344 7845 8400 7851
rect 8086 7785 8344 7805
rect 8396 7785 8400 7845
rect 8030 7775 8400 7785
rect 8430 8105 8800 8115
rect 8430 8045 8434 8105
rect 8486 8085 8744 8105
rect 8430 8039 8486 8045
rect 8430 7851 8460 8039
rect 8515 8030 8715 8055
rect 8796 8045 8800 8105
rect 8744 8039 8800 8045
rect 8515 8010 8585 8030
rect 8490 7970 8585 8010
rect 8645 8010 8715 8030
rect 8645 7970 8740 8010
rect 8490 7920 8740 7970
rect 8490 7880 8585 7920
rect 8515 7860 8585 7880
rect 8645 7880 8740 7920
rect 8645 7860 8715 7880
rect 8430 7845 8486 7851
rect 8430 7785 8434 7845
rect 8515 7835 8715 7860
rect 8770 7851 8800 8039
rect 8744 7845 8800 7851
rect 8486 7785 8744 7805
rect 8796 7785 8800 7845
rect 8430 7775 8800 7785
rect 8830 8105 9200 8115
rect 8830 8045 8834 8105
rect 8886 8085 9144 8105
rect 8830 8039 8886 8045
rect 8830 7851 8860 8039
rect 8915 8030 9115 8055
rect 9196 8045 9200 8105
rect 9144 8039 9200 8045
rect 8915 8010 8985 8030
rect 8890 7970 8985 8010
rect 9045 8010 9115 8030
rect 9045 7970 9140 8010
rect 8890 7920 9140 7970
rect 8890 7880 8985 7920
rect 8915 7860 8985 7880
rect 9045 7880 9140 7920
rect 9045 7860 9115 7880
rect 8830 7845 8886 7851
rect 8830 7785 8834 7845
rect 8915 7835 9115 7860
rect 9170 7851 9200 8039
rect 9144 7845 9200 7851
rect 8886 7785 9144 7805
rect 9196 7785 9200 7845
rect 8830 7775 9200 7785
rect 9230 8105 9600 8115
rect 9230 8045 9234 8105
rect 9286 8085 9544 8105
rect 9230 8039 9286 8045
rect 9230 7851 9260 8039
rect 9315 8030 9515 8055
rect 9596 8045 9600 8105
rect 9544 8039 9600 8045
rect 9315 8010 9385 8030
rect 9290 7970 9385 8010
rect 9445 8010 9515 8030
rect 9445 7970 9540 8010
rect 9290 7920 9540 7970
rect 9290 7880 9385 7920
rect 9315 7860 9385 7880
rect 9445 7880 9540 7920
rect 9445 7860 9515 7880
rect 9230 7845 9286 7851
rect 9230 7785 9234 7845
rect 9315 7835 9515 7860
rect 9570 7851 9600 8039
rect 9544 7845 9600 7851
rect 9286 7785 9544 7805
rect 9596 7785 9600 7845
rect 9230 7775 9600 7785
rect 9630 8105 10000 8115
rect 9630 8045 9634 8105
rect 9686 8085 9944 8105
rect 9630 8039 9686 8045
rect 9630 7851 9660 8039
rect 9715 8030 9915 8055
rect 9996 8045 10000 8105
rect 9944 8039 10000 8045
rect 9715 8010 9785 8030
rect 9690 7970 9785 8010
rect 9845 8010 9915 8030
rect 9845 7970 9940 8010
rect 9690 7920 9940 7970
rect 9690 7880 9785 7920
rect 9715 7860 9785 7880
rect 9845 7880 9940 7920
rect 9845 7860 9915 7880
rect 9630 7845 9686 7851
rect 9630 7785 9634 7845
rect 9715 7835 9915 7860
rect 9970 7851 10000 8039
rect 9944 7845 10000 7851
rect 9686 7785 9944 7805
rect 9996 7785 10000 7845
rect 9630 7775 10000 7785
rect 10030 8105 10400 8115
rect 10030 8045 10034 8105
rect 10086 8085 10344 8105
rect 10030 8039 10086 8045
rect 10030 7851 10060 8039
rect 10115 8030 10315 8055
rect 10396 8045 10400 8105
rect 10344 8039 10400 8045
rect 10115 8010 10185 8030
rect 10090 7970 10185 8010
rect 10245 8010 10315 8030
rect 10245 7970 10340 8010
rect 10090 7920 10340 7970
rect 10090 7880 10185 7920
rect 10115 7860 10185 7880
rect 10245 7880 10340 7920
rect 10245 7860 10315 7880
rect 10030 7845 10086 7851
rect 10030 7785 10034 7845
rect 10115 7835 10315 7860
rect 10370 7851 10400 8039
rect 10344 7845 10400 7851
rect 10086 7785 10344 7805
rect 10396 7785 10400 7845
rect 10030 7775 10400 7785
rect 10430 8105 10800 8115
rect 10430 8045 10434 8105
rect 10486 8085 10744 8105
rect 10430 8039 10486 8045
rect 10430 7851 10460 8039
rect 10515 8030 10715 8055
rect 10796 8045 10800 8105
rect 10744 8039 10800 8045
rect 10515 8010 10585 8030
rect 10490 7970 10585 8010
rect 10645 8010 10715 8030
rect 10645 7970 10740 8010
rect 10490 7920 10740 7970
rect 10490 7880 10585 7920
rect 10515 7860 10585 7880
rect 10645 7880 10740 7920
rect 10645 7860 10715 7880
rect 10430 7845 10486 7851
rect 10430 7785 10434 7845
rect 10515 7835 10715 7860
rect 10770 7851 10800 8039
rect 10744 7845 10800 7851
rect 10486 7785 10744 7805
rect 10796 7785 10800 7845
rect 10430 7775 10800 7785
rect 10830 8105 11200 8115
rect 10830 8045 10834 8105
rect 10886 8085 11144 8105
rect 10830 8039 10886 8045
rect 10830 7851 10860 8039
rect 10915 8030 11115 8055
rect 11196 8045 11200 8105
rect 11144 8039 11200 8045
rect 10915 8010 10985 8030
rect 10890 7970 10985 8010
rect 11045 8010 11115 8030
rect 11045 7970 11140 8010
rect 10890 7920 11140 7970
rect 10890 7880 10985 7920
rect 10915 7860 10985 7880
rect 11045 7880 11140 7920
rect 11045 7860 11115 7880
rect 10830 7845 10886 7851
rect 10830 7785 10834 7845
rect 10915 7835 11115 7860
rect 11170 7851 11200 8039
rect 11144 7845 11200 7851
rect 10886 7785 11144 7805
rect 11196 7785 11200 7845
rect 10830 7775 11200 7785
rect 11230 8105 11600 8115
rect 11230 8045 11234 8105
rect 11286 8085 11544 8105
rect 11230 8039 11286 8045
rect 11230 7851 11260 8039
rect 11315 8030 11515 8055
rect 11596 8045 11600 8105
rect 11544 8039 11600 8045
rect 11315 8010 11385 8030
rect 11290 7970 11385 8010
rect 11445 8010 11515 8030
rect 11445 7970 11540 8010
rect 11290 7920 11540 7970
rect 11290 7880 11385 7920
rect 11315 7860 11385 7880
rect 11445 7880 11540 7920
rect 11445 7860 11515 7880
rect 11230 7845 11286 7851
rect 11230 7785 11234 7845
rect 11315 7835 11515 7860
rect 11570 7851 11600 8039
rect 11544 7845 11600 7851
rect 11286 7785 11544 7805
rect 11596 7785 11600 7845
rect 11230 7775 11600 7785
rect 11630 8105 12000 8115
rect 11630 8045 11634 8105
rect 11686 8085 11944 8105
rect 11630 8039 11686 8045
rect 11630 7851 11660 8039
rect 11715 8030 11915 8055
rect 11996 8045 12000 8105
rect 11944 8039 12000 8045
rect 11715 8010 11785 8030
rect 11690 7970 11785 8010
rect 11845 8010 11915 8030
rect 11845 7970 11940 8010
rect 11690 7920 11940 7970
rect 11690 7880 11785 7920
rect 11715 7860 11785 7880
rect 11845 7880 11940 7920
rect 11845 7860 11915 7880
rect 11630 7845 11686 7851
rect 11630 7785 11634 7845
rect 11715 7835 11915 7860
rect 11970 7851 12000 8039
rect 11944 7845 12000 7851
rect 11686 7785 11944 7805
rect 11996 7785 12000 7845
rect 11630 7775 12000 7785
rect 12030 8105 12400 8115
rect 12030 8045 12034 8105
rect 12086 8085 12344 8105
rect 12030 8039 12086 8045
rect 12030 7851 12060 8039
rect 12115 8030 12315 8055
rect 12396 8045 12400 8105
rect 12344 8039 12400 8045
rect 12115 8010 12185 8030
rect 12090 7970 12185 8010
rect 12245 8010 12315 8030
rect 12245 7970 12340 8010
rect 12090 7920 12340 7970
rect 12090 7880 12185 7920
rect 12115 7860 12185 7880
rect 12245 7880 12340 7920
rect 12245 7860 12315 7880
rect 12030 7845 12086 7851
rect 12030 7785 12034 7845
rect 12115 7835 12315 7860
rect 12370 7851 12400 8039
rect 12344 7845 12400 7851
rect 12086 7785 12344 7805
rect 12396 7785 12400 7845
rect 12030 7775 12400 7785
rect 12430 8105 12800 8115
rect 12430 8045 12434 8105
rect 12486 8085 12744 8105
rect 12430 8039 12486 8045
rect 12430 7851 12460 8039
rect 12515 8030 12715 8055
rect 12796 8045 12800 8105
rect 12744 8039 12800 8045
rect 12515 8010 12585 8030
rect 12490 7970 12585 8010
rect 12645 8010 12715 8030
rect 12645 7970 12740 8010
rect 12490 7920 12740 7970
rect 12490 7880 12585 7920
rect 12515 7860 12585 7880
rect 12645 7880 12740 7920
rect 12645 7860 12715 7880
rect 12430 7845 12486 7851
rect 12430 7785 12434 7845
rect 12515 7835 12715 7860
rect 12770 7851 12800 8039
rect 12744 7845 12800 7851
rect 12486 7785 12744 7805
rect 12796 7785 12800 7845
rect 12430 7775 12800 7785
rect 12830 8105 13200 8115
rect 12830 8045 12834 8105
rect 12886 8085 13144 8105
rect 12830 8039 12886 8045
rect 12830 7851 12860 8039
rect 12915 8030 13115 8055
rect 13196 8045 13200 8105
rect 13144 8039 13200 8045
rect 12915 8010 12985 8030
rect 12890 7970 12985 8010
rect 13045 8010 13115 8030
rect 13045 7970 13140 8010
rect 12890 7920 13140 7970
rect 12890 7880 12985 7920
rect 12915 7860 12985 7880
rect 13045 7880 13140 7920
rect 13045 7860 13115 7880
rect 12830 7845 12886 7851
rect 12830 7785 12834 7845
rect 12915 7835 13115 7860
rect 13170 7851 13200 8039
rect 13144 7845 13200 7851
rect 12886 7785 13144 7805
rect 13196 7785 13200 7845
rect 12830 7775 13200 7785
rect -370 7735 0 7745
rect -370 7675 -366 7735
rect -314 7715 -56 7735
rect -370 7669 -314 7675
rect -370 7481 -340 7669
rect -285 7660 -85 7685
rect -4 7675 0 7735
rect -56 7669 0 7675
rect -285 7640 -215 7660
rect -310 7600 -215 7640
rect -155 7640 -85 7660
rect -155 7600 -60 7640
rect -310 7550 -60 7600
rect -310 7510 -215 7550
rect -285 7490 -215 7510
rect -155 7510 -60 7550
rect -155 7490 -85 7510
rect -370 7475 -314 7481
rect -370 7415 -366 7475
rect -285 7465 -85 7490
rect -30 7481 0 7669
rect -56 7475 0 7481
rect -314 7415 -56 7435
rect -4 7415 0 7475
rect -370 7405 0 7415
rect 30 7735 400 7745
rect 30 7675 34 7735
rect 86 7715 344 7735
rect 30 7669 86 7675
rect 30 7481 60 7669
rect 115 7660 315 7685
rect 396 7675 400 7735
rect 344 7669 400 7675
rect 115 7640 185 7660
rect 90 7600 185 7640
rect 245 7640 315 7660
rect 245 7600 340 7640
rect 90 7550 340 7600
rect 90 7510 185 7550
rect 115 7490 185 7510
rect 245 7510 340 7550
rect 245 7490 315 7510
rect 30 7475 86 7481
rect 30 7415 34 7475
rect 115 7465 315 7490
rect 370 7481 400 7669
rect 344 7475 400 7481
rect 86 7415 344 7435
rect 396 7415 400 7475
rect 30 7405 400 7415
rect 430 7735 800 7745
rect 430 7675 434 7735
rect 486 7715 744 7735
rect 430 7669 486 7675
rect 430 7481 460 7669
rect 515 7660 715 7685
rect 796 7675 800 7735
rect 744 7669 800 7675
rect 515 7640 585 7660
rect 490 7600 585 7640
rect 645 7640 715 7660
rect 645 7600 740 7640
rect 490 7550 740 7600
rect 490 7510 585 7550
rect 515 7490 585 7510
rect 645 7510 740 7550
rect 645 7490 715 7510
rect 430 7475 486 7481
rect 430 7415 434 7475
rect 515 7465 715 7490
rect 770 7481 800 7669
rect 744 7475 800 7481
rect 486 7415 744 7435
rect 796 7415 800 7475
rect 430 7405 800 7415
rect 830 7735 1200 7745
rect 830 7675 834 7735
rect 886 7715 1144 7735
rect 830 7669 886 7675
rect 830 7481 860 7669
rect 915 7660 1115 7685
rect 1196 7675 1200 7735
rect 1144 7669 1200 7675
rect 915 7640 985 7660
rect 890 7600 985 7640
rect 1045 7640 1115 7660
rect 1045 7600 1140 7640
rect 890 7550 1140 7600
rect 890 7510 985 7550
rect 915 7490 985 7510
rect 1045 7510 1140 7550
rect 1045 7490 1115 7510
rect 830 7475 886 7481
rect 830 7415 834 7475
rect 915 7465 1115 7490
rect 1170 7481 1200 7669
rect 1144 7475 1200 7481
rect 886 7415 1144 7435
rect 1196 7415 1200 7475
rect 830 7405 1200 7415
rect 1230 7735 1600 7745
rect 1230 7675 1234 7735
rect 1286 7715 1544 7735
rect 1230 7669 1286 7675
rect 1230 7481 1260 7669
rect 1315 7660 1515 7685
rect 1596 7675 1600 7735
rect 1544 7669 1600 7675
rect 1315 7640 1385 7660
rect 1290 7600 1385 7640
rect 1445 7640 1515 7660
rect 1445 7600 1540 7640
rect 1290 7550 1540 7600
rect 1290 7510 1385 7550
rect 1315 7490 1385 7510
rect 1445 7510 1540 7550
rect 1445 7490 1515 7510
rect 1230 7475 1286 7481
rect 1230 7415 1234 7475
rect 1315 7465 1515 7490
rect 1570 7481 1600 7669
rect 1544 7475 1600 7481
rect 1286 7415 1544 7435
rect 1596 7415 1600 7475
rect 1230 7405 1600 7415
rect 1630 7735 2000 7745
rect 1630 7675 1634 7735
rect 1686 7715 1944 7735
rect 1630 7669 1686 7675
rect 1630 7481 1660 7669
rect 1715 7660 1915 7685
rect 1996 7675 2000 7735
rect 1944 7669 2000 7675
rect 1715 7640 1785 7660
rect 1690 7600 1785 7640
rect 1845 7640 1915 7660
rect 1845 7600 1940 7640
rect 1690 7550 1940 7600
rect 1690 7510 1785 7550
rect 1715 7490 1785 7510
rect 1845 7510 1940 7550
rect 1845 7490 1915 7510
rect 1630 7475 1686 7481
rect 1630 7415 1634 7475
rect 1715 7465 1915 7490
rect 1970 7481 2000 7669
rect 1944 7475 2000 7481
rect 1686 7415 1944 7435
rect 1996 7415 2000 7475
rect 1630 7405 2000 7415
rect 2030 7735 2400 7745
rect 2030 7675 2034 7735
rect 2086 7715 2344 7735
rect 2030 7669 2086 7675
rect 2030 7481 2060 7669
rect 2115 7660 2315 7685
rect 2396 7675 2400 7735
rect 2344 7669 2400 7675
rect 2115 7640 2185 7660
rect 2090 7600 2185 7640
rect 2245 7640 2315 7660
rect 2245 7600 2340 7640
rect 2090 7550 2340 7600
rect 2090 7510 2185 7550
rect 2115 7490 2185 7510
rect 2245 7510 2340 7550
rect 2245 7490 2315 7510
rect 2030 7475 2086 7481
rect 2030 7415 2034 7475
rect 2115 7465 2315 7490
rect 2370 7481 2400 7669
rect 2344 7475 2400 7481
rect 2086 7415 2344 7435
rect 2396 7415 2400 7475
rect 2030 7405 2400 7415
rect 2430 7735 2800 7745
rect 2430 7675 2434 7735
rect 2486 7715 2744 7735
rect 2430 7669 2486 7675
rect 2430 7481 2460 7669
rect 2515 7660 2715 7685
rect 2796 7675 2800 7735
rect 2744 7669 2800 7675
rect 2515 7640 2585 7660
rect 2490 7600 2585 7640
rect 2645 7640 2715 7660
rect 2645 7600 2740 7640
rect 2490 7550 2740 7600
rect 2490 7510 2585 7550
rect 2515 7490 2585 7510
rect 2645 7510 2740 7550
rect 2645 7490 2715 7510
rect 2430 7475 2486 7481
rect 2430 7415 2434 7475
rect 2515 7465 2715 7490
rect 2770 7481 2800 7669
rect 2744 7475 2800 7481
rect 2486 7415 2744 7435
rect 2796 7415 2800 7475
rect 2430 7405 2800 7415
rect 2830 7735 3200 7745
rect 2830 7675 2834 7735
rect 2886 7715 3144 7735
rect 2830 7669 2886 7675
rect 2830 7481 2860 7669
rect 2915 7660 3115 7685
rect 3196 7675 3200 7735
rect 3144 7669 3200 7675
rect 2915 7640 2985 7660
rect 2890 7600 2985 7640
rect 3045 7640 3115 7660
rect 3045 7600 3140 7640
rect 2890 7550 3140 7600
rect 2890 7510 2985 7550
rect 2915 7490 2985 7510
rect 3045 7510 3140 7550
rect 3045 7490 3115 7510
rect 2830 7475 2886 7481
rect 2830 7415 2834 7475
rect 2915 7465 3115 7490
rect 3170 7481 3200 7669
rect 3144 7475 3200 7481
rect 2886 7415 3144 7435
rect 3196 7415 3200 7475
rect 2830 7405 3200 7415
rect 3230 7735 3600 7745
rect 3230 7675 3234 7735
rect 3286 7715 3544 7735
rect 3230 7669 3286 7675
rect 3230 7481 3260 7669
rect 3315 7660 3515 7685
rect 3596 7675 3600 7735
rect 3544 7669 3600 7675
rect 3315 7640 3385 7660
rect 3290 7600 3385 7640
rect 3445 7640 3515 7660
rect 3445 7600 3540 7640
rect 3290 7550 3540 7600
rect 3290 7510 3385 7550
rect 3315 7490 3385 7510
rect 3445 7510 3540 7550
rect 3445 7490 3515 7510
rect 3230 7475 3286 7481
rect 3230 7415 3234 7475
rect 3315 7465 3515 7490
rect 3570 7481 3600 7669
rect 3544 7475 3600 7481
rect 3286 7415 3544 7435
rect 3596 7415 3600 7475
rect 3230 7405 3600 7415
rect 3630 7735 4000 7745
rect 3630 7675 3634 7735
rect 3686 7715 3944 7735
rect 3630 7669 3686 7675
rect 3630 7481 3660 7669
rect 3715 7660 3915 7685
rect 3996 7675 4000 7735
rect 3944 7669 4000 7675
rect 3715 7640 3785 7660
rect 3690 7600 3785 7640
rect 3845 7640 3915 7660
rect 3845 7600 3940 7640
rect 3690 7550 3940 7600
rect 3690 7510 3785 7550
rect 3715 7490 3785 7510
rect 3845 7510 3940 7550
rect 3845 7490 3915 7510
rect 3630 7475 3686 7481
rect 3630 7415 3634 7475
rect 3715 7465 3915 7490
rect 3970 7481 4000 7669
rect 3944 7475 4000 7481
rect 3686 7415 3944 7435
rect 3996 7415 4000 7475
rect 3630 7405 4000 7415
rect 4030 7735 4400 7745
rect 4030 7675 4034 7735
rect 4086 7715 4344 7735
rect 4030 7669 4086 7675
rect 4030 7481 4060 7669
rect 4115 7660 4315 7685
rect 4396 7675 4400 7735
rect 4344 7669 4400 7675
rect 4115 7640 4185 7660
rect 4090 7600 4185 7640
rect 4245 7640 4315 7660
rect 4245 7600 4340 7640
rect 4090 7550 4340 7600
rect 4090 7510 4185 7550
rect 4115 7490 4185 7510
rect 4245 7510 4340 7550
rect 4245 7490 4315 7510
rect 4030 7475 4086 7481
rect 4030 7415 4034 7475
rect 4115 7465 4315 7490
rect 4370 7481 4400 7669
rect 4344 7475 4400 7481
rect 4086 7415 4344 7435
rect 4396 7415 4400 7475
rect 4030 7405 4400 7415
rect 4430 7735 4800 7745
rect 4430 7675 4434 7735
rect 4486 7715 4744 7735
rect 4430 7669 4486 7675
rect 4430 7481 4460 7669
rect 4515 7660 4715 7685
rect 4796 7675 4800 7735
rect 4744 7669 4800 7675
rect 4515 7640 4585 7660
rect 4490 7600 4585 7640
rect 4645 7640 4715 7660
rect 4645 7600 4740 7640
rect 4490 7550 4740 7600
rect 4490 7510 4585 7550
rect 4515 7490 4585 7510
rect 4645 7510 4740 7550
rect 4645 7490 4715 7510
rect 4430 7475 4486 7481
rect 4430 7415 4434 7475
rect 4515 7465 4715 7490
rect 4770 7481 4800 7669
rect 4744 7475 4800 7481
rect 4486 7415 4744 7435
rect 4796 7415 4800 7475
rect 4430 7405 4800 7415
rect 4830 7735 5200 7745
rect 4830 7675 4834 7735
rect 4886 7715 5144 7735
rect 4830 7669 4886 7675
rect 4830 7481 4860 7669
rect 4915 7660 5115 7685
rect 5196 7675 5200 7735
rect 5144 7669 5200 7675
rect 4915 7640 4985 7660
rect 4890 7600 4985 7640
rect 5045 7640 5115 7660
rect 5045 7600 5140 7640
rect 4890 7550 5140 7600
rect 4890 7510 4985 7550
rect 4915 7490 4985 7510
rect 5045 7510 5140 7550
rect 5045 7490 5115 7510
rect 4830 7475 4886 7481
rect 4830 7415 4834 7475
rect 4915 7465 5115 7490
rect 5170 7481 5200 7669
rect 5144 7475 5200 7481
rect 4886 7415 5144 7435
rect 5196 7415 5200 7475
rect 4830 7405 5200 7415
rect 5230 7735 5600 7745
rect 5230 7675 5234 7735
rect 5286 7715 5544 7735
rect 5230 7669 5286 7675
rect 5230 7481 5260 7669
rect 5315 7660 5515 7685
rect 5596 7675 5600 7735
rect 5544 7669 5600 7675
rect 5315 7640 5385 7660
rect 5290 7600 5385 7640
rect 5445 7640 5515 7660
rect 5445 7600 5540 7640
rect 5290 7550 5540 7600
rect 5290 7510 5385 7550
rect 5315 7490 5385 7510
rect 5445 7510 5540 7550
rect 5445 7490 5515 7510
rect 5230 7475 5286 7481
rect 5230 7415 5234 7475
rect 5315 7465 5515 7490
rect 5570 7481 5600 7669
rect 5544 7475 5600 7481
rect 5286 7415 5544 7435
rect 5596 7415 5600 7475
rect 5230 7405 5600 7415
rect 5630 7735 6000 7745
rect 5630 7675 5634 7735
rect 5686 7715 5944 7735
rect 5630 7669 5686 7675
rect 5630 7481 5660 7669
rect 5715 7660 5915 7685
rect 5996 7675 6000 7735
rect 5944 7669 6000 7675
rect 5715 7640 5785 7660
rect 5690 7600 5785 7640
rect 5845 7640 5915 7660
rect 5845 7600 5940 7640
rect 5690 7550 5940 7600
rect 5690 7510 5785 7550
rect 5715 7490 5785 7510
rect 5845 7510 5940 7550
rect 5845 7490 5915 7510
rect 5630 7475 5686 7481
rect 5630 7415 5634 7475
rect 5715 7465 5915 7490
rect 5970 7481 6000 7669
rect 5944 7475 6000 7481
rect 5686 7415 5944 7435
rect 5996 7415 6000 7475
rect 5630 7405 6000 7415
rect 6030 7735 6400 7745
rect 6030 7675 6034 7735
rect 6086 7715 6344 7735
rect 6030 7669 6086 7675
rect 6030 7481 6060 7669
rect 6115 7660 6315 7685
rect 6396 7675 6400 7735
rect 6344 7669 6400 7675
rect 6115 7640 6185 7660
rect 6090 7600 6185 7640
rect 6245 7640 6315 7660
rect 6245 7600 6340 7640
rect 6090 7550 6340 7600
rect 6090 7510 6185 7550
rect 6115 7490 6185 7510
rect 6245 7510 6340 7550
rect 6245 7490 6315 7510
rect 6030 7475 6086 7481
rect 6030 7415 6034 7475
rect 6115 7465 6315 7490
rect 6370 7481 6400 7669
rect 6344 7475 6400 7481
rect 6086 7415 6344 7435
rect 6396 7415 6400 7475
rect 6030 7405 6400 7415
rect 6430 7735 6800 7745
rect 6430 7675 6434 7735
rect 6486 7715 6744 7735
rect 6430 7669 6486 7675
rect 6430 7481 6460 7669
rect 6515 7660 6715 7685
rect 6796 7675 6800 7735
rect 6744 7669 6800 7675
rect 6515 7640 6585 7660
rect 6490 7600 6585 7640
rect 6645 7640 6715 7660
rect 6645 7600 6740 7640
rect 6490 7550 6740 7600
rect 6490 7510 6585 7550
rect 6515 7490 6585 7510
rect 6645 7510 6740 7550
rect 6645 7490 6715 7510
rect 6430 7475 6486 7481
rect 6430 7415 6434 7475
rect 6515 7465 6715 7490
rect 6770 7481 6800 7669
rect 6744 7475 6800 7481
rect 6486 7415 6744 7435
rect 6796 7415 6800 7475
rect 6430 7405 6800 7415
rect 6830 7735 7200 7745
rect 6830 7675 6834 7735
rect 6886 7715 7144 7735
rect 6830 7669 6886 7675
rect 6830 7481 6860 7669
rect 6915 7660 7115 7685
rect 7196 7675 7200 7735
rect 7144 7669 7200 7675
rect 6915 7640 6985 7660
rect 6890 7600 6985 7640
rect 7045 7640 7115 7660
rect 7045 7600 7140 7640
rect 6890 7550 7140 7600
rect 6890 7510 6985 7550
rect 6915 7490 6985 7510
rect 7045 7510 7140 7550
rect 7045 7490 7115 7510
rect 6830 7475 6886 7481
rect 6830 7415 6834 7475
rect 6915 7465 7115 7490
rect 7170 7481 7200 7669
rect 7144 7475 7200 7481
rect 6886 7415 7144 7435
rect 7196 7415 7200 7475
rect 6830 7405 7200 7415
rect 7230 7735 7600 7745
rect 7230 7675 7234 7735
rect 7286 7715 7544 7735
rect 7230 7669 7286 7675
rect 7230 7481 7260 7669
rect 7315 7660 7515 7685
rect 7596 7675 7600 7735
rect 7544 7669 7600 7675
rect 7315 7640 7385 7660
rect 7290 7600 7385 7640
rect 7445 7640 7515 7660
rect 7445 7600 7540 7640
rect 7290 7550 7540 7600
rect 7290 7510 7385 7550
rect 7315 7490 7385 7510
rect 7445 7510 7540 7550
rect 7445 7490 7515 7510
rect 7230 7475 7286 7481
rect 7230 7415 7234 7475
rect 7315 7465 7515 7490
rect 7570 7481 7600 7669
rect 7544 7475 7600 7481
rect 7286 7415 7544 7435
rect 7596 7415 7600 7475
rect 7230 7405 7600 7415
rect 7630 7735 8000 7745
rect 7630 7675 7634 7735
rect 7686 7715 7944 7735
rect 7630 7669 7686 7675
rect 7630 7481 7660 7669
rect 7715 7660 7915 7685
rect 7996 7675 8000 7735
rect 7944 7669 8000 7675
rect 7715 7640 7785 7660
rect 7690 7600 7785 7640
rect 7845 7640 7915 7660
rect 7845 7600 7940 7640
rect 7690 7550 7940 7600
rect 7690 7510 7785 7550
rect 7715 7490 7785 7510
rect 7845 7510 7940 7550
rect 7845 7490 7915 7510
rect 7630 7475 7686 7481
rect 7630 7415 7634 7475
rect 7715 7465 7915 7490
rect 7970 7481 8000 7669
rect 7944 7475 8000 7481
rect 7686 7415 7944 7435
rect 7996 7415 8000 7475
rect 7630 7405 8000 7415
rect 8030 7735 8400 7745
rect 8030 7675 8034 7735
rect 8086 7715 8344 7735
rect 8030 7669 8086 7675
rect 8030 7481 8060 7669
rect 8115 7660 8315 7685
rect 8396 7675 8400 7735
rect 8344 7669 8400 7675
rect 8115 7640 8185 7660
rect 8090 7600 8185 7640
rect 8245 7640 8315 7660
rect 8245 7600 8340 7640
rect 8090 7550 8340 7600
rect 8090 7510 8185 7550
rect 8115 7490 8185 7510
rect 8245 7510 8340 7550
rect 8245 7490 8315 7510
rect 8030 7475 8086 7481
rect 8030 7415 8034 7475
rect 8115 7465 8315 7490
rect 8370 7481 8400 7669
rect 8344 7475 8400 7481
rect 8086 7415 8344 7435
rect 8396 7415 8400 7475
rect 8030 7405 8400 7415
rect 8430 7735 8800 7745
rect 8430 7675 8434 7735
rect 8486 7715 8744 7735
rect 8430 7669 8486 7675
rect 8430 7481 8460 7669
rect 8515 7660 8715 7685
rect 8796 7675 8800 7735
rect 8744 7669 8800 7675
rect 8515 7640 8585 7660
rect 8490 7600 8585 7640
rect 8645 7640 8715 7660
rect 8645 7600 8740 7640
rect 8490 7550 8740 7600
rect 8490 7510 8585 7550
rect 8515 7490 8585 7510
rect 8645 7510 8740 7550
rect 8645 7490 8715 7510
rect 8430 7475 8486 7481
rect 8430 7415 8434 7475
rect 8515 7465 8715 7490
rect 8770 7481 8800 7669
rect 8744 7475 8800 7481
rect 8486 7415 8744 7435
rect 8796 7415 8800 7475
rect 8430 7405 8800 7415
rect 8830 7735 9200 7745
rect 8830 7675 8834 7735
rect 8886 7715 9144 7735
rect 8830 7669 8886 7675
rect 8830 7481 8860 7669
rect 8915 7660 9115 7685
rect 9196 7675 9200 7735
rect 9144 7669 9200 7675
rect 8915 7640 8985 7660
rect 8890 7600 8985 7640
rect 9045 7640 9115 7660
rect 9045 7600 9140 7640
rect 8890 7550 9140 7600
rect 8890 7510 8985 7550
rect 8915 7490 8985 7510
rect 9045 7510 9140 7550
rect 9045 7490 9115 7510
rect 8830 7475 8886 7481
rect 8830 7415 8834 7475
rect 8915 7465 9115 7490
rect 9170 7481 9200 7669
rect 9144 7475 9200 7481
rect 8886 7415 9144 7435
rect 9196 7415 9200 7475
rect 8830 7405 9200 7415
rect 9230 7735 9600 7745
rect 9230 7675 9234 7735
rect 9286 7715 9544 7735
rect 9230 7669 9286 7675
rect 9230 7481 9260 7669
rect 9315 7660 9515 7685
rect 9596 7675 9600 7735
rect 9544 7669 9600 7675
rect 9315 7640 9385 7660
rect 9290 7600 9385 7640
rect 9445 7640 9515 7660
rect 9445 7600 9540 7640
rect 9290 7550 9540 7600
rect 9290 7510 9385 7550
rect 9315 7490 9385 7510
rect 9445 7510 9540 7550
rect 9445 7490 9515 7510
rect 9230 7475 9286 7481
rect 9230 7415 9234 7475
rect 9315 7465 9515 7490
rect 9570 7481 9600 7669
rect 9544 7475 9600 7481
rect 9286 7415 9544 7435
rect 9596 7415 9600 7475
rect 9230 7405 9600 7415
rect 9630 7735 10000 7745
rect 9630 7675 9634 7735
rect 9686 7715 9944 7735
rect 9630 7669 9686 7675
rect 9630 7481 9660 7669
rect 9715 7660 9915 7685
rect 9996 7675 10000 7735
rect 9944 7669 10000 7675
rect 9715 7640 9785 7660
rect 9690 7600 9785 7640
rect 9845 7640 9915 7660
rect 9845 7600 9940 7640
rect 9690 7550 9940 7600
rect 9690 7510 9785 7550
rect 9715 7490 9785 7510
rect 9845 7510 9940 7550
rect 9845 7490 9915 7510
rect 9630 7475 9686 7481
rect 9630 7415 9634 7475
rect 9715 7465 9915 7490
rect 9970 7481 10000 7669
rect 9944 7475 10000 7481
rect 9686 7415 9944 7435
rect 9996 7415 10000 7475
rect 9630 7405 10000 7415
rect 10030 7735 10400 7745
rect 10030 7675 10034 7735
rect 10086 7715 10344 7735
rect 10030 7669 10086 7675
rect 10030 7481 10060 7669
rect 10115 7660 10315 7685
rect 10396 7675 10400 7735
rect 10344 7669 10400 7675
rect 10115 7640 10185 7660
rect 10090 7600 10185 7640
rect 10245 7640 10315 7660
rect 10245 7600 10340 7640
rect 10090 7550 10340 7600
rect 10090 7510 10185 7550
rect 10115 7490 10185 7510
rect 10245 7510 10340 7550
rect 10245 7490 10315 7510
rect 10030 7475 10086 7481
rect 10030 7415 10034 7475
rect 10115 7465 10315 7490
rect 10370 7481 10400 7669
rect 10344 7475 10400 7481
rect 10086 7415 10344 7435
rect 10396 7415 10400 7475
rect 10030 7405 10400 7415
rect 10430 7735 10800 7745
rect 10430 7675 10434 7735
rect 10486 7715 10744 7735
rect 10430 7669 10486 7675
rect 10430 7481 10460 7669
rect 10515 7660 10715 7685
rect 10796 7675 10800 7735
rect 10744 7669 10800 7675
rect 10515 7640 10585 7660
rect 10490 7600 10585 7640
rect 10645 7640 10715 7660
rect 10645 7600 10740 7640
rect 10490 7550 10740 7600
rect 10490 7510 10585 7550
rect 10515 7490 10585 7510
rect 10645 7510 10740 7550
rect 10645 7490 10715 7510
rect 10430 7475 10486 7481
rect 10430 7415 10434 7475
rect 10515 7465 10715 7490
rect 10770 7481 10800 7669
rect 10744 7475 10800 7481
rect 10486 7415 10744 7435
rect 10796 7415 10800 7475
rect 10430 7405 10800 7415
rect 10830 7735 11200 7745
rect 10830 7675 10834 7735
rect 10886 7715 11144 7735
rect 10830 7669 10886 7675
rect 10830 7481 10860 7669
rect 10915 7660 11115 7685
rect 11196 7675 11200 7735
rect 11144 7669 11200 7675
rect 10915 7640 10985 7660
rect 10890 7600 10985 7640
rect 11045 7640 11115 7660
rect 11045 7600 11140 7640
rect 10890 7550 11140 7600
rect 10890 7510 10985 7550
rect 10915 7490 10985 7510
rect 11045 7510 11140 7550
rect 11045 7490 11115 7510
rect 10830 7475 10886 7481
rect 10830 7415 10834 7475
rect 10915 7465 11115 7490
rect 11170 7481 11200 7669
rect 11144 7475 11200 7481
rect 10886 7415 11144 7435
rect 11196 7415 11200 7475
rect 10830 7405 11200 7415
rect 11230 7735 11600 7745
rect 11230 7675 11234 7735
rect 11286 7715 11544 7735
rect 11230 7669 11286 7675
rect 11230 7481 11260 7669
rect 11315 7660 11515 7685
rect 11596 7675 11600 7735
rect 11544 7669 11600 7675
rect 11315 7640 11385 7660
rect 11290 7600 11385 7640
rect 11445 7640 11515 7660
rect 11445 7600 11540 7640
rect 11290 7550 11540 7600
rect 11290 7510 11385 7550
rect 11315 7490 11385 7510
rect 11445 7510 11540 7550
rect 11445 7490 11515 7510
rect 11230 7475 11286 7481
rect 11230 7415 11234 7475
rect 11315 7465 11515 7490
rect 11570 7481 11600 7669
rect 11544 7475 11600 7481
rect 11286 7415 11544 7435
rect 11596 7415 11600 7475
rect 11230 7405 11600 7415
rect 11630 7735 12000 7745
rect 11630 7675 11634 7735
rect 11686 7715 11944 7735
rect 11630 7669 11686 7675
rect 11630 7481 11660 7669
rect 11715 7660 11915 7685
rect 11996 7675 12000 7735
rect 11944 7669 12000 7675
rect 11715 7640 11785 7660
rect 11690 7600 11785 7640
rect 11845 7640 11915 7660
rect 11845 7600 11940 7640
rect 11690 7550 11940 7600
rect 11690 7510 11785 7550
rect 11715 7490 11785 7510
rect 11845 7510 11940 7550
rect 11845 7490 11915 7510
rect 11630 7475 11686 7481
rect 11630 7415 11634 7475
rect 11715 7465 11915 7490
rect 11970 7481 12000 7669
rect 11944 7475 12000 7481
rect 11686 7415 11944 7435
rect 11996 7415 12000 7475
rect 11630 7405 12000 7415
rect 12030 7735 12400 7745
rect 12030 7675 12034 7735
rect 12086 7715 12344 7735
rect 12030 7669 12086 7675
rect 12030 7481 12060 7669
rect 12115 7660 12315 7685
rect 12396 7675 12400 7735
rect 12344 7669 12400 7675
rect 12115 7640 12185 7660
rect 12090 7600 12185 7640
rect 12245 7640 12315 7660
rect 12245 7600 12340 7640
rect 12090 7550 12340 7600
rect 12090 7510 12185 7550
rect 12115 7490 12185 7510
rect 12245 7510 12340 7550
rect 12245 7490 12315 7510
rect 12030 7475 12086 7481
rect 12030 7415 12034 7475
rect 12115 7465 12315 7490
rect 12370 7481 12400 7669
rect 12344 7475 12400 7481
rect 12086 7415 12344 7435
rect 12396 7415 12400 7475
rect 12030 7405 12400 7415
rect 12430 7735 12800 7745
rect 12430 7675 12434 7735
rect 12486 7715 12744 7735
rect 12430 7669 12486 7675
rect 12430 7481 12460 7669
rect 12515 7660 12715 7685
rect 12796 7675 12800 7735
rect 12744 7669 12800 7675
rect 12515 7640 12585 7660
rect 12490 7600 12585 7640
rect 12645 7640 12715 7660
rect 12645 7600 12740 7640
rect 12490 7550 12740 7600
rect 12490 7510 12585 7550
rect 12515 7490 12585 7510
rect 12645 7510 12740 7550
rect 12645 7490 12715 7510
rect 12430 7475 12486 7481
rect 12430 7415 12434 7475
rect 12515 7465 12715 7490
rect 12770 7481 12800 7669
rect 12744 7475 12800 7481
rect 12486 7415 12744 7435
rect 12796 7415 12800 7475
rect 12430 7405 12800 7415
rect 12830 7735 13200 7745
rect 12830 7675 12834 7735
rect 12886 7715 13144 7735
rect 12830 7669 12886 7675
rect 12830 7481 12860 7669
rect 12915 7660 13115 7685
rect 13196 7675 13200 7735
rect 13144 7669 13200 7675
rect 12915 7640 12985 7660
rect 12890 7600 12985 7640
rect 13045 7640 13115 7660
rect 13045 7600 13140 7640
rect 12890 7550 13140 7600
rect 12890 7510 12985 7550
rect 12915 7490 12985 7510
rect 13045 7510 13140 7550
rect 13045 7490 13115 7510
rect 12830 7475 12886 7481
rect 12830 7415 12834 7475
rect 12915 7465 13115 7490
rect 13170 7481 13200 7669
rect 13144 7475 13200 7481
rect 12886 7415 13144 7435
rect 13196 7415 13200 7475
rect 12830 7405 13200 7415
rect -370 7365 0 7375
rect -370 7305 -366 7365
rect -314 7345 -56 7365
rect -370 7299 -314 7305
rect -370 7111 -340 7299
rect -285 7290 -85 7315
rect -4 7305 0 7365
rect -56 7299 0 7305
rect -285 7270 -215 7290
rect -310 7230 -215 7270
rect -155 7270 -85 7290
rect -155 7230 -60 7270
rect -310 7180 -60 7230
rect -310 7140 -215 7180
rect -285 7120 -215 7140
rect -155 7140 -60 7180
rect -155 7120 -85 7140
rect -370 7105 -314 7111
rect -370 7045 -366 7105
rect -285 7095 -85 7120
rect -30 7111 0 7299
rect -56 7105 0 7111
rect -314 7045 -56 7065
rect -4 7045 0 7105
rect -370 7035 0 7045
rect 30 7365 400 7375
rect 30 7305 34 7365
rect 86 7345 344 7365
rect 30 7299 86 7305
rect 30 7111 60 7299
rect 115 7290 315 7315
rect 396 7305 400 7365
rect 344 7299 400 7305
rect 115 7270 185 7290
rect 90 7230 185 7270
rect 245 7270 315 7290
rect 245 7230 340 7270
rect 90 7180 340 7230
rect 90 7140 185 7180
rect 115 7120 185 7140
rect 245 7140 340 7180
rect 245 7120 315 7140
rect 30 7105 86 7111
rect 30 7045 34 7105
rect 115 7095 315 7120
rect 370 7111 400 7299
rect 344 7105 400 7111
rect 86 7045 344 7065
rect 396 7045 400 7105
rect 30 7035 400 7045
rect 430 7365 800 7375
rect 430 7305 434 7365
rect 486 7345 744 7365
rect 430 7299 486 7305
rect 430 7111 460 7299
rect 515 7290 715 7315
rect 796 7305 800 7365
rect 744 7299 800 7305
rect 515 7270 585 7290
rect 490 7230 585 7270
rect 645 7270 715 7290
rect 645 7230 740 7270
rect 490 7180 740 7230
rect 490 7140 585 7180
rect 515 7120 585 7140
rect 645 7140 740 7180
rect 645 7120 715 7140
rect 430 7105 486 7111
rect 430 7045 434 7105
rect 515 7095 715 7120
rect 770 7111 800 7299
rect 744 7105 800 7111
rect 486 7045 744 7065
rect 796 7045 800 7105
rect 430 7035 800 7045
rect 830 7365 1200 7375
rect 830 7305 834 7365
rect 886 7345 1144 7365
rect 830 7299 886 7305
rect 830 7111 860 7299
rect 915 7290 1115 7315
rect 1196 7305 1200 7365
rect 1144 7299 1200 7305
rect 915 7270 985 7290
rect 890 7230 985 7270
rect 1045 7270 1115 7290
rect 1045 7230 1140 7270
rect 890 7180 1140 7230
rect 890 7140 985 7180
rect 915 7120 985 7140
rect 1045 7140 1140 7180
rect 1045 7120 1115 7140
rect 830 7105 886 7111
rect 830 7045 834 7105
rect 915 7095 1115 7120
rect 1170 7111 1200 7299
rect 1144 7105 1200 7111
rect 886 7045 1144 7065
rect 1196 7045 1200 7105
rect 830 7035 1200 7045
rect 1230 7365 1600 7375
rect 1230 7305 1234 7365
rect 1286 7345 1544 7365
rect 1230 7299 1286 7305
rect 1230 7111 1260 7299
rect 1315 7290 1515 7315
rect 1596 7305 1600 7365
rect 1544 7299 1600 7305
rect 1315 7270 1385 7290
rect 1290 7230 1385 7270
rect 1445 7270 1515 7290
rect 1445 7230 1540 7270
rect 1290 7180 1540 7230
rect 1290 7140 1385 7180
rect 1315 7120 1385 7140
rect 1445 7140 1540 7180
rect 1445 7120 1515 7140
rect 1230 7105 1286 7111
rect 1230 7045 1234 7105
rect 1315 7095 1515 7120
rect 1570 7111 1600 7299
rect 1544 7105 1600 7111
rect 1286 7045 1544 7065
rect 1596 7045 1600 7105
rect 1230 7035 1600 7045
rect 1630 7365 2000 7375
rect 1630 7305 1634 7365
rect 1686 7345 1944 7365
rect 1630 7299 1686 7305
rect 1630 7111 1660 7299
rect 1715 7290 1915 7315
rect 1996 7305 2000 7365
rect 1944 7299 2000 7305
rect 1715 7270 1785 7290
rect 1690 7230 1785 7270
rect 1845 7270 1915 7290
rect 1845 7230 1940 7270
rect 1690 7180 1940 7230
rect 1690 7140 1785 7180
rect 1715 7120 1785 7140
rect 1845 7140 1940 7180
rect 1845 7120 1915 7140
rect 1630 7105 1686 7111
rect 1630 7045 1634 7105
rect 1715 7095 1915 7120
rect 1970 7111 2000 7299
rect 1944 7105 2000 7111
rect 1686 7045 1944 7065
rect 1996 7045 2000 7105
rect 1630 7035 2000 7045
rect 2030 7365 2400 7375
rect 2030 7305 2034 7365
rect 2086 7345 2344 7365
rect 2030 7299 2086 7305
rect 2030 7111 2060 7299
rect 2115 7290 2315 7315
rect 2396 7305 2400 7365
rect 2344 7299 2400 7305
rect 2115 7270 2185 7290
rect 2090 7230 2185 7270
rect 2245 7270 2315 7290
rect 2245 7230 2340 7270
rect 2090 7180 2340 7230
rect 2090 7140 2185 7180
rect 2115 7120 2185 7140
rect 2245 7140 2340 7180
rect 2245 7120 2315 7140
rect 2030 7105 2086 7111
rect 2030 7045 2034 7105
rect 2115 7095 2315 7120
rect 2370 7111 2400 7299
rect 2344 7105 2400 7111
rect 2086 7045 2344 7065
rect 2396 7045 2400 7105
rect 2030 7035 2400 7045
rect 2430 7365 2800 7375
rect 2430 7305 2434 7365
rect 2486 7345 2744 7365
rect 2430 7299 2486 7305
rect 2430 7111 2460 7299
rect 2515 7290 2715 7315
rect 2796 7305 2800 7365
rect 2744 7299 2800 7305
rect 2515 7270 2585 7290
rect 2490 7230 2585 7270
rect 2645 7270 2715 7290
rect 2645 7230 2740 7270
rect 2490 7180 2740 7230
rect 2490 7140 2585 7180
rect 2515 7120 2585 7140
rect 2645 7140 2740 7180
rect 2645 7120 2715 7140
rect 2430 7105 2486 7111
rect 2430 7045 2434 7105
rect 2515 7095 2715 7120
rect 2770 7111 2800 7299
rect 2744 7105 2800 7111
rect 2486 7045 2744 7065
rect 2796 7045 2800 7105
rect 2430 7035 2800 7045
rect 2830 7365 3200 7375
rect 2830 7305 2834 7365
rect 2886 7345 3144 7365
rect 2830 7299 2886 7305
rect 2830 7111 2860 7299
rect 2915 7290 3115 7315
rect 3196 7305 3200 7365
rect 3144 7299 3200 7305
rect 2915 7270 2985 7290
rect 2890 7230 2985 7270
rect 3045 7270 3115 7290
rect 3045 7230 3140 7270
rect 2890 7180 3140 7230
rect 2890 7140 2985 7180
rect 2915 7120 2985 7140
rect 3045 7140 3140 7180
rect 3045 7120 3115 7140
rect 2830 7105 2886 7111
rect 2830 7045 2834 7105
rect 2915 7095 3115 7120
rect 3170 7111 3200 7299
rect 3144 7105 3200 7111
rect 2886 7045 3144 7065
rect 3196 7045 3200 7105
rect 2830 7035 3200 7045
rect 3230 7365 3600 7375
rect 3230 7305 3234 7365
rect 3286 7345 3544 7365
rect 3230 7299 3286 7305
rect 3230 7111 3260 7299
rect 3315 7290 3515 7315
rect 3596 7305 3600 7365
rect 3544 7299 3600 7305
rect 3315 7270 3385 7290
rect 3290 7230 3385 7270
rect 3445 7270 3515 7290
rect 3445 7230 3540 7270
rect 3290 7180 3540 7230
rect 3290 7140 3385 7180
rect 3315 7120 3385 7140
rect 3445 7140 3540 7180
rect 3445 7120 3515 7140
rect 3230 7105 3286 7111
rect 3230 7045 3234 7105
rect 3315 7095 3515 7120
rect 3570 7111 3600 7299
rect 3544 7105 3600 7111
rect 3286 7045 3544 7065
rect 3596 7045 3600 7105
rect 3230 7035 3600 7045
rect 3630 7365 4000 7375
rect 3630 7305 3634 7365
rect 3686 7345 3944 7365
rect 3630 7299 3686 7305
rect 3630 7111 3660 7299
rect 3715 7290 3915 7315
rect 3996 7305 4000 7365
rect 3944 7299 4000 7305
rect 3715 7270 3785 7290
rect 3690 7230 3785 7270
rect 3845 7270 3915 7290
rect 3845 7230 3940 7270
rect 3690 7180 3940 7230
rect 3690 7140 3785 7180
rect 3715 7120 3785 7140
rect 3845 7140 3940 7180
rect 3845 7120 3915 7140
rect 3630 7105 3686 7111
rect 3630 7045 3634 7105
rect 3715 7095 3915 7120
rect 3970 7111 4000 7299
rect 3944 7105 4000 7111
rect 3686 7045 3944 7065
rect 3996 7045 4000 7105
rect 3630 7035 4000 7045
rect 4030 7365 4400 7375
rect 4030 7305 4034 7365
rect 4086 7345 4344 7365
rect 4030 7299 4086 7305
rect 4030 7111 4060 7299
rect 4115 7290 4315 7315
rect 4396 7305 4400 7365
rect 4344 7299 4400 7305
rect 4115 7270 4185 7290
rect 4090 7230 4185 7270
rect 4245 7270 4315 7290
rect 4245 7230 4340 7270
rect 4090 7180 4340 7230
rect 4090 7140 4185 7180
rect 4115 7120 4185 7140
rect 4245 7140 4340 7180
rect 4245 7120 4315 7140
rect 4030 7105 4086 7111
rect 4030 7045 4034 7105
rect 4115 7095 4315 7120
rect 4370 7111 4400 7299
rect 4344 7105 4400 7111
rect 4086 7045 4344 7065
rect 4396 7045 4400 7105
rect 4030 7035 4400 7045
rect 4430 7365 4800 7375
rect 4430 7305 4434 7365
rect 4486 7345 4744 7365
rect 4430 7299 4486 7305
rect 4430 7111 4460 7299
rect 4515 7290 4715 7315
rect 4796 7305 4800 7365
rect 4744 7299 4800 7305
rect 4515 7270 4585 7290
rect 4490 7230 4585 7270
rect 4645 7270 4715 7290
rect 4645 7230 4740 7270
rect 4490 7180 4740 7230
rect 4490 7140 4585 7180
rect 4515 7120 4585 7140
rect 4645 7140 4740 7180
rect 4645 7120 4715 7140
rect 4430 7105 4486 7111
rect 4430 7045 4434 7105
rect 4515 7095 4715 7120
rect 4770 7111 4800 7299
rect 4744 7105 4800 7111
rect 4486 7045 4744 7065
rect 4796 7045 4800 7105
rect 4430 7035 4800 7045
rect 4830 7365 5200 7375
rect 4830 7305 4834 7365
rect 4886 7345 5144 7365
rect 4830 7299 4886 7305
rect 4830 7111 4860 7299
rect 4915 7290 5115 7315
rect 5196 7305 5200 7365
rect 5144 7299 5200 7305
rect 4915 7270 4985 7290
rect 4890 7230 4985 7270
rect 5045 7270 5115 7290
rect 5045 7230 5140 7270
rect 4890 7180 5140 7230
rect 4890 7140 4985 7180
rect 4915 7120 4985 7140
rect 5045 7140 5140 7180
rect 5045 7120 5115 7140
rect 4830 7105 4886 7111
rect 4830 7045 4834 7105
rect 4915 7095 5115 7120
rect 5170 7111 5200 7299
rect 5144 7105 5200 7111
rect 4886 7045 5144 7065
rect 5196 7045 5200 7105
rect 4830 7035 5200 7045
rect 5230 7365 5600 7375
rect 5230 7305 5234 7365
rect 5286 7345 5544 7365
rect 5230 7299 5286 7305
rect 5230 7111 5260 7299
rect 5315 7290 5515 7315
rect 5596 7305 5600 7365
rect 5544 7299 5600 7305
rect 5315 7270 5385 7290
rect 5290 7230 5385 7270
rect 5445 7270 5515 7290
rect 5445 7230 5540 7270
rect 5290 7180 5540 7230
rect 5290 7140 5385 7180
rect 5315 7120 5385 7140
rect 5445 7140 5540 7180
rect 5445 7120 5515 7140
rect 5230 7105 5286 7111
rect 5230 7045 5234 7105
rect 5315 7095 5515 7120
rect 5570 7111 5600 7299
rect 5544 7105 5600 7111
rect 5286 7045 5544 7065
rect 5596 7045 5600 7105
rect 5230 7035 5600 7045
rect 5630 7365 6000 7375
rect 5630 7305 5634 7365
rect 5686 7345 5944 7365
rect 5630 7299 5686 7305
rect 5630 7111 5660 7299
rect 5715 7290 5915 7315
rect 5996 7305 6000 7365
rect 5944 7299 6000 7305
rect 5715 7270 5785 7290
rect 5690 7230 5785 7270
rect 5845 7270 5915 7290
rect 5845 7230 5940 7270
rect 5690 7180 5940 7230
rect 5690 7140 5785 7180
rect 5715 7120 5785 7140
rect 5845 7140 5940 7180
rect 5845 7120 5915 7140
rect 5630 7105 5686 7111
rect 5630 7045 5634 7105
rect 5715 7095 5915 7120
rect 5970 7111 6000 7299
rect 5944 7105 6000 7111
rect 5686 7045 5944 7065
rect 5996 7045 6000 7105
rect 5630 7035 6000 7045
rect 6030 7365 6400 7375
rect 6030 7305 6034 7365
rect 6086 7345 6344 7365
rect 6030 7299 6086 7305
rect 6030 7111 6060 7299
rect 6115 7290 6315 7315
rect 6396 7305 6400 7365
rect 6344 7299 6400 7305
rect 6115 7270 6185 7290
rect 6090 7230 6185 7270
rect 6245 7270 6315 7290
rect 6245 7230 6340 7270
rect 6090 7180 6340 7230
rect 6090 7140 6185 7180
rect 6115 7120 6185 7140
rect 6245 7140 6340 7180
rect 6245 7120 6315 7140
rect 6030 7105 6086 7111
rect 6030 7045 6034 7105
rect 6115 7095 6315 7120
rect 6370 7111 6400 7299
rect 6344 7105 6400 7111
rect 6086 7045 6344 7065
rect 6396 7045 6400 7105
rect 6030 7035 6400 7045
rect 6430 7365 6800 7375
rect 6430 7305 6434 7365
rect 6486 7345 6744 7365
rect 6430 7299 6486 7305
rect 6430 7111 6460 7299
rect 6515 7290 6715 7315
rect 6796 7305 6800 7365
rect 6744 7299 6800 7305
rect 6515 7270 6585 7290
rect 6490 7230 6585 7270
rect 6645 7270 6715 7290
rect 6645 7230 6740 7270
rect 6490 7180 6740 7230
rect 6490 7140 6585 7180
rect 6515 7120 6585 7140
rect 6645 7140 6740 7180
rect 6645 7120 6715 7140
rect 6430 7105 6486 7111
rect 6430 7045 6434 7105
rect 6515 7095 6715 7120
rect 6770 7111 6800 7299
rect 6744 7105 6800 7111
rect 6486 7045 6744 7065
rect 6796 7045 6800 7105
rect 6430 7035 6800 7045
rect 6830 7365 7200 7375
rect 6830 7305 6834 7365
rect 6886 7345 7144 7365
rect 6830 7299 6886 7305
rect 6830 7111 6860 7299
rect 6915 7290 7115 7315
rect 7196 7305 7200 7365
rect 7144 7299 7200 7305
rect 6915 7270 6985 7290
rect 6890 7230 6985 7270
rect 7045 7270 7115 7290
rect 7045 7230 7140 7270
rect 6890 7180 7140 7230
rect 6890 7140 6985 7180
rect 6915 7120 6985 7140
rect 7045 7140 7140 7180
rect 7045 7120 7115 7140
rect 6830 7105 6886 7111
rect 6830 7045 6834 7105
rect 6915 7095 7115 7120
rect 7170 7111 7200 7299
rect 7144 7105 7200 7111
rect 6886 7045 7144 7065
rect 7196 7045 7200 7105
rect 6830 7035 7200 7045
rect 7230 7365 7600 7375
rect 7230 7305 7234 7365
rect 7286 7345 7544 7365
rect 7230 7299 7286 7305
rect 7230 7111 7260 7299
rect 7315 7290 7515 7315
rect 7596 7305 7600 7365
rect 7544 7299 7600 7305
rect 7315 7270 7385 7290
rect 7290 7230 7385 7270
rect 7445 7270 7515 7290
rect 7445 7230 7540 7270
rect 7290 7180 7540 7230
rect 7290 7140 7385 7180
rect 7315 7120 7385 7140
rect 7445 7140 7540 7180
rect 7445 7120 7515 7140
rect 7230 7105 7286 7111
rect 7230 7045 7234 7105
rect 7315 7095 7515 7120
rect 7570 7111 7600 7299
rect 7544 7105 7600 7111
rect 7286 7045 7544 7065
rect 7596 7045 7600 7105
rect 7230 7035 7600 7045
rect 7630 7365 8000 7375
rect 7630 7305 7634 7365
rect 7686 7345 7944 7365
rect 7630 7299 7686 7305
rect 7630 7111 7660 7299
rect 7715 7290 7915 7315
rect 7996 7305 8000 7365
rect 7944 7299 8000 7305
rect 7715 7270 7785 7290
rect 7690 7230 7785 7270
rect 7845 7270 7915 7290
rect 7845 7230 7940 7270
rect 7690 7180 7940 7230
rect 7690 7140 7785 7180
rect 7715 7120 7785 7140
rect 7845 7140 7940 7180
rect 7845 7120 7915 7140
rect 7630 7105 7686 7111
rect 7630 7045 7634 7105
rect 7715 7095 7915 7120
rect 7970 7111 8000 7299
rect 7944 7105 8000 7111
rect 7686 7045 7944 7065
rect 7996 7045 8000 7105
rect 7630 7035 8000 7045
rect 8030 7365 8400 7375
rect 8030 7305 8034 7365
rect 8086 7345 8344 7365
rect 8030 7299 8086 7305
rect 8030 7111 8060 7299
rect 8115 7290 8315 7315
rect 8396 7305 8400 7365
rect 8344 7299 8400 7305
rect 8115 7270 8185 7290
rect 8090 7230 8185 7270
rect 8245 7270 8315 7290
rect 8245 7230 8340 7270
rect 8090 7180 8340 7230
rect 8090 7140 8185 7180
rect 8115 7120 8185 7140
rect 8245 7140 8340 7180
rect 8245 7120 8315 7140
rect 8030 7105 8086 7111
rect 8030 7045 8034 7105
rect 8115 7095 8315 7120
rect 8370 7111 8400 7299
rect 8344 7105 8400 7111
rect 8086 7045 8344 7065
rect 8396 7045 8400 7105
rect 8030 7035 8400 7045
rect 8430 7365 8800 7375
rect 8430 7305 8434 7365
rect 8486 7345 8744 7365
rect 8430 7299 8486 7305
rect 8430 7111 8460 7299
rect 8515 7290 8715 7315
rect 8796 7305 8800 7365
rect 8744 7299 8800 7305
rect 8515 7270 8585 7290
rect 8490 7230 8585 7270
rect 8645 7270 8715 7290
rect 8645 7230 8740 7270
rect 8490 7180 8740 7230
rect 8490 7140 8585 7180
rect 8515 7120 8585 7140
rect 8645 7140 8740 7180
rect 8645 7120 8715 7140
rect 8430 7105 8486 7111
rect 8430 7045 8434 7105
rect 8515 7095 8715 7120
rect 8770 7111 8800 7299
rect 8744 7105 8800 7111
rect 8486 7045 8744 7065
rect 8796 7045 8800 7105
rect 8430 7035 8800 7045
rect 8830 7365 9200 7375
rect 8830 7305 8834 7365
rect 8886 7345 9144 7365
rect 8830 7299 8886 7305
rect 8830 7111 8860 7299
rect 8915 7290 9115 7315
rect 9196 7305 9200 7365
rect 9144 7299 9200 7305
rect 8915 7270 8985 7290
rect 8890 7230 8985 7270
rect 9045 7270 9115 7290
rect 9045 7230 9140 7270
rect 8890 7180 9140 7230
rect 8890 7140 8985 7180
rect 8915 7120 8985 7140
rect 9045 7140 9140 7180
rect 9045 7120 9115 7140
rect 8830 7105 8886 7111
rect 8830 7045 8834 7105
rect 8915 7095 9115 7120
rect 9170 7111 9200 7299
rect 9144 7105 9200 7111
rect 8886 7045 9144 7065
rect 9196 7045 9200 7105
rect 8830 7035 9200 7045
rect 9230 7365 9600 7375
rect 9230 7305 9234 7365
rect 9286 7345 9544 7365
rect 9230 7299 9286 7305
rect 9230 7111 9260 7299
rect 9315 7290 9515 7315
rect 9596 7305 9600 7365
rect 9544 7299 9600 7305
rect 9315 7270 9385 7290
rect 9290 7230 9385 7270
rect 9445 7270 9515 7290
rect 9445 7230 9540 7270
rect 9290 7180 9540 7230
rect 9290 7140 9385 7180
rect 9315 7120 9385 7140
rect 9445 7140 9540 7180
rect 9445 7120 9515 7140
rect 9230 7105 9286 7111
rect 9230 7045 9234 7105
rect 9315 7095 9515 7120
rect 9570 7111 9600 7299
rect 9544 7105 9600 7111
rect 9286 7045 9544 7065
rect 9596 7045 9600 7105
rect 9230 7035 9600 7045
rect 9630 7365 10000 7375
rect 9630 7305 9634 7365
rect 9686 7345 9944 7365
rect 9630 7299 9686 7305
rect 9630 7111 9660 7299
rect 9715 7290 9915 7315
rect 9996 7305 10000 7365
rect 9944 7299 10000 7305
rect 9715 7270 9785 7290
rect 9690 7230 9785 7270
rect 9845 7270 9915 7290
rect 9845 7230 9940 7270
rect 9690 7180 9940 7230
rect 9690 7140 9785 7180
rect 9715 7120 9785 7140
rect 9845 7140 9940 7180
rect 9845 7120 9915 7140
rect 9630 7105 9686 7111
rect 9630 7045 9634 7105
rect 9715 7095 9915 7120
rect 9970 7111 10000 7299
rect 9944 7105 10000 7111
rect 9686 7045 9944 7065
rect 9996 7045 10000 7105
rect 9630 7035 10000 7045
rect 10030 7365 10400 7375
rect 10030 7305 10034 7365
rect 10086 7345 10344 7365
rect 10030 7299 10086 7305
rect 10030 7111 10060 7299
rect 10115 7290 10315 7315
rect 10396 7305 10400 7365
rect 10344 7299 10400 7305
rect 10115 7270 10185 7290
rect 10090 7230 10185 7270
rect 10245 7270 10315 7290
rect 10245 7230 10340 7270
rect 10090 7180 10340 7230
rect 10090 7140 10185 7180
rect 10115 7120 10185 7140
rect 10245 7140 10340 7180
rect 10245 7120 10315 7140
rect 10030 7105 10086 7111
rect 10030 7045 10034 7105
rect 10115 7095 10315 7120
rect 10370 7111 10400 7299
rect 10344 7105 10400 7111
rect 10086 7045 10344 7065
rect 10396 7045 10400 7105
rect 10030 7035 10400 7045
rect 10430 7365 10800 7375
rect 10430 7305 10434 7365
rect 10486 7345 10744 7365
rect 10430 7299 10486 7305
rect 10430 7111 10460 7299
rect 10515 7290 10715 7315
rect 10796 7305 10800 7365
rect 10744 7299 10800 7305
rect 10515 7270 10585 7290
rect 10490 7230 10585 7270
rect 10645 7270 10715 7290
rect 10645 7230 10740 7270
rect 10490 7180 10740 7230
rect 10490 7140 10585 7180
rect 10515 7120 10585 7140
rect 10645 7140 10740 7180
rect 10645 7120 10715 7140
rect 10430 7105 10486 7111
rect 10430 7045 10434 7105
rect 10515 7095 10715 7120
rect 10770 7111 10800 7299
rect 10744 7105 10800 7111
rect 10486 7045 10744 7065
rect 10796 7045 10800 7105
rect 10430 7035 10800 7045
rect 10830 7365 11200 7375
rect 10830 7305 10834 7365
rect 10886 7345 11144 7365
rect 10830 7299 10886 7305
rect 10830 7111 10860 7299
rect 10915 7290 11115 7315
rect 11196 7305 11200 7365
rect 11144 7299 11200 7305
rect 10915 7270 10985 7290
rect 10890 7230 10985 7270
rect 11045 7270 11115 7290
rect 11045 7230 11140 7270
rect 10890 7180 11140 7230
rect 10890 7140 10985 7180
rect 10915 7120 10985 7140
rect 11045 7140 11140 7180
rect 11045 7120 11115 7140
rect 10830 7105 10886 7111
rect 10830 7045 10834 7105
rect 10915 7095 11115 7120
rect 11170 7111 11200 7299
rect 11144 7105 11200 7111
rect 10886 7045 11144 7065
rect 11196 7045 11200 7105
rect 10830 7035 11200 7045
rect 11230 7365 11600 7375
rect 11230 7305 11234 7365
rect 11286 7345 11544 7365
rect 11230 7299 11286 7305
rect 11230 7111 11260 7299
rect 11315 7290 11515 7315
rect 11596 7305 11600 7365
rect 11544 7299 11600 7305
rect 11315 7270 11385 7290
rect 11290 7230 11385 7270
rect 11445 7270 11515 7290
rect 11445 7230 11540 7270
rect 11290 7180 11540 7230
rect 11290 7140 11385 7180
rect 11315 7120 11385 7140
rect 11445 7140 11540 7180
rect 11445 7120 11515 7140
rect 11230 7105 11286 7111
rect 11230 7045 11234 7105
rect 11315 7095 11515 7120
rect 11570 7111 11600 7299
rect 11544 7105 11600 7111
rect 11286 7045 11544 7065
rect 11596 7045 11600 7105
rect 11230 7035 11600 7045
rect 11630 7365 12000 7375
rect 11630 7305 11634 7365
rect 11686 7345 11944 7365
rect 11630 7299 11686 7305
rect 11630 7111 11660 7299
rect 11715 7290 11915 7315
rect 11996 7305 12000 7365
rect 11944 7299 12000 7305
rect 11715 7270 11785 7290
rect 11690 7230 11785 7270
rect 11845 7270 11915 7290
rect 11845 7230 11940 7270
rect 11690 7180 11940 7230
rect 11690 7140 11785 7180
rect 11715 7120 11785 7140
rect 11845 7140 11940 7180
rect 11845 7120 11915 7140
rect 11630 7105 11686 7111
rect 11630 7045 11634 7105
rect 11715 7095 11915 7120
rect 11970 7111 12000 7299
rect 11944 7105 12000 7111
rect 11686 7045 11944 7065
rect 11996 7045 12000 7105
rect 11630 7035 12000 7045
rect 12030 7365 12400 7375
rect 12030 7305 12034 7365
rect 12086 7345 12344 7365
rect 12030 7299 12086 7305
rect 12030 7111 12060 7299
rect 12115 7290 12315 7315
rect 12396 7305 12400 7365
rect 12344 7299 12400 7305
rect 12115 7270 12185 7290
rect 12090 7230 12185 7270
rect 12245 7270 12315 7290
rect 12245 7230 12340 7270
rect 12090 7180 12340 7230
rect 12090 7140 12185 7180
rect 12115 7120 12185 7140
rect 12245 7140 12340 7180
rect 12245 7120 12315 7140
rect 12030 7105 12086 7111
rect 12030 7045 12034 7105
rect 12115 7095 12315 7120
rect 12370 7111 12400 7299
rect 12344 7105 12400 7111
rect 12086 7045 12344 7065
rect 12396 7045 12400 7105
rect 12030 7035 12400 7045
rect 12430 7365 12800 7375
rect 12430 7305 12434 7365
rect 12486 7345 12744 7365
rect 12430 7299 12486 7305
rect 12430 7111 12460 7299
rect 12515 7290 12715 7315
rect 12796 7305 12800 7365
rect 12744 7299 12800 7305
rect 12515 7270 12585 7290
rect 12490 7230 12585 7270
rect 12645 7270 12715 7290
rect 12645 7230 12740 7270
rect 12490 7180 12740 7230
rect 12490 7140 12585 7180
rect 12515 7120 12585 7140
rect 12645 7140 12740 7180
rect 12645 7120 12715 7140
rect 12430 7105 12486 7111
rect 12430 7045 12434 7105
rect 12515 7095 12715 7120
rect 12770 7111 12800 7299
rect 12744 7105 12800 7111
rect 12486 7045 12744 7065
rect 12796 7045 12800 7105
rect 12430 7035 12800 7045
rect 12830 7365 13200 7375
rect 12830 7305 12834 7365
rect 12886 7345 13144 7365
rect 12830 7299 12886 7305
rect 12830 7111 12860 7299
rect 12915 7290 13115 7315
rect 13196 7305 13200 7365
rect 13144 7299 13200 7305
rect 12915 7270 12985 7290
rect 12890 7230 12985 7270
rect 13045 7270 13115 7290
rect 13045 7230 13140 7270
rect 12890 7180 13140 7230
rect 12890 7140 12985 7180
rect 12915 7120 12985 7140
rect 13045 7140 13140 7180
rect 13045 7120 13115 7140
rect 12830 7105 12886 7111
rect 12830 7045 12834 7105
rect 12915 7095 13115 7120
rect 13170 7111 13200 7299
rect 13144 7105 13200 7111
rect 12886 7045 13144 7065
rect 13196 7045 13200 7105
rect 12830 7035 13200 7045
rect -370 6995 0 7005
rect -370 6935 -366 6995
rect -314 6975 -56 6995
rect -370 6929 -314 6935
rect -370 6741 -340 6929
rect -285 6920 -85 6945
rect -4 6935 0 6995
rect -56 6929 0 6935
rect -285 6900 -215 6920
rect -310 6860 -215 6900
rect -155 6900 -85 6920
rect -155 6860 -60 6900
rect -310 6810 -60 6860
rect -310 6770 -215 6810
rect -285 6750 -215 6770
rect -155 6770 -60 6810
rect -155 6750 -85 6770
rect -370 6735 -314 6741
rect -370 6675 -366 6735
rect -285 6725 -85 6750
rect -30 6741 0 6929
rect -56 6735 0 6741
rect -314 6675 -56 6695
rect -4 6675 0 6735
rect -370 6665 0 6675
rect 30 6995 400 7005
rect 30 6935 34 6995
rect 86 6975 344 6995
rect 30 6929 86 6935
rect 30 6741 60 6929
rect 115 6920 315 6945
rect 396 6935 400 6995
rect 344 6929 400 6935
rect 115 6900 185 6920
rect 90 6860 185 6900
rect 245 6900 315 6920
rect 245 6860 340 6900
rect 90 6810 340 6860
rect 90 6770 185 6810
rect 115 6750 185 6770
rect 245 6770 340 6810
rect 245 6750 315 6770
rect 30 6735 86 6741
rect 30 6675 34 6735
rect 115 6725 315 6750
rect 370 6741 400 6929
rect 344 6735 400 6741
rect 86 6675 344 6695
rect 396 6675 400 6735
rect 30 6665 400 6675
rect 430 6995 800 7005
rect 430 6935 434 6995
rect 486 6975 744 6995
rect 430 6929 486 6935
rect 430 6741 460 6929
rect 515 6920 715 6945
rect 796 6935 800 6995
rect 744 6929 800 6935
rect 515 6900 585 6920
rect 490 6860 585 6900
rect 645 6900 715 6920
rect 645 6860 740 6900
rect 490 6810 740 6860
rect 490 6770 585 6810
rect 515 6750 585 6770
rect 645 6770 740 6810
rect 645 6750 715 6770
rect 430 6735 486 6741
rect 430 6675 434 6735
rect 515 6725 715 6750
rect 770 6741 800 6929
rect 744 6735 800 6741
rect 486 6675 744 6695
rect 796 6675 800 6735
rect 430 6665 800 6675
rect 830 6995 1200 7005
rect 830 6935 834 6995
rect 886 6975 1144 6995
rect 830 6929 886 6935
rect 830 6741 860 6929
rect 915 6920 1115 6945
rect 1196 6935 1200 6995
rect 1144 6929 1200 6935
rect 915 6900 985 6920
rect 890 6860 985 6900
rect 1045 6900 1115 6920
rect 1045 6860 1140 6900
rect 890 6810 1140 6860
rect 890 6770 985 6810
rect 915 6750 985 6770
rect 1045 6770 1140 6810
rect 1045 6750 1115 6770
rect 830 6735 886 6741
rect 830 6675 834 6735
rect 915 6725 1115 6750
rect 1170 6741 1200 6929
rect 1144 6735 1200 6741
rect 886 6675 1144 6695
rect 1196 6675 1200 6735
rect 830 6665 1200 6675
rect 1230 6995 1600 7005
rect 1230 6935 1234 6995
rect 1286 6975 1544 6995
rect 1230 6929 1286 6935
rect 1230 6741 1260 6929
rect 1315 6920 1515 6945
rect 1596 6935 1600 6995
rect 1544 6929 1600 6935
rect 1315 6900 1385 6920
rect 1290 6860 1385 6900
rect 1445 6900 1515 6920
rect 1445 6860 1540 6900
rect 1290 6810 1540 6860
rect 1290 6770 1385 6810
rect 1315 6750 1385 6770
rect 1445 6770 1540 6810
rect 1445 6750 1515 6770
rect 1230 6735 1286 6741
rect 1230 6675 1234 6735
rect 1315 6725 1515 6750
rect 1570 6741 1600 6929
rect 1544 6735 1600 6741
rect 1286 6675 1544 6695
rect 1596 6675 1600 6735
rect 1230 6665 1600 6675
rect 1630 6995 2000 7005
rect 1630 6935 1634 6995
rect 1686 6975 1944 6995
rect 1630 6929 1686 6935
rect 1630 6741 1660 6929
rect 1715 6920 1915 6945
rect 1996 6935 2000 6995
rect 1944 6929 2000 6935
rect 1715 6900 1785 6920
rect 1690 6860 1785 6900
rect 1845 6900 1915 6920
rect 1845 6860 1940 6900
rect 1690 6810 1940 6860
rect 1690 6770 1785 6810
rect 1715 6750 1785 6770
rect 1845 6770 1940 6810
rect 1845 6750 1915 6770
rect 1630 6735 1686 6741
rect 1630 6675 1634 6735
rect 1715 6725 1915 6750
rect 1970 6741 2000 6929
rect 1944 6735 2000 6741
rect 1686 6675 1944 6695
rect 1996 6675 2000 6735
rect 1630 6665 2000 6675
rect 2030 6995 2400 7005
rect 2030 6935 2034 6995
rect 2086 6975 2344 6995
rect 2030 6929 2086 6935
rect 2030 6741 2060 6929
rect 2115 6920 2315 6945
rect 2396 6935 2400 6995
rect 2344 6929 2400 6935
rect 2115 6900 2185 6920
rect 2090 6860 2185 6900
rect 2245 6900 2315 6920
rect 2245 6860 2340 6900
rect 2090 6810 2340 6860
rect 2090 6770 2185 6810
rect 2115 6750 2185 6770
rect 2245 6770 2340 6810
rect 2245 6750 2315 6770
rect 2030 6735 2086 6741
rect 2030 6675 2034 6735
rect 2115 6725 2315 6750
rect 2370 6741 2400 6929
rect 2344 6735 2400 6741
rect 2086 6675 2344 6695
rect 2396 6675 2400 6735
rect 2030 6665 2400 6675
rect 2430 6995 2800 7005
rect 2430 6935 2434 6995
rect 2486 6975 2744 6995
rect 2430 6929 2486 6935
rect 2430 6741 2460 6929
rect 2515 6920 2715 6945
rect 2796 6935 2800 6995
rect 2744 6929 2800 6935
rect 2515 6900 2585 6920
rect 2490 6860 2585 6900
rect 2645 6900 2715 6920
rect 2645 6860 2740 6900
rect 2490 6810 2740 6860
rect 2490 6770 2585 6810
rect 2515 6750 2585 6770
rect 2645 6770 2740 6810
rect 2645 6750 2715 6770
rect 2430 6735 2486 6741
rect 2430 6675 2434 6735
rect 2515 6725 2715 6750
rect 2770 6741 2800 6929
rect 2744 6735 2800 6741
rect 2486 6675 2744 6695
rect 2796 6675 2800 6735
rect 2430 6665 2800 6675
rect 2830 6995 3200 7005
rect 2830 6935 2834 6995
rect 2886 6975 3144 6995
rect 2830 6929 2886 6935
rect 2830 6741 2860 6929
rect 2915 6920 3115 6945
rect 3196 6935 3200 6995
rect 3144 6929 3200 6935
rect 2915 6900 2985 6920
rect 2890 6860 2985 6900
rect 3045 6900 3115 6920
rect 3045 6860 3140 6900
rect 2890 6810 3140 6860
rect 2890 6770 2985 6810
rect 2915 6750 2985 6770
rect 3045 6770 3140 6810
rect 3045 6750 3115 6770
rect 2830 6735 2886 6741
rect 2830 6675 2834 6735
rect 2915 6725 3115 6750
rect 3170 6741 3200 6929
rect 3144 6735 3200 6741
rect 2886 6675 3144 6695
rect 3196 6675 3200 6735
rect 2830 6665 3200 6675
rect 3230 6995 3600 7005
rect 3230 6935 3234 6995
rect 3286 6975 3544 6995
rect 3230 6929 3286 6935
rect 3230 6741 3260 6929
rect 3315 6920 3515 6945
rect 3596 6935 3600 6995
rect 3544 6929 3600 6935
rect 3315 6900 3385 6920
rect 3290 6860 3385 6900
rect 3445 6900 3515 6920
rect 3445 6860 3540 6900
rect 3290 6810 3540 6860
rect 3290 6770 3385 6810
rect 3315 6750 3385 6770
rect 3445 6770 3540 6810
rect 3445 6750 3515 6770
rect 3230 6735 3286 6741
rect 3230 6675 3234 6735
rect 3315 6725 3515 6750
rect 3570 6741 3600 6929
rect 3544 6735 3600 6741
rect 3286 6675 3544 6695
rect 3596 6675 3600 6735
rect 3230 6665 3600 6675
rect 3630 6995 4000 7005
rect 3630 6935 3634 6995
rect 3686 6975 3944 6995
rect 3630 6929 3686 6935
rect 3630 6741 3660 6929
rect 3715 6920 3915 6945
rect 3996 6935 4000 6995
rect 3944 6929 4000 6935
rect 3715 6900 3785 6920
rect 3690 6860 3785 6900
rect 3845 6900 3915 6920
rect 3845 6860 3940 6900
rect 3690 6810 3940 6860
rect 3690 6770 3785 6810
rect 3715 6750 3785 6770
rect 3845 6770 3940 6810
rect 3845 6750 3915 6770
rect 3630 6735 3686 6741
rect 3630 6675 3634 6735
rect 3715 6725 3915 6750
rect 3970 6741 4000 6929
rect 3944 6735 4000 6741
rect 3686 6675 3944 6695
rect 3996 6675 4000 6735
rect 3630 6665 4000 6675
rect 4030 6995 4400 7005
rect 4030 6935 4034 6995
rect 4086 6975 4344 6995
rect 4030 6929 4086 6935
rect 4030 6741 4060 6929
rect 4115 6920 4315 6945
rect 4396 6935 4400 6995
rect 4344 6929 4400 6935
rect 4115 6900 4185 6920
rect 4090 6860 4185 6900
rect 4245 6900 4315 6920
rect 4245 6860 4340 6900
rect 4090 6810 4340 6860
rect 4090 6770 4185 6810
rect 4115 6750 4185 6770
rect 4245 6770 4340 6810
rect 4245 6750 4315 6770
rect 4030 6735 4086 6741
rect 4030 6675 4034 6735
rect 4115 6725 4315 6750
rect 4370 6741 4400 6929
rect 4344 6735 4400 6741
rect 4086 6675 4344 6695
rect 4396 6675 4400 6735
rect 4030 6665 4400 6675
rect 4430 6995 4800 7005
rect 4430 6935 4434 6995
rect 4486 6975 4744 6995
rect 4430 6929 4486 6935
rect 4430 6741 4460 6929
rect 4515 6920 4715 6945
rect 4796 6935 4800 6995
rect 4744 6929 4800 6935
rect 4515 6900 4585 6920
rect 4490 6860 4585 6900
rect 4645 6900 4715 6920
rect 4645 6860 4740 6900
rect 4490 6810 4740 6860
rect 4490 6770 4585 6810
rect 4515 6750 4585 6770
rect 4645 6770 4740 6810
rect 4645 6750 4715 6770
rect 4430 6735 4486 6741
rect 4430 6675 4434 6735
rect 4515 6725 4715 6750
rect 4770 6741 4800 6929
rect 4744 6735 4800 6741
rect 4486 6675 4744 6695
rect 4796 6675 4800 6735
rect 4430 6665 4800 6675
rect 4830 6995 5200 7005
rect 4830 6935 4834 6995
rect 4886 6975 5144 6995
rect 4830 6929 4886 6935
rect 4830 6741 4860 6929
rect 4915 6920 5115 6945
rect 5196 6935 5200 6995
rect 5144 6929 5200 6935
rect 4915 6900 4985 6920
rect 4890 6860 4985 6900
rect 5045 6900 5115 6920
rect 5045 6860 5140 6900
rect 4890 6810 5140 6860
rect 4890 6770 4985 6810
rect 4915 6750 4985 6770
rect 5045 6770 5140 6810
rect 5045 6750 5115 6770
rect 4830 6735 4886 6741
rect 4830 6675 4834 6735
rect 4915 6725 5115 6750
rect 5170 6741 5200 6929
rect 5144 6735 5200 6741
rect 4886 6675 5144 6695
rect 5196 6675 5200 6735
rect 4830 6665 5200 6675
rect 5230 6995 5600 7005
rect 5230 6935 5234 6995
rect 5286 6975 5544 6995
rect 5230 6929 5286 6935
rect 5230 6741 5260 6929
rect 5315 6920 5515 6945
rect 5596 6935 5600 6995
rect 5544 6929 5600 6935
rect 5315 6900 5385 6920
rect 5290 6860 5385 6900
rect 5445 6900 5515 6920
rect 5445 6860 5540 6900
rect 5290 6810 5540 6860
rect 5290 6770 5385 6810
rect 5315 6750 5385 6770
rect 5445 6770 5540 6810
rect 5445 6750 5515 6770
rect 5230 6735 5286 6741
rect 5230 6675 5234 6735
rect 5315 6725 5515 6750
rect 5570 6741 5600 6929
rect 5544 6735 5600 6741
rect 5286 6675 5544 6695
rect 5596 6675 5600 6735
rect 5230 6665 5600 6675
rect 5630 6995 6000 7005
rect 5630 6935 5634 6995
rect 5686 6975 5944 6995
rect 5630 6929 5686 6935
rect 5630 6741 5660 6929
rect 5715 6920 5915 6945
rect 5996 6935 6000 6995
rect 5944 6929 6000 6935
rect 5715 6900 5785 6920
rect 5690 6860 5785 6900
rect 5845 6900 5915 6920
rect 5845 6860 5940 6900
rect 5690 6810 5940 6860
rect 5690 6770 5785 6810
rect 5715 6750 5785 6770
rect 5845 6770 5940 6810
rect 5845 6750 5915 6770
rect 5630 6735 5686 6741
rect 5630 6675 5634 6735
rect 5715 6725 5915 6750
rect 5970 6741 6000 6929
rect 5944 6735 6000 6741
rect 5686 6675 5944 6695
rect 5996 6675 6000 6735
rect 5630 6665 6000 6675
rect 6030 6995 6400 7005
rect 6030 6935 6034 6995
rect 6086 6975 6344 6995
rect 6030 6929 6086 6935
rect 6030 6741 6060 6929
rect 6115 6920 6315 6945
rect 6396 6935 6400 6995
rect 6344 6929 6400 6935
rect 6115 6900 6185 6920
rect 6090 6860 6185 6900
rect 6245 6900 6315 6920
rect 6245 6860 6340 6900
rect 6090 6810 6340 6860
rect 6090 6770 6185 6810
rect 6115 6750 6185 6770
rect 6245 6770 6340 6810
rect 6245 6750 6315 6770
rect 6030 6735 6086 6741
rect 6030 6675 6034 6735
rect 6115 6725 6315 6750
rect 6370 6741 6400 6929
rect 6344 6735 6400 6741
rect 6086 6675 6344 6695
rect 6396 6675 6400 6735
rect 6030 6665 6400 6675
rect 6430 6995 6800 7005
rect 6430 6935 6434 6995
rect 6486 6975 6744 6995
rect 6430 6929 6486 6935
rect 6430 6741 6460 6929
rect 6515 6920 6715 6945
rect 6796 6935 6800 6995
rect 6744 6929 6800 6935
rect 6515 6900 6585 6920
rect 6490 6860 6585 6900
rect 6645 6900 6715 6920
rect 6645 6860 6740 6900
rect 6490 6810 6740 6860
rect 6490 6770 6585 6810
rect 6515 6750 6585 6770
rect 6645 6770 6740 6810
rect 6645 6750 6715 6770
rect 6430 6735 6486 6741
rect 6430 6675 6434 6735
rect 6515 6725 6715 6750
rect 6770 6741 6800 6929
rect 6744 6735 6800 6741
rect 6486 6675 6744 6695
rect 6796 6675 6800 6735
rect 6430 6665 6800 6675
rect 6830 6995 7200 7005
rect 6830 6935 6834 6995
rect 6886 6975 7144 6995
rect 6830 6929 6886 6935
rect 6830 6741 6860 6929
rect 6915 6920 7115 6945
rect 7196 6935 7200 6995
rect 7144 6929 7200 6935
rect 6915 6900 6985 6920
rect 6890 6860 6985 6900
rect 7045 6900 7115 6920
rect 7045 6860 7140 6900
rect 6890 6810 7140 6860
rect 6890 6770 6985 6810
rect 6915 6750 6985 6770
rect 7045 6770 7140 6810
rect 7045 6750 7115 6770
rect 6830 6735 6886 6741
rect 6830 6675 6834 6735
rect 6915 6725 7115 6750
rect 7170 6741 7200 6929
rect 7144 6735 7200 6741
rect 6886 6675 7144 6695
rect 7196 6675 7200 6735
rect 6830 6665 7200 6675
rect 7230 6995 7600 7005
rect 7230 6935 7234 6995
rect 7286 6975 7544 6995
rect 7230 6929 7286 6935
rect 7230 6741 7260 6929
rect 7315 6920 7515 6945
rect 7596 6935 7600 6995
rect 7544 6929 7600 6935
rect 7315 6900 7385 6920
rect 7290 6860 7385 6900
rect 7445 6900 7515 6920
rect 7445 6860 7540 6900
rect 7290 6810 7540 6860
rect 7290 6770 7385 6810
rect 7315 6750 7385 6770
rect 7445 6770 7540 6810
rect 7445 6750 7515 6770
rect 7230 6735 7286 6741
rect 7230 6675 7234 6735
rect 7315 6725 7515 6750
rect 7570 6741 7600 6929
rect 7544 6735 7600 6741
rect 7286 6675 7544 6695
rect 7596 6675 7600 6735
rect 7230 6665 7600 6675
rect 7630 6995 8000 7005
rect 7630 6935 7634 6995
rect 7686 6975 7944 6995
rect 7630 6929 7686 6935
rect 7630 6741 7660 6929
rect 7715 6920 7915 6945
rect 7996 6935 8000 6995
rect 7944 6929 8000 6935
rect 7715 6900 7785 6920
rect 7690 6860 7785 6900
rect 7845 6900 7915 6920
rect 7845 6860 7940 6900
rect 7690 6810 7940 6860
rect 7690 6770 7785 6810
rect 7715 6750 7785 6770
rect 7845 6770 7940 6810
rect 7845 6750 7915 6770
rect 7630 6735 7686 6741
rect 7630 6675 7634 6735
rect 7715 6725 7915 6750
rect 7970 6741 8000 6929
rect 7944 6735 8000 6741
rect 7686 6675 7944 6695
rect 7996 6675 8000 6735
rect 7630 6665 8000 6675
rect 8030 6995 8400 7005
rect 8030 6935 8034 6995
rect 8086 6975 8344 6995
rect 8030 6929 8086 6935
rect 8030 6741 8060 6929
rect 8115 6920 8315 6945
rect 8396 6935 8400 6995
rect 8344 6929 8400 6935
rect 8115 6900 8185 6920
rect 8090 6860 8185 6900
rect 8245 6900 8315 6920
rect 8245 6860 8340 6900
rect 8090 6810 8340 6860
rect 8090 6770 8185 6810
rect 8115 6750 8185 6770
rect 8245 6770 8340 6810
rect 8245 6750 8315 6770
rect 8030 6735 8086 6741
rect 8030 6675 8034 6735
rect 8115 6725 8315 6750
rect 8370 6741 8400 6929
rect 8344 6735 8400 6741
rect 8086 6675 8344 6695
rect 8396 6675 8400 6735
rect 8030 6665 8400 6675
rect 8430 6995 8800 7005
rect 8430 6935 8434 6995
rect 8486 6975 8744 6995
rect 8430 6929 8486 6935
rect 8430 6741 8460 6929
rect 8515 6920 8715 6945
rect 8796 6935 8800 6995
rect 8744 6929 8800 6935
rect 8515 6900 8585 6920
rect 8490 6860 8585 6900
rect 8645 6900 8715 6920
rect 8645 6860 8740 6900
rect 8490 6810 8740 6860
rect 8490 6770 8585 6810
rect 8515 6750 8585 6770
rect 8645 6770 8740 6810
rect 8645 6750 8715 6770
rect 8430 6735 8486 6741
rect 8430 6675 8434 6735
rect 8515 6725 8715 6750
rect 8770 6741 8800 6929
rect 8744 6735 8800 6741
rect 8486 6675 8744 6695
rect 8796 6675 8800 6735
rect 8430 6665 8800 6675
rect 8830 6995 9200 7005
rect 8830 6935 8834 6995
rect 8886 6975 9144 6995
rect 8830 6929 8886 6935
rect 8830 6741 8860 6929
rect 8915 6920 9115 6945
rect 9196 6935 9200 6995
rect 9144 6929 9200 6935
rect 8915 6900 8985 6920
rect 8890 6860 8985 6900
rect 9045 6900 9115 6920
rect 9045 6860 9140 6900
rect 8890 6810 9140 6860
rect 8890 6770 8985 6810
rect 8915 6750 8985 6770
rect 9045 6770 9140 6810
rect 9045 6750 9115 6770
rect 8830 6735 8886 6741
rect 8830 6675 8834 6735
rect 8915 6725 9115 6750
rect 9170 6741 9200 6929
rect 9144 6735 9200 6741
rect 8886 6675 9144 6695
rect 9196 6675 9200 6735
rect 8830 6665 9200 6675
rect 9230 6995 9600 7005
rect 9230 6935 9234 6995
rect 9286 6975 9544 6995
rect 9230 6929 9286 6935
rect 9230 6741 9260 6929
rect 9315 6920 9515 6945
rect 9596 6935 9600 6995
rect 9544 6929 9600 6935
rect 9315 6900 9385 6920
rect 9290 6860 9385 6900
rect 9445 6900 9515 6920
rect 9445 6860 9540 6900
rect 9290 6810 9540 6860
rect 9290 6770 9385 6810
rect 9315 6750 9385 6770
rect 9445 6770 9540 6810
rect 9445 6750 9515 6770
rect 9230 6735 9286 6741
rect 9230 6675 9234 6735
rect 9315 6725 9515 6750
rect 9570 6741 9600 6929
rect 9544 6735 9600 6741
rect 9286 6675 9544 6695
rect 9596 6675 9600 6735
rect 9230 6665 9600 6675
rect 9630 6995 10000 7005
rect 9630 6935 9634 6995
rect 9686 6975 9944 6995
rect 9630 6929 9686 6935
rect 9630 6741 9660 6929
rect 9715 6920 9915 6945
rect 9996 6935 10000 6995
rect 9944 6929 10000 6935
rect 9715 6900 9785 6920
rect 9690 6860 9785 6900
rect 9845 6900 9915 6920
rect 9845 6860 9940 6900
rect 9690 6810 9940 6860
rect 9690 6770 9785 6810
rect 9715 6750 9785 6770
rect 9845 6770 9940 6810
rect 9845 6750 9915 6770
rect 9630 6735 9686 6741
rect 9630 6675 9634 6735
rect 9715 6725 9915 6750
rect 9970 6741 10000 6929
rect 9944 6735 10000 6741
rect 9686 6675 9944 6695
rect 9996 6675 10000 6735
rect 9630 6665 10000 6675
rect 10030 6995 10400 7005
rect 10030 6935 10034 6995
rect 10086 6975 10344 6995
rect 10030 6929 10086 6935
rect 10030 6741 10060 6929
rect 10115 6920 10315 6945
rect 10396 6935 10400 6995
rect 10344 6929 10400 6935
rect 10115 6900 10185 6920
rect 10090 6860 10185 6900
rect 10245 6900 10315 6920
rect 10245 6860 10340 6900
rect 10090 6810 10340 6860
rect 10090 6770 10185 6810
rect 10115 6750 10185 6770
rect 10245 6770 10340 6810
rect 10245 6750 10315 6770
rect 10030 6735 10086 6741
rect 10030 6675 10034 6735
rect 10115 6725 10315 6750
rect 10370 6741 10400 6929
rect 10344 6735 10400 6741
rect 10086 6675 10344 6695
rect 10396 6675 10400 6735
rect 10030 6665 10400 6675
rect 10430 6995 10800 7005
rect 10430 6935 10434 6995
rect 10486 6975 10744 6995
rect 10430 6929 10486 6935
rect 10430 6741 10460 6929
rect 10515 6920 10715 6945
rect 10796 6935 10800 6995
rect 10744 6929 10800 6935
rect 10515 6900 10585 6920
rect 10490 6860 10585 6900
rect 10645 6900 10715 6920
rect 10645 6860 10740 6900
rect 10490 6810 10740 6860
rect 10490 6770 10585 6810
rect 10515 6750 10585 6770
rect 10645 6770 10740 6810
rect 10645 6750 10715 6770
rect 10430 6735 10486 6741
rect 10430 6675 10434 6735
rect 10515 6725 10715 6750
rect 10770 6741 10800 6929
rect 10744 6735 10800 6741
rect 10486 6675 10744 6695
rect 10796 6675 10800 6735
rect 10430 6665 10800 6675
rect 10830 6995 11200 7005
rect 10830 6935 10834 6995
rect 10886 6975 11144 6995
rect 10830 6929 10886 6935
rect 10830 6741 10860 6929
rect 10915 6920 11115 6945
rect 11196 6935 11200 6995
rect 11144 6929 11200 6935
rect 10915 6900 10985 6920
rect 10890 6860 10985 6900
rect 11045 6900 11115 6920
rect 11045 6860 11140 6900
rect 10890 6810 11140 6860
rect 10890 6770 10985 6810
rect 10915 6750 10985 6770
rect 11045 6770 11140 6810
rect 11045 6750 11115 6770
rect 10830 6735 10886 6741
rect 10830 6675 10834 6735
rect 10915 6725 11115 6750
rect 11170 6741 11200 6929
rect 11144 6735 11200 6741
rect 10886 6675 11144 6695
rect 11196 6675 11200 6735
rect 10830 6665 11200 6675
rect 11230 6995 11600 7005
rect 11230 6935 11234 6995
rect 11286 6975 11544 6995
rect 11230 6929 11286 6935
rect 11230 6741 11260 6929
rect 11315 6920 11515 6945
rect 11596 6935 11600 6995
rect 11544 6929 11600 6935
rect 11315 6900 11385 6920
rect 11290 6860 11385 6900
rect 11445 6900 11515 6920
rect 11445 6860 11540 6900
rect 11290 6810 11540 6860
rect 11290 6770 11385 6810
rect 11315 6750 11385 6770
rect 11445 6770 11540 6810
rect 11445 6750 11515 6770
rect 11230 6735 11286 6741
rect 11230 6675 11234 6735
rect 11315 6725 11515 6750
rect 11570 6741 11600 6929
rect 11544 6735 11600 6741
rect 11286 6675 11544 6695
rect 11596 6675 11600 6735
rect 11230 6665 11600 6675
rect 11630 6995 12000 7005
rect 11630 6935 11634 6995
rect 11686 6975 11944 6995
rect 11630 6929 11686 6935
rect 11630 6741 11660 6929
rect 11715 6920 11915 6945
rect 11996 6935 12000 6995
rect 11944 6929 12000 6935
rect 11715 6900 11785 6920
rect 11690 6860 11785 6900
rect 11845 6900 11915 6920
rect 11845 6860 11940 6900
rect 11690 6810 11940 6860
rect 11690 6770 11785 6810
rect 11715 6750 11785 6770
rect 11845 6770 11940 6810
rect 11845 6750 11915 6770
rect 11630 6735 11686 6741
rect 11630 6675 11634 6735
rect 11715 6725 11915 6750
rect 11970 6741 12000 6929
rect 11944 6735 12000 6741
rect 11686 6675 11944 6695
rect 11996 6675 12000 6735
rect 11630 6665 12000 6675
rect 12030 6995 12400 7005
rect 12030 6935 12034 6995
rect 12086 6975 12344 6995
rect 12030 6929 12086 6935
rect 12030 6741 12060 6929
rect 12115 6920 12315 6945
rect 12396 6935 12400 6995
rect 12344 6929 12400 6935
rect 12115 6900 12185 6920
rect 12090 6860 12185 6900
rect 12245 6900 12315 6920
rect 12245 6860 12340 6900
rect 12090 6810 12340 6860
rect 12090 6770 12185 6810
rect 12115 6750 12185 6770
rect 12245 6770 12340 6810
rect 12245 6750 12315 6770
rect 12030 6735 12086 6741
rect 12030 6675 12034 6735
rect 12115 6725 12315 6750
rect 12370 6741 12400 6929
rect 12344 6735 12400 6741
rect 12086 6675 12344 6695
rect 12396 6675 12400 6735
rect 12030 6665 12400 6675
rect 12430 6995 12800 7005
rect 12430 6935 12434 6995
rect 12486 6975 12744 6995
rect 12430 6929 12486 6935
rect 12430 6741 12460 6929
rect 12515 6920 12715 6945
rect 12796 6935 12800 6995
rect 12744 6929 12800 6935
rect 12515 6900 12585 6920
rect 12490 6860 12585 6900
rect 12645 6900 12715 6920
rect 12645 6860 12740 6900
rect 12490 6810 12740 6860
rect 12490 6770 12585 6810
rect 12515 6750 12585 6770
rect 12645 6770 12740 6810
rect 12645 6750 12715 6770
rect 12430 6735 12486 6741
rect 12430 6675 12434 6735
rect 12515 6725 12715 6750
rect 12770 6741 12800 6929
rect 12744 6735 12800 6741
rect 12486 6675 12744 6695
rect 12796 6675 12800 6735
rect 12430 6665 12800 6675
rect 12830 6995 13200 7005
rect 12830 6935 12834 6995
rect 12886 6975 13144 6995
rect 12830 6929 12886 6935
rect 12830 6741 12860 6929
rect 12915 6920 13115 6945
rect 13196 6935 13200 6995
rect 13144 6929 13200 6935
rect 12915 6900 12985 6920
rect 12890 6860 12985 6900
rect 13045 6900 13115 6920
rect 13045 6860 13140 6900
rect 12890 6810 13140 6860
rect 12890 6770 12985 6810
rect 12915 6750 12985 6770
rect 13045 6770 13140 6810
rect 13045 6750 13115 6770
rect 12830 6735 12886 6741
rect 12830 6675 12834 6735
rect 12915 6725 13115 6750
rect 13170 6741 13200 6929
rect 13144 6735 13200 6741
rect 12886 6675 13144 6695
rect 13196 6675 13200 6735
rect 12830 6665 13200 6675
rect -370 6625 0 6635
rect -370 6565 -366 6625
rect -314 6605 -56 6625
rect -370 6559 -314 6565
rect -370 6371 -340 6559
rect -285 6550 -85 6575
rect -4 6565 0 6625
rect -56 6559 0 6565
rect -285 6530 -215 6550
rect -310 6490 -215 6530
rect -155 6530 -85 6550
rect -155 6490 -60 6530
rect -310 6440 -60 6490
rect -310 6400 -215 6440
rect -285 6380 -215 6400
rect -155 6400 -60 6440
rect -155 6380 -85 6400
rect -370 6365 -314 6371
rect -370 6305 -366 6365
rect -285 6355 -85 6380
rect -30 6371 0 6559
rect -56 6365 0 6371
rect -314 6305 -56 6325
rect -4 6305 0 6365
rect -370 6295 0 6305
rect 30 6625 400 6635
rect 30 6565 34 6625
rect 86 6605 344 6625
rect 30 6559 86 6565
rect 30 6371 60 6559
rect 115 6550 315 6575
rect 396 6565 400 6625
rect 344 6559 400 6565
rect 115 6530 185 6550
rect 90 6490 185 6530
rect 245 6530 315 6550
rect 245 6490 340 6530
rect 90 6440 340 6490
rect 90 6400 185 6440
rect 115 6380 185 6400
rect 245 6400 340 6440
rect 245 6380 315 6400
rect 30 6365 86 6371
rect 30 6305 34 6365
rect 115 6355 315 6380
rect 370 6371 400 6559
rect 344 6365 400 6371
rect 86 6305 344 6325
rect 396 6305 400 6365
rect 30 6295 400 6305
rect 430 6625 800 6635
rect 430 6565 434 6625
rect 486 6605 744 6625
rect 430 6559 486 6565
rect 430 6371 460 6559
rect 515 6550 715 6575
rect 796 6565 800 6625
rect 744 6559 800 6565
rect 515 6530 585 6550
rect 490 6490 585 6530
rect 645 6530 715 6550
rect 645 6490 740 6530
rect 490 6440 740 6490
rect 490 6400 585 6440
rect 515 6380 585 6400
rect 645 6400 740 6440
rect 645 6380 715 6400
rect 430 6365 486 6371
rect 430 6305 434 6365
rect 515 6355 715 6380
rect 770 6371 800 6559
rect 744 6365 800 6371
rect 486 6305 744 6325
rect 796 6305 800 6365
rect 430 6295 800 6305
rect 830 6625 1200 6635
rect 830 6565 834 6625
rect 886 6605 1144 6625
rect 830 6559 886 6565
rect 830 6371 860 6559
rect 915 6550 1115 6575
rect 1196 6565 1200 6625
rect 1144 6559 1200 6565
rect 915 6530 985 6550
rect 890 6490 985 6530
rect 1045 6530 1115 6550
rect 1045 6490 1140 6530
rect 890 6440 1140 6490
rect 890 6400 985 6440
rect 915 6380 985 6400
rect 1045 6400 1140 6440
rect 1045 6380 1115 6400
rect 830 6365 886 6371
rect 830 6305 834 6365
rect 915 6355 1115 6380
rect 1170 6371 1200 6559
rect 1144 6365 1200 6371
rect 886 6305 1144 6325
rect 1196 6305 1200 6365
rect 830 6295 1200 6305
rect 1230 6625 1600 6635
rect 1230 6565 1234 6625
rect 1286 6605 1544 6625
rect 1230 6559 1286 6565
rect 1230 6371 1260 6559
rect 1315 6550 1515 6575
rect 1596 6565 1600 6625
rect 1544 6559 1600 6565
rect 1315 6530 1385 6550
rect 1290 6490 1385 6530
rect 1445 6530 1515 6550
rect 1445 6490 1540 6530
rect 1290 6440 1540 6490
rect 1290 6400 1385 6440
rect 1315 6380 1385 6400
rect 1445 6400 1540 6440
rect 1445 6380 1515 6400
rect 1230 6365 1286 6371
rect 1230 6305 1234 6365
rect 1315 6355 1515 6380
rect 1570 6371 1600 6559
rect 1544 6365 1600 6371
rect 1286 6305 1544 6325
rect 1596 6305 1600 6365
rect 1230 6295 1600 6305
rect 1630 6625 2000 6635
rect 1630 6565 1634 6625
rect 1686 6605 1944 6625
rect 1630 6559 1686 6565
rect 1630 6371 1660 6559
rect 1715 6550 1915 6575
rect 1996 6565 2000 6625
rect 1944 6559 2000 6565
rect 1715 6530 1785 6550
rect 1690 6490 1785 6530
rect 1845 6530 1915 6550
rect 1845 6490 1940 6530
rect 1690 6440 1940 6490
rect 1690 6400 1785 6440
rect 1715 6380 1785 6400
rect 1845 6400 1940 6440
rect 1845 6380 1915 6400
rect 1630 6365 1686 6371
rect 1630 6305 1634 6365
rect 1715 6355 1915 6380
rect 1970 6371 2000 6559
rect 1944 6365 2000 6371
rect 1686 6305 1944 6325
rect 1996 6305 2000 6365
rect 1630 6295 2000 6305
rect 2030 6625 2400 6635
rect 2030 6565 2034 6625
rect 2086 6605 2344 6625
rect 2030 6559 2086 6565
rect 2030 6371 2060 6559
rect 2115 6550 2315 6575
rect 2396 6565 2400 6625
rect 2344 6559 2400 6565
rect 2115 6530 2185 6550
rect 2090 6490 2185 6530
rect 2245 6530 2315 6550
rect 2245 6490 2340 6530
rect 2090 6440 2340 6490
rect 2090 6400 2185 6440
rect 2115 6380 2185 6400
rect 2245 6400 2340 6440
rect 2245 6380 2315 6400
rect 2030 6365 2086 6371
rect 2030 6305 2034 6365
rect 2115 6355 2315 6380
rect 2370 6371 2400 6559
rect 2344 6365 2400 6371
rect 2086 6305 2344 6325
rect 2396 6305 2400 6365
rect 2030 6295 2400 6305
rect 2430 6625 2800 6635
rect 2430 6565 2434 6625
rect 2486 6605 2744 6625
rect 2430 6559 2486 6565
rect 2430 6371 2460 6559
rect 2515 6550 2715 6575
rect 2796 6565 2800 6625
rect 2744 6559 2800 6565
rect 2515 6530 2585 6550
rect 2490 6490 2585 6530
rect 2645 6530 2715 6550
rect 2645 6490 2740 6530
rect 2490 6440 2740 6490
rect 2490 6400 2585 6440
rect 2515 6380 2585 6400
rect 2645 6400 2740 6440
rect 2645 6380 2715 6400
rect 2430 6365 2486 6371
rect 2430 6305 2434 6365
rect 2515 6355 2715 6380
rect 2770 6371 2800 6559
rect 2744 6365 2800 6371
rect 2486 6305 2744 6325
rect 2796 6305 2800 6365
rect 2430 6295 2800 6305
rect 2830 6625 3200 6635
rect 2830 6565 2834 6625
rect 2886 6605 3144 6625
rect 2830 6559 2886 6565
rect 2830 6371 2860 6559
rect 2915 6550 3115 6575
rect 3196 6565 3200 6625
rect 3144 6559 3200 6565
rect 2915 6530 2985 6550
rect 2890 6490 2985 6530
rect 3045 6530 3115 6550
rect 3045 6490 3140 6530
rect 2890 6440 3140 6490
rect 2890 6400 2985 6440
rect 2915 6380 2985 6400
rect 3045 6400 3140 6440
rect 3045 6380 3115 6400
rect 2830 6365 2886 6371
rect 2830 6305 2834 6365
rect 2915 6355 3115 6380
rect 3170 6371 3200 6559
rect 3144 6365 3200 6371
rect 2886 6305 3144 6325
rect 3196 6305 3200 6365
rect 2830 6295 3200 6305
rect 3230 6625 3600 6635
rect 3230 6565 3234 6625
rect 3286 6605 3544 6625
rect 3230 6559 3286 6565
rect 3230 6371 3260 6559
rect 3315 6550 3515 6575
rect 3596 6565 3600 6625
rect 3544 6559 3600 6565
rect 3315 6530 3385 6550
rect 3290 6490 3385 6530
rect 3445 6530 3515 6550
rect 3445 6490 3540 6530
rect 3290 6440 3540 6490
rect 3290 6400 3385 6440
rect 3315 6380 3385 6400
rect 3445 6400 3540 6440
rect 3445 6380 3515 6400
rect 3230 6365 3286 6371
rect 3230 6305 3234 6365
rect 3315 6355 3515 6380
rect 3570 6371 3600 6559
rect 3544 6365 3600 6371
rect 3286 6305 3544 6325
rect 3596 6305 3600 6365
rect 3230 6295 3600 6305
rect 3630 6625 4000 6635
rect 3630 6565 3634 6625
rect 3686 6605 3944 6625
rect 3630 6559 3686 6565
rect 3630 6371 3660 6559
rect 3715 6550 3915 6575
rect 3996 6565 4000 6625
rect 3944 6559 4000 6565
rect 3715 6530 3785 6550
rect 3690 6490 3785 6530
rect 3845 6530 3915 6550
rect 3845 6490 3940 6530
rect 3690 6440 3940 6490
rect 3690 6400 3785 6440
rect 3715 6380 3785 6400
rect 3845 6400 3940 6440
rect 3845 6380 3915 6400
rect 3630 6365 3686 6371
rect 3630 6305 3634 6365
rect 3715 6355 3915 6380
rect 3970 6371 4000 6559
rect 3944 6365 4000 6371
rect 3686 6305 3944 6325
rect 3996 6305 4000 6365
rect 3630 6295 4000 6305
rect 4030 6625 4400 6635
rect 4030 6565 4034 6625
rect 4086 6605 4344 6625
rect 4030 6559 4086 6565
rect 4030 6371 4060 6559
rect 4115 6550 4315 6575
rect 4396 6565 4400 6625
rect 4344 6559 4400 6565
rect 4115 6530 4185 6550
rect 4090 6490 4185 6530
rect 4245 6530 4315 6550
rect 4245 6490 4340 6530
rect 4090 6440 4340 6490
rect 4090 6400 4185 6440
rect 4115 6380 4185 6400
rect 4245 6400 4340 6440
rect 4245 6380 4315 6400
rect 4030 6365 4086 6371
rect 4030 6305 4034 6365
rect 4115 6355 4315 6380
rect 4370 6371 4400 6559
rect 4344 6365 4400 6371
rect 4086 6305 4344 6325
rect 4396 6305 4400 6365
rect 4030 6295 4400 6305
rect 4430 6625 4800 6635
rect 4430 6565 4434 6625
rect 4486 6605 4744 6625
rect 4430 6559 4486 6565
rect 4430 6371 4460 6559
rect 4515 6550 4715 6575
rect 4796 6565 4800 6625
rect 4744 6559 4800 6565
rect 4515 6530 4585 6550
rect 4490 6490 4585 6530
rect 4645 6530 4715 6550
rect 4645 6490 4740 6530
rect 4490 6440 4740 6490
rect 4490 6400 4585 6440
rect 4515 6380 4585 6400
rect 4645 6400 4740 6440
rect 4645 6380 4715 6400
rect 4430 6365 4486 6371
rect 4430 6305 4434 6365
rect 4515 6355 4715 6380
rect 4770 6371 4800 6559
rect 4744 6365 4800 6371
rect 4486 6305 4744 6325
rect 4796 6305 4800 6365
rect 4430 6295 4800 6305
rect 4830 6625 5200 6635
rect 4830 6565 4834 6625
rect 4886 6605 5144 6625
rect 4830 6559 4886 6565
rect 4830 6371 4860 6559
rect 4915 6550 5115 6575
rect 5196 6565 5200 6625
rect 5144 6559 5200 6565
rect 4915 6530 4985 6550
rect 4890 6490 4985 6530
rect 5045 6530 5115 6550
rect 5045 6490 5140 6530
rect 4890 6440 5140 6490
rect 4890 6400 4985 6440
rect 4915 6380 4985 6400
rect 5045 6400 5140 6440
rect 5045 6380 5115 6400
rect 4830 6365 4886 6371
rect 4830 6305 4834 6365
rect 4915 6355 5115 6380
rect 5170 6371 5200 6559
rect 5144 6365 5200 6371
rect 4886 6305 5144 6325
rect 5196 6305 5200 6365
rect 4830 6295 5200 6305
rect 5230 6625 5600 6635
rect 5230 6565 5234 6625
rect 5286 6605 5544 6625
rect 5230 6559 5286 6565
rect 5230 6371 5260 6559
rect 5315 6550 5515 6575
rect 5596 6565 5600 6625
rect 5544 6559 5600 6565
rect 5315 6530 5385 6550
rect 5290 6490 5385 6530
rect 5445 6530 5515 6550
rect 5445 6490 5540 6530
rect 5290 6440 5540 6490
rect 5290 6400 5385 6440
rect 5315 6380 5385 6400
rect 5445 6400 5540 6440
rect 5445 6380 5515 6400
rect 5230 6365 5286 6371
rect 5230 6305 5234 6365
rect 5315 6355 5515 6380
rect 5570 6371 5600 6559
rect 5544 6365 5600 6371
rect 5286 6305 5544 6325
rect 5596 6305 5600 6365
rect 5230 6295 5600 6305
rect 5630 6625 6000 6635
rect 5630 6565 5634 6625
rect 5686 6605 5944 6625
rect 5630 6559 5686 6565
rect 5630 6371 5660 6559
rect 5715 6550 5915 6575
rect 5996 6565 6000 6625
rect 5944 6559 6000 6565
rect 5715 6530 5785 6550
rect 5690 6490 5785 6530
rect 5845 6530 5915 6550
rect 5845 6490 5940 6530
rect 5690 6440 5940 6490
rect 5690 6400 5785 6440
rect 5715 6380 5785 6400
rect 5845 6400 5940 6440
rect 5845 6380 5915 6400
rect 5630 6365 5686 6371
rect 5630 6305 5634 6365
rect 5715 6355 5915 6380
rect 5970 6371 6000 6559
rect 5944 6365 6000 6371
rect 5686 6305 5944 6325
rect 5996 6305 6000 6365
rect 5630 6295 6000 6305
rect 6030 6625 6400 6635
rect 6030 6565 6034 6625
rect 6086 6605 6344 6625
rect 6030 6559 6086 6565
rect 6030 6371 6060 6559
rect 6115 6550 6315 6575
rect 6396 6565 6400 6625
rect 6344 6559 6400 6565
rect 6115 6530 6185 6550
rect 6090 6490 6185 6530
rect 6245 6530 6315 6550
rect 6245 6490 6340 6530
rect 6090 6440 6340 6490
rect 6090 6400 6185 6440
rect 6115 6380 6185 6400
rect 6245 6400 6340 6440
rect 6245 6380 6315 6400
rect 6030 6365 6086 6371
rect 6030 6305 6034 6365
rect 6115 6355 6315 6380
rect 6370 6371 6400 6559
rect 6344 6365 6400 6371
rect 6086 6305 6344 6325
rect 6396 6305 6400 6365
rect 6030 6295 6400 6305
rect 6430 6625 6800 6635
rect 6430 6565 6434 6625
rect 6486 6605 6744 6625
rect 6430 6559 6486 6565
rect 6430 6371 6460 6559
rect 6515 6550 6715 6575
rect 6796 6565 6800 6625
rect 6744 6559 6800 6565
rect 6515 6530 6585 6550
rect 6490 6490 6585 6530
rect 6645 6530 6715 6550
rect 6645 6490 6740 6530
rect 6490 6440 6740 6490
rect 6490 6400 6585 6440
rect 6515 6380 6585 6400
rect 6645 6400 6740 6440
rect 6645 6380 6715 6400
rect 6430 6365 6486 6371
rect 6430 6305 6434 6365
rect 6515 6355 6715 6380
rect 6770 6371 6800 6559
rect 6744 6365 6800 6371
rect 6486 6305 6744 6325
rect 6796 6305 6800 6365
rect 6430 6295 6800 6305
rect 6830 6625 7200 6635
rect 6830 6565 6834 6625
rect 6886 6605 7144 6625
rect 6830 6559 6886 6565
rect 6830 6371 6860 6559
rect 6915 6550 7115 6575
rect 7196 6565 7200 6625
rect 7144 6559 7200 6565
rect 6915 6530 6985 6550
rect 6890 6490 6985 6530
rect 7045 6530 7115 6550
rect 7045 6490 7140 6530
rect 6890 6440 7140 6490
rect 6890 6400 6985 6440
rect 6915 6380 6985 6400
rect 7045 6400 7140 6440
rect 7045 6380 7115 6400
rect 6830 6365 6886 6371
rect 6830 6305 6834 6365
rect 6915 6355 7115 6380
rect 7170 6371 7200 6559
rect 7144 6365 7200 6371
rect 6886 6305 7144 6325
rect 7196 6305 7200 6365
rect 6830 6295 7200 6305
rect 7230 6625 7600 6635
rect 7230 6565 7234 6625
rect 7286 6605 7544 6625
rect 7230 6559 7286 6565
rect 7230 6371 7260 6559
rect 7315 6550 7515 6575
rect 7596 6565 7600 6625
rect 7544 6559 7600 6565
rect 7315 6530 7385 6550
rect 7290 6490 7385 6530
rect 7445 6530 7515 6550
rect 7445 6490 7540 6530
rect 7290 6440 7540 6490
rect 7290 6400 7385 6440
rect 7315 6380 7385 6400
rect 7445 6400 7540 6440
rect 7445 6380 7515 6400
rect 7230 6365 7286 6371
rect 7230 6305 7234 6365
rect 7315 6355 7515 6380
rect 7570 6371 7600 6559
rect 7544 6365 7600 6371
rect 7286 6305 7544 6325
rect 7596 6305 7600 6365
rect 7230 6295 7600 6305
rect 7630 6625 8000 6635
rect 7630 6565 7634 6625
rect 7686 6605 7944 6625
rect 7630 6559 7686 6565
rect 7630 6371 7660 6559
rect 7715 6550 7915 6575
rect 7996 6565 8000 6625
rect 7944 6559 8000 6565
rect 7715 6530 7785 6550
rect 7690 6490 7785 6530
rect 7845 6530 7915 6550
rect 7845 6490 7940 6530
rect 7690 6440 7940 6490
rect 7690 6400 7785 6440
rect 7715 6380 7785 6400
rect 7845 6400 7940 6440
rect 7845 6380 7915 6400
rect 7630 6365 7686 6371
rect 7630 6305 7634 6365
rect 7715 6355 7915 6380
rect 7970 6371 8000 6559
rect 7944 6365 8000 6371
rect 7686 6305 7944 6325
rect 7996 6305 8000 6365
rect 7630 6295 8000 6305
rect 8030 6625 8400 6635
rect 8030 6565 8034 6625
rect 8086 6605 8344 6625
rect 8030 6559 8086 6565
rect 8030 6371 8060 6559
rect 8115 6550 8315 6575
rect 8396 6565 8400 6625
rect 8344 6559 8400 6565
rect 8115 6530 8185 6550
rect 8090 6490 8185 6530
rect 8245 6530 8315 6550
rect 8245 6490 8340 6530
rect 8090 6440 8340 6490
rect 8090 6400 8185 6440
rect 8115 6380 8185 6400
rect 8245 6400 8340 6440
rect 8245 6380 8315 6400
rect 8030 6365 8086 6371
rect 8030 6305 8034 6365
rect 8115 6355 8315 6380
rect 8370 6371 8400 6559
rect 8344 6365 8400 6371
rect 8086 6305 8344 6325
rect 8396 6305 8400 6365
rect 8030 6295 8400 6305
rect 8430 6625 8800 6635
rect 8430 6565 8434 6625
rect 8486 6605 8744 6625
rect 8430 6559 8486 6565
rect 8430 6371 8460 6559
rect 8515 6550 8715 6575
rect 8796 6565 8800 6625
rect 8744 6559 8800 6565
rect 8515 6530 8585 6550
rect 8490 6490 8585 6530
rect 8645 6530 8715 6550
rect 8645 6490 8740 6530
rect 8490 6440 8740 6490
rect 8490 6400 8585 6440
rect 8515 6380 8585 6400
rect 8645 6400 8740 6440
rect 8645 6380 8715 6400
rect 8430 6365 8486 6371
rect 8430 6305 8434 6365
rect 8515 6355 8715 6380
rect 8770 6371 8800 6559
rect 8744 6365 8800 6371
rect 8486 6305 8744 6325
rect 8796 6305 8800 6365
rect 8430 6295 8800 6305
rect 8830 6625 9200 6635
rect 8830 6565 8834 6625
rect 8886 6605 9144 6625
rect 8830 6559 8886 6565
rect 8830 6371 8860 6559
rect 8915 6550 9115 6575
rect 9196 6565 9200 6625
rect 9144 6559 9200 6565
rect 8915 6530 8985 6550
rect 8890 6490 8985 6530
rect 9045 6530 9115 6550
rect 9045 6490 9140 6530
rect 8890 6440 9140 6490
rect 8890 6400 8985 6440
rect 8915 6380 8985 6400
rect 9045 6400 9140 6440
rect 9045 6380 9115 6400
rect 8830 6365 8886 6371
rect 8830 6305 8834 6365
rect 8915 6355 9115 6380
rect 9170 6371 9200 6559
rect 9144 6365 9200 6371
rect 8886 6305 9144 6325
rect 9196 6305 9200 6365
rect 8830 6295 9200 6305
rect 9230 6625 9600 6635
rect 9230 6565 9234 6625
rect 9286 6605 9544 6625
rect 9230 6559 9286 6565
rect 9230 6371 9260 6559
rect 9315 6550 9515 6575
rect 9596 6565 9600 6625
rect 9544 6559 9600 6565
rect 9315 6530 9385 6550
rect 9290 6490 9385 6530
rect 9445 6530 9515 6550
rect 9445 6490 9540 6530
rect 9290 6440 9540 6490
rect 9290 6400 9385 6440
rect 9315 6380 9385 6400
rect 9445 6400 9540 6440
rect 9445 6380 9515 6400
rect 9230 6365 9286 6371
rect 9230 6305 9234 6365
rect 9315 6355 9515 6380
rect 9570 6371 9600 6559
rect 9544 6365 9600 6371
rect 9286 6305 9544 6325
rect 9596 6305 9600 6365
rect 9230 6295 9600 6305
rect 9630 6625 10000 6635
rect 9630 6565 9634 6625
rect 9686 6605 9944 6625
rect 9630 6559 9686 6565
rect 9630 6371 9660 6559
rect 9715 6550 9915 6575
rect 9996 6565 10000 6625
rect 9944 6559 10000 6565
rect 9715 6530 9785 6550
rect 9690 6490 9785 6530
rect 9845 6530 9915 6550
rect 9845 6490 9940 6530
rect 9690 6440 9940 6490
rect 9690 6400 9785 6440
rect 9715 6380 9785 6400
rect 9845 6400 9940 6440
rect 9845 6380 9915 6400
rect 9630 6365 9686 6371
rect 9630 6305 9634 6365
rect 9715 6355 9915 6380
rect 9970 6371 10000 6559
rect 9944 6365 10000 6371
rect 9686 6305 9944 6325
rect 9996 6305 10000 6365
rect 9630 6295 10000 6305
rect 10030 6625 10400 6635
rect 10030 6565 10034 6625
rect 10086 6605 10344 6625
rect 10030 6559 10086 6565
rect 10030 6371 10060 6559
rect 10115 6550 10315 6575
rect 10396 6565 10400 6625
rect 10344 6559 10400 6565
rect 10115 6530 10185 6550
rect 10090 6490 10185 6530
rect 10245 6530 10315 6550
rect 10245 6490 10340 6530
rect 10090 6440 10340 6490
rect 10090 6400 10185 6440
rect 10115 6380 10185 6400
rect 10245 6400 10340 6440
rect 10245 6380 10315 6400
rect 10030 6365 10086 6371
rect 10030 6305 10034 6365
rect 10115 6355 10315 6380
rect 10370 6371 10400 6559
rect 10344 6365 10400 6371
rect 10086 6305 10344 6325
rect 10396 6305 10400 6365
rect 10030 6295 10400 6305
rect 10430 6625 10800 6635
rect 10430 6565 10434 6625
rect 10486 6605 10744 6625
rect 10430 6559 10486 6565
rect 10430 6371 10460 6559
rect 10515 6550 10715 6575
rect 10796 6565 10800 6625
rect 10744 6559 10800 6565
rect 10515 6530 10585 6550
rect 10490 6490 10585 6530
rect 10645 6530 10715 6550
rect 10645 6490 10740 6530
rect 10490 6440 10740 6490
rect 10490 6400 10585 6440
rect 10515 6380 10585 6400
rect 10645 6400 10740 6440
rect 10645 6380 10715 6400
rect 10430 6365 10486 6371
rect 10430 6305 10434 6365
rect 10515 6355 10715 6380
rect 10770 6371 10800 6559
rect 10744 6365 10800 6371
rect 10486 6305 10744 6325
rect 10796 6305 10800 6365
rect 10430 6295 10800 6305
rect 10830 6625 11200 6635
rect 10830 6565 10834 6625
rect 10886 6605 11144 6625
rect 10830 6559 10886 6565
rect 10830 6371 10860 6559
rect 10915 6550 11115 6575
rect 11196 6565 11200 6625
rect 11144 6559 11200 6565
rect 10915 6530 10985 6550
rect 10890 6490 10985 6530
rect 11045 6530 11115 6550
rect 11045 6490 11140 6530
rect 10890 6440 11140 6490
rect 10890 6400 10985 6440
rect 10915 6380 10985 6400
rect 11045 6400 11140 6440
rect 11045 6380 11115 6400
rect 10830 6365 10886 6371
rect 10830 6305 10834 6365
rect 10915 6355 11115 6380
rect 11170 6371 11200 6559
rect 11144 6365 11200 6371
rect 10886 6305 11144 6325
rect 11196 6305 11200 6365
rect 10830 6295 11200 6305
rect 11230 6625 11600 6635
rect 11230 6565 11234 6625
rect 11286 6605 11544 6625
rect 11230 6559 11286 6565
rect 11230 6371 11260 6559
rect 11315 6550 11515 6575
rect 11596 6565 11600 6625
rect 11544 6559 11600 6565
rect 11315 6530 11385 6550
rect 11290 6490 11385 6530
rect 11445 6530 11515 6550
rect 11445 6490 11540 6530
rect 11290 6440 11540 6490
rect 11290 6400 11385 6440
rect 11315 6380 11385 6400
rect 11445 6400 11540 6440
rect 11445 6380 11515 6400
rect 11230 6365 11286 6371
rect 11230 6305 11234 6365
rect 11315 6355 11515 6380
rect 11570 6371 11600 6559
rect 11544 6365 11600 6371
rect 11286 6305 11544 6325
rect 11596 6305 11600 6365
rect 11230 6295 11600 6305
rect 11630 6625 12000 6635
rect 11630 6565 11634 6625
rect 11686 6605 11944 6625
rect 11630 6559 11686 6565
rect 11630 6371 11660 6559
rect 11715 6550 11915 6575
rect 11996 6565 12000 6625
rect 11944 6559 12000 6565
rect 11715 6530 11785 6550
rect 11690 6490 11785 6530
rect 11845 6530 11915 6550
rect 11845 6490 11940 6530
rect 11690 6440 11940 6490
rect 11690 6400 11785 6440
rect 11715 6380 11785 6400
rect 11845 6400 11940 6440
rect 11845 6380 11915 6400
rect 11630 6365 11686 6371
rect 11630 6305 11634 6365
rect 11715 6355 11915 6380
rect 11970 6371 12000 6559
rect 11944 6365 12000 6371
rect 11686 6305 11944 6325
rect 11996 6305 12000 6365
rect 11630 6295 12000 6305
rect 12030 6625 12400 6635
rect 12030 6565 12034 6625
rect 12086 6605 12344 6625
rect 12030 6559 12086 6565
rect 12030 6371 12060 6559
rect 12115 6550 12315 6575
rect 12396 6565 12400 6625
rect 12344 6559 12400 6565
rect 12115 6530 12185 6550
rect 12090 6490 12185 6530
rect 12245 6530 12315 6550
rect 12245 6490 12340 6530
rect 12090 6440 12340 6490
rect 12090 6400 12185 6440
rect 12115 6380 12185 6400
rect 12245 6400 12340 6440
rect 12245 6380 12315 6400
rect 12030 6365 12086 6371
rect 12030 6305 12034 6365
rect 12115 6355 12315 6380
rect 12370 6371 12400 6559
rect 12344 6365 12400 6371
rect 12086 6305 12344 6325
rect 12396 6305 12400 6365
rect 12030 6295 12400 6305
rect 12430 6625 12800 6635
rect 12430 6565 12434 6625
rect 12486 6605 12744 6625
rect 12430 6559 12486 6565
rect 12430 6371 12460 6559
rect 12515 6550 12715 6575
rect 12796 6565 12800 6625
rect 12744 6559 12800 6565
rect 12515 6530 12585 6550
rect 12490 6490 12585 6530
rect 12645 6530 12715 6550
rect 12645 6490 12740 6530
rect 12490 6440 12740 6490
rect 12490 6400 12585 6440
rect 12515 6380 12585 6400
rect 12645 6400 12740 6440
rect 12645 6380 12715 6400
rect 12430 6365 12486 6371
rect 12430 6305 12434 6365
rect 12515 6355 12715 6380
rect 12770 6371 12800 6559
rect 12744 6365 12800 6371
rect 12486 6305 12744 6325
rect 12796 6305 12800 6365
rect 12430 6295 12800 6305
rect 12830 6625 13200 6635
rect 12830 6565 12834 6625
rect 12886 6605 13144 6625
rect 12830 6559 12886 6565
rect 12830 6371 12860 6559
rect 12915 6550 13115 6575
rect 13196 6565 13200 6625
rect 13144 6559 13200 6565
rect 12915 6530 12985 6550
rect 12890 6490 12985 6530
rect 13045 6530 13115 6550
rect 13045 6490 13140 6530
rect 12890 6440 13140 6490
rect 12890 6400 12985 6440
rect 12915 6380 12985 6400
rect 13045 6400 13140 6440
rect 13045 6380 13115 6400
rect 12830 6365 12886 6371
rect 12830 6305 12834 6365
rect 12915 6355 13115 6380
rect 13170 6371 13200 6559
rect 13144 6365 13200 6371
rect 12886 6305 13144 6325
rect 13196 6305 13200 6365
rect 12830 6295 13200 6305
rect -370 6255 0 6265
rect -370 6195 -366 6255
rect -314 6235 -56 6255
rect -370 6189 -314 6195
rect -370 6001 -340 6189
rect -285 6180 -85 6205
rect -4 6195 0 6255
rect -56 6189 0 6195
rect -285 6160 -215 6180
rect -310 6120 -215 6160
rect -155 6160 -85 6180
rect -155 6120 -60 6160
rect -310 6070 -60 6120
rect -310 6030 -215 6070
rect -285 6010 -215 6030
rect -155 6030 -60 6070
rect -155 6010 -85 6030
rect -370 5995 -314 6001
rect -370 5935 -366 5995
rect -285 5985 -85 6010
rect -30 6001 0 6189
rect -56 5995 0 6001
rect -314 5935 -56 5955
rect -4 5935 0 5995
rect -370 5925 0 5935
rect 30 6255 400 6265
rect 30 6195 34 6255
rect 86 6235 344 6255
rect 30 6189 86 6195
rect 30 6001 60 6189
rect 115 6180 315 6205
rect 396 6195 400 6255
rect 344 6189 400 6195
rect 115 6160 185 6180
rect 90 6120 185 6160
rect 245 6160 315 6180
rect 245 6120 340 6160
rect 90 6070 340 6120
rect 90 6030 185 6070
rect 115 6010 185 6030
rect 245 6030 340 6070
rect 245 6010 315 6030
rect 30 5995 86 6001
rect 30 5935 34 5995
rect 115 5985 315 6010
rect 370 6001 400 6189
rect 344 5995 400 6001
rect 86 5935 344 5955
rect 396 5935 400 5995
rect 30 5925 400 5935
rect 430 6255 800 6265
rect 430 6195 434 6255
rect 486 6235 744 6255
rect 430 6189 486 6195
rect 430 6001 460 6189
rect 515 6180 715 6205
rect 796 6195 800 6255
rect 744 6189 800 6195
rect 515 6160 585 6180
rect 490 6120 585 6160
rect 645 6160 715 6180
rect 645 6120 740 6160
rect 490 6070 740 6120
rect 490 6030 585 6070
rect 515 6010 585 6030
rect 645 6030 740 6070
rect 645 6010 715 6030
rect 430 5995 486 6001
rect 430 5935 434 5995
rect 515 5985 715 6010
rect 770 6001 800 6189
rect 744 5995 800 6001
rect 486 5935 744 5955
rect 796 5935 800 5995
rect 430 5925 800 5935
rect 830 6255 1200 6265
rect 830 6195 834 6255
rect 886 6235 1144 6255
rect 830 6189 886 6195
rect 830 6001 860 6189
rect 915 6180 1115 6205
rect 1196 6195 1200 6255
rect 1144 6189 1200 6195
rect 915 6160 985 6180
rect 890 6120 985 6160
rect 1045 6160 1115 6180
rect 1045 6120 1140 6160
rect 890 6070 1140 6120
rect 890 6030 985 6070
rect 915 6010 985 6030
rect 1045 6030 1140 6070
rect 1045 6010 1115 6030
rect 830 5995 886 6001
rect 830 5935 834 5995
rect 915 5985 1115 6010
rect 1170 6001 1200 6189
rect 1144 5995 1200 6001
rect 886 5935 1144 5955
rect 1196 5935 1200 5995
rect 830 5925 1200 5935
rect 1230 6255 1600 6265
rect 1230 6195 1234 6255
rect 1286 6235 1544 6255
rect 1230 6189 1286 6195
rect 1230 6001 1260 6189
rect 1315 6180 1515 6205
rect 1596 6195 1600 6255
rect 1544 6189 1600 6195
rect 1315 6160 1385 6180
rect 1290 6120 1385 6160
rect 1445 6160 1515 6180
rect 1445 6120 1540 6160
rect 1290 6070 1540 6120
rect 1290 6030 1385 6070
rect 1315 6010 1385 6030
rect 1445 6030 1540 6070
rect 1445 6010 1515 6030
rect 1230 5995 1286 6001
rect 1230 5935 1234 5995
rect 1315 5985 1515 6010
rect 1570 6001 1600 6189
rect 1544 5995 1600 6001
rect 1286 5935 1544 5955
rect 1596 5935 1600 5995
rect 1230 5925 1600 5935
rect 1630 6255 2000 6265
rect 1630 6195 1634 6255
rect 1686 6235 1944 6255
rect 1630 6189 1686 6195
rect 1630 6001 1660 6189
rect 1715 6180 1915 6205
rect 1996 6195 2000 6255
rect 1944 6189 2000 6195
rect 1715 6160 1785 6180
rect 1690 6120 1785 6160
rect 1845 6160 1915 6180
rect 1845 6120 1940 6160
rect 1690 6070 1940 6120
rect 1690 6030 1785 6070
rect 1715 6010 1785 6030
rect 1845 6030 1940 6070
rect 1845 6010 1915 6030
rect 1630 5995 1686 6001
rect 1630 5935 1634 5995
rect 1715 5985 1915 6010
rect 1970 6001 2000 6189
rect 1944 5995 2000 6001
rect 1686 5935 1944 5955
rect 1996 5935 2000 5995
rect 1630 5925 2000 5935
rect 2030 6255 2400 6265
rect 2030 6195 2034 6255
rect 2086 6235 2344 6255
rect 2030 6189 2086 6195
rect 2030 6001 2060 6189
rect 2115 6180 2315 6205
rect 2396 6195 2400 6255
rect 2344 6189 2400 6195
rect 2115 6160 2185 6180
rect 2090 6120 2185 6160
rect 2245 6160 2315 6180
rect 2245 6120 2340 6160
rect 2090 6070 2340 6120
rect 2090 6030 2185 6070
rect 2115 6010 2185 6030
rect 2245 6030 2340 6070
rect 2245 6010 2315 6030
rect 2030 5995 2086 6001
rect 2030 5935 2034 5995
rect 2115 5985 2315 6010
rect 2370 6001 2400 6189
rect 2344 5995 2400 6001
rect 2086 5935 2344 5955
rect 2396 5935 2400 5995
rect 2030 5925 2400 5935
rect 2430 6255 2800 6265
rect 2430 6195 2434 6255
rect 2486 6235 2744 6255
rect 2430 6189 2486 6195
rect 2430 6001 2460 6189
rect 2515 6180 2715 6205
rect 2796 6195 2800 6255
rect 2744 6189 2800 6195
rect 2515 6160 2585 6180
rect 2490 6120 2585 6160
rect 2645 6160 2715 6180
rect 2645 6120 2740 6160
rect 2490 6070 2740 6120
rect 2490 6030 2585 6070
rect 2515 6010 2585 6030
rect 2645 6030 2740 6070
rect 2645 6010 2715 6030
rect 2430 5995 2486 6001
rect 2430 5935 2434 5995
rect 2515 5985 2715 6010
rect 2770 6001 2800 6189
rect 2744 5995 2800 6001
rect 2486 5935 2744 5955
rect 2796 5935 2800 5995
rect 2430 5925 2800 5935
rect 2830 6255 3200 6265
rect 2830 6195 2834 6255
rect 2886 6235 3144 6255
rect 2830 6189 2886 6195
rect 2830 6001 2860 6189
rect 2915 6180 3115 6205
rect 3196 6195 3200 6255
rect 3144 6189 3200 6195
rect 2915 6160 2985 6180
rect 2890 6120 2985 6160
rect 3045 6160 3115 6180
rect 3045 6120 3140 6160
rect 2890 6070 3140 6120
rect 2890 6030 2985 6070
rect 2915 6010 2985 6030
rect 3045 6030 3140 6070
rect 3045 6010 3115 6030
rect 2830 5995 2886 6001
rect 2830 5935 2834 5995
rect 2915 5985 3115 6010
rect 3170 6001 3200 6189
rect 3144 5995 3200 6001
rect 2886 5935 3144 5955
rect 3196 5935 3200 5995
rect 2830 5925 3200 5935
rect 3230 6255 3600 6265
rect 3230 6195 3234 6255
rect 3286 6235 3544 6255
rect 3230 6189 3286 6195
rect 3230 6001 3260 6189
rect 3315 6180 3515 6205
rect 3596 6195 3600 6255
rect 3544 6189 3600 6195
rect 3315 6160 3385 6180
rect 3290 6120 3385 6160
rect 3445 6160 3515 6180
rect 3445 6120 3540 6160
rect 3290 6070 3540 6120
rect 3290 6030 3385 6070
rect 3315 6010 3385 6030
rect 3445 6030 3540 6070
rect 3445 6010 3515 6030
rect 3230 5995 3286 6001
rect 3230 5935 3234 5995
rect 3315 5985 3515 6010
rect 3570 6001 3600 6189
rect 3544 5995 3600 6001
rect 3286 5935 3544 5955
rect 3596 5935 3600 5995
rect 3230 5925 3600 5935
rect 3630 6255 4000 6265
rect 3630 6195 3634 6255
rect 3686 6235 3944 6255
rect 3630 6189 3686 6195
rect 3630 6001 3660 6189
rect 3715 6180 3915 6205
rect 3996 6195 4000 6255
rect 3944 6189 4000 6195
rect 3715 6160 3785 6180
rect 3690 6120 3785 6160
rect 3845 6160 3915 6180
rect 3845 6120 3940 6160
rect 3690 6070 3940 6120
rect 3690 6030 3785 6070
rect 3715 6010 3785 6030
rect 3845 6030 3940 6070
rect 3845 6010 3915 6030
rect 3630 5995 3686 6001
rect 3630 5935 3634 5995
rect 3715 5985 3915 6010
rect 3970 6001 4000 6189
rect 3944 5995 4000 6001
rect 3686 5935 3944 5955
rect 3996 5935 4000 5995
rect 3630 5925 4000 5935
rect 4030 6255 4400 6265
rect 4030 6195 4034 6255
rect 4086 6235 4344 6255
rect 4030 6189 4086 6195
rect 4030 6001 4060 6189
rect 4115 6180 4315 6205
rect 4396 6195 4400 6255
rect 4344 6189 4400 6195
rect 4115 6160 4185 6180
rect 4090 6120 4185 6160
rect 4245 6160 4315 6180
rect 4245 6120 4340 6160
rect 4090 6070 4340 6120
rect 4090 6030 4185 6070
rect 4115 6010 4185 6030
rect 4245 6030 4340 6070
rect 4245 6010 4315 6030
rect 4030 5995 4086 6001
rect 4030 5935 4034 5995
rect 4115 5985 4315 6010
rect 4370 6001 4400 6189
rect 4344 5995 4400 6001
rect 4086 5935 4344 5955
rect 4396 5935 4400 5995
rect 4030 5925 4400 5935
rect 4430 6255 4800 6265
rect 4430 6195 4434 6255
rect 4486 6235 4744 6255
rect 4430 6189 4486 6195
rect 4430 6001 4460 6189
rect 4515 6180 4715 6205
rect 4796 6195 4800 6255
rect 4744 6189 4800 6195
rect 4515 6160 4585 6180
rect 4490 6120 4585 6160
rect 4645 6160 4715 6180
rect 4645 6120 4740 6160
rect 4490 6070 4740 6120
rect 4490 6030 4585 6070
rect 4515 6010 4585 6030
rect 4645 6030 4740 6070
rect 4645 6010 4715 6030
rect 4430 5995 4486 6001
rect 4430 5935 4434 5995
rect 4515 5985 4715 6010
rect 4770 6001 4800 6189
rect 4744 5995 4800 6001
rect 4486 5935 4744 5955
rect 4796 5935 4800 5995
rect 4430 5925 4800 5935
rect 4830 6255 5200 6265
rect 4830 6195 4834 6255
rect 4886 6235 5144 6255
rect 4830 6189 4886 6195
rect 4830 6001 4860 6189
rect 4915 6180 5115 6205
rect 5196 6195 5200 6255
rect 5144 6189 5200 6195
rect 4915 6160 4985 6180
rect 4890 6120 4985 6160
rect 5045 6160 5115 6180
rect 5045 6120 5140 6160
rect 4890 6070 5140 6120
rect 4890 6030 4985 6070
rect 4915 6010 4985 6030
rect 5045 6030 5140 6070
rect 5045 6010 5115 6030
rect 4830 5995 4886 6001
rect 4830 5935 4834 5995
rect 4915 5985 5115 6010
rect 5170 6001 5200 6189
rect 5144 5995 5200 6001
rect 4886 5935 5144 5955
rect 5196 5935 5200 5995
rect 4830 5925 5200 5935
rect 5230 6255 5600 6265
rect 5230 6195 5234 6255
rect 5286 6235 5544 6255
rect 5230 6189 5286 6195
rect 5230 6001 5260 6189
rect 5315 6180 5515 6205
rect 5596 6195 5600 6255
rect 5544 6189 5600 6195
rect 5315 6160 5385 6180
rect 5290 6120 5385 6160
rect 5445 6160 5515 6180
rect 5445 6120 5540 6160
rect 5290 6070 5540 6120
rect 5290 6030 5385 6070
rect 5315 6010 5385 6030
rect 5445 6030 5540 6070
rect 5445 6010 5515 6030
rect 5230 5995 5286 6001
rect 5230 5935 5234 5995
rect 5315 5985 5515 6010
rect 5570 6001 5600 6189
rect 5544 5995 5600 6001
rect 5286 5935 5544 5955
rect 5596 5935 5600 5995
rect 5230 5925 5600 5935
rect 5630 6255 6000 6265
rect 5630 6195 5634 6255
rect 5686 6235 5944 6255
rect 5630 6189 5686 6195
rect 5630 6001 5660 6189
rect 5715 6180 5915 6205
rect 5996 6195 6000 6255
rect 5944 6189 6000 6195
rect 5715 6160 5785 6180
rect 5690 6120 5785 6160
rect 5845 6160 5915 6180
rect 5845 6120 5940 6160
rect 5690 6070 5940 6120
rect 5690 6030 5785 6070
rect 5715 6010 5785 6030
rect 5845 6030 5940 6070
rect 5845 6010 5915 6030
rect 5630 5995 5686 6001
rect 5630 5935 5634 5995
rect 5715 5985 5915 6010
rect 5970 6001 6000 6189
rect 5944 5995 6000 6001
rect 5686 5935 5944 5955
rect 5996 5935 6000 5995
rect 5630 5925 6000 5935
rect 6030 6255 6400 6265
rect 6030 6195 6034 6255
rect 6086 6235 6344 6255
rect 6030 6189 6086 6195
rect 6030 6001 6060 6189
rect 6115 6180 6315 6205
rect 6396 6195 6400 6255
rect 6344 6189 6400 6195
rect 6115 6160 6185 6180
rect 6090 6120 6185 6160
rect 6245 6160 6315 6180
rect 6245 6120 6340 6160
rect 6090 6070 6340 6120
rect 6090 6030 6185 6070
rect 6115 6010 6185 6030
rect 6245 6030 6340 6070
rect 6245 6010 6315 6030
rect 6030 5995 6086 6001
rect 6030 5935 6034 5995
rect 6115 5985 6315 6010
rect 6370 6001 6400 6189
rect 6344 5995 6400 6001
rect 6086 5935 6344 5955
rect 6396 5935 6400 5995
rect 6030 5925 6400 5935
rect 6430 6255 6800 6265
rect 6430 6195 6434 6255
rect 6486 6235 6744 6255
rect 6430 6189 6486 6195
rect 6430 6001 6460 6189
rect 6515 6180 6715 6205
rect 6796 6195 6800 6255
rect 6744 6189 6800 6195
rect 6515 6160 6585 6180
rect 6490 6120 6585 6160
rect 6645 6160 6715 6180
rect 6645 6120 6740 6160
rect 6490 6070 6740 6120
rect 6490 6030 6585 6070
rect 6515 6010 6585 6030
rect 6645 6030 6740 6070
rect 6645 6010 6715 6030
rect 6430 5995 6486 6001
rect 6430 5935 6434 5995
rect 6515 5985 6715 6010
rect 6770 6001 6800 6189
rect 6744 5995 6800 6001
rect 6486 5935 6744 5955
rect 6796 5935 6800 5995
rect 6430 5925 6800 5935
rect 6830 6255 7200 6265
rect 6830 6195 6834 6255
rect 6886 6235 7144 6255
rect 6830 6189 6886 6195
rect 6830 6001 6860 6189
rect 6915 6180 7115 6205
rect 7196 6195 7200 6255
rect 7144 6189 7200 6195
rect 6915 6160 6985 6180
rect 6890 6120 6985 6160
rect 7045 6160 7115 6180
rect 7045 6120 7140 6160
rect 6890 6070 7140 6120
rect 6890 6030 6985 6070
rect 6915 6010 6985 6030
rect 7045 6030 7140 6070
rect 7045 6010 7115 6030
rect 6830 5995 6886 6001
rect 6830 5935 6834 5995
rect 6915 5985 7115 6010
rect 7170 6001 7200 6189
rect 7144 5995 7200 6001
rect 6886 5935 7144 5955
rect 7196 5935 7200 5995
rect 6830 5925 7200 5935
rect 7230 6255 7600 6265
rect 7230 6195 7234 6255
rect 7286 6235 7544 6255
rect 7230 6189 7286 6195
rect 7230 6001 7260 6189
rect 7315 6180 7515 6205
rect 7596 6195 7600 6255
rect 7544 6189 7600 6195
rect 7315 6160 7385 6180
rect 7290 6120 7385 6160
rect 7445 6160 7515 6180
rect 7445 6120 7540 6160
rect 7290 6070 7540 6120
rect 7290 6030 7385 6070
rect 7315 6010 7385 6030
rect 7445 6030 7540 6070
rect 7445 6010 7515 6030
rect 7230 5995 7286 6001
rect 7230 5935 7234 5995
rect 7315 5985 7515 6010
rect 7570 6001 7600 6189
rect 7544 5995 7600 6001
rect 7286 5935 7544 5955
rect 7596 5935 7600 5995
rect 7230 5925 7600 5935
rect 7630 6255 8000 6265
rect 7630 6195 7634 6255
rect 7686 6235 7944 6255
rect 7630 6189 7686 6195
rect 7630 6001 7660 6189
rect 7715 6180 7915 6205
rect 7996 6195 8000 6255
rect 7944 6189 8000 6195
rect 7715 6160 7785 6180
rect 7690 6120 7785 6160
rect 7845 6160 7915 6180
rect 7845 6120 7940 6160
rect 7690 6070 7940 6120
rect 7690 6030 7785 6070
rect 7715 6010 7785 6030
rect 7845 6030 7940 6070
rect 7845 6010 7915 6030
rect 7630 5995 7686 6001
rect 7630 5935 7634 5995
rect 7715 5985 7915 6010
rect 7970 6001 8000 6189
rect 7944 5995 8000 6001
rect 7686 5935 7944 5955
rect 7996 5935 8000 5995
rect 7630 5925 8000 5935
rect 8030 6255 8400 6265
rect 8030 6195 8034 6255
rect 8086 6235 8344 6255
rect 8030 6189 8086 6195
rect 8030 6001 8060 6189
rect 8115 6180 8315 6205
rect 8396 6195 8400 6255
rect 8344 6189 8400 6195
rect 8115 6160 8185 6180
rect 8090 6120 8185 6160
rect 8245 6160 8315 6180
rect 8245 6120 8340 6160
rect 8090 6070 8340 6120
rect 8090 6030 8185 6070
rect 8115 6010 8185 6030
rect 8245 6030 8340 6070
rect 8245 6010 8315 6030
rect 8030 5995 8086 6001
rect 8030 5935 8034 5995
rect 8115 5985 8315 6010
rect 8370 6001 8400 6189
rect 8344 5995 8400 6001
rect 8086 5935 8344 5955
rect 8396 5935 8400 5995
rect 8030 5925 8400 5935
rect 8430 6255 8800 6265
rect 8430 6195 8434 6255
rect 8486 6235 8744 6255
rect 8430 6189 8486 6195
rect 8430 6001 8460 6189
rect 8515 6180 8715 6205
rect 8796 6195 8800 6255
rect 8744 6189 8800 6195
rect 8515 6160 8585 6180
rect 8490 6120 8585 6160
rect 8645 6160 8715 6180
rect 8645 6120 8740 6160
rect 8490 6070 8740 6120
rect 8490 6030 8585 6070
rect 8515 6010 8585 6030
rect 8645 6030 8740 6070
rect 8645 6010 8715 6030
rect 8430 5995 8486 6001
rect 8430 5935 8434 5995
rect 8515 5985 8715 6010
rect 8770 6001 8800 6189
rect 8744 5995 8800 6001
rect 8486 5935 8744 5955
rect 8796 5935 8800 5995
rect 8430 5925 8800 5935
rect 8830 6255 9200 6265
rect 8830 6195 8834 6255
rect 8886 6235 9144 6255
rect 8830 6189 8886 6195
rect 8830 6001 8860 6189
rect 8915 6180 9115 6205
rect 9196 6195 9200 6255
rect 9144 6189 9200 6195
rect 8915 6160 8985 6180
rect 8890 6120 8985 6160
rect 9045 6160 9115 6180
rect 9045 6120 9140 6160
rect 8890 6070 9140 6120
rect 8890 6030 8985 6070
rect 8915 6010 8985 6030
rect 9045 6030 9140 6070
rect 9045 6010 9115 6030
rect 8830 5995 8886 6001
rect 8830 5935 8834 5995
rect 8915 5985 9115 6010
rect 9170 6001 9200 6189
rect 9144 5995 9200 6001
rect 8886 5935 9144 5955
rect 9196 5935 9200 5995
rect 8830 5925 9200 5935
rect 9230 6255 9600 6265
rect 9230 6195 9234 6255
rect 9286 6235 9544 6255
rect 9230 6189 9286 6195
rect 9230 6001 9260 6189
rect 9315 6180 9515 6205
rect 9596 6195 9600 6255
rect 9544 6189 9600 6195
rect 9315 6160 9385 6180
rect 9290 6120 9385 6160
rect 9445 6160 9515 6180
rect 9445 6120 9540 6160
rect 9290 6070 9540 6120
rect 9290 6030 9385 6070
rect 9315 6010 9385 6030
rect 9445 6030 9540 6070
rect 9445 6010 9515 6030
rect 9230 5995 9286 6001
rect 9230 5935 9234 5995
rect 9315 5985 9515 6010
rect 9570 6001 9600 6189
rect 9544 5995 9600 6001
rect 9286 5935 9544 5955
rect 9596 5935 9600 5995
rect 9230 5925 9600 5935
rect 9630 6255 10000 6265
rect 9630 6195 9634 6255
rect 9686 6235 9944 6255
rect 9630 6189 9686 6195
rect 9630 6001 9660 6189
rect 9715 6180 9915 6205
rect 9996 6195 10000 6255
rect 9944 6189 10000 6195
rect 9715 6160 9785 6180
rect 9690 6120 9785 6160
rect 9845 6160 9915 6180
rect 9845 6120 9940 6160
rect 9690 6070 9940 6120
rect 9690 6030 9785 6070
rect 9715 6010 9785 6030
rect 9845 6030 9940 6070
rect 9845 6010 9915 6030
rect 9630 5995 9686 6001
rect 9630 5935 9634 5995
rect 9715 5985 9915 6010
rect 9970 6001 10000 6189
rect 9944 5995 10000 6001
rect 9686 5935 9944 5955
rect 9996 5935 10000 5995
rect 9630 5925 10000 5935
rect 10030 6255 10400 6265
rect 10030 6195 10034 6255
rect 10086 6235 10344 6255
rect 10030 6189 10086 6195
rect 10030 6001 10060 6189
rect 10115 6180 10315 6205
rect 10396 6195 10400 6255
rect 10344 6189 10400 6195
rect 10115 6160 10185 6180
rect 10090 6120 10185 6160
rect 10245 6160 10315 6180
rect 10245 6120 10340 6160
rect 10090 6070 10340 6120
rect 10090 6030 10185 6070
rect 10115 6010 10185 6030
rect 10245 6030 10340 6070
rect 10245 6010 10315 6030
rect 10030 5995 10086 6001
rect 10030 5935 10034 5995
rect 10115 5985 10315 6010
rect 10370 6001 10400 6189
rect 10344 5995 10400 6001
rect 10086 5935 10344 5955
rect 10396 5935 10400 5995
rect 10030 5925 10400 5935
rect 10430 6255 10800 6265
rect 10430 6195 10434 6255
rect 10486 6235 10744 6255
rect 10430 6189 10486 6195
rect 10430 6001 10460 6189
rect 10515 6180 10715 6205
rect 10796 6195 10800 6255
rect 10744 6189 10800 6195
rect 10515 6160 10585 6180
rect 10490 6120 10585 6160
rect 10645 6160 10715 6180
rect 10645 6120 10740 6160
rect 10490 6070 10740 6120
rect 10490 6030 10585 6070
rect 10515 6010 10585 6030
rect 10645 6030 10740 6070
rect 10645 6010 10715 6030
rect 10430 5995 10486 6001
rect 10430 5935 10434 5995
rect 10515 5985 10715 6010
rect 10770 6001 10800 6189
rect 10744 5995 10800 6001
rect 10486 5935 10744 5955
rect 10796 5935 10800 5995
rect 10430 5925 10800 5935
rect 10830 6255 11200 6265
rect 10830 6195 10834 6255
rect 10886 6235 11144 6255
rect 10830 6189 10886 6195
rect 10830 6001 10860 6189
rect 10915 6180 11115 6205
rect 11196 6195 11200 6255
rect 11144 6189 11200 6195
rect 10915 6160 10985 6180
rect 10890 6120 10985 6160
rect 11045 6160 11115 6180
rect 11045 6120 11140 6160
rect 10890 6070 11140 6120
rect 10890 6030 10985 6070
rect 10915 6010 10985 6030
rect 11045 6030 11140 6070
rect 11045 6010 11115 6030
rect 10830 5995 10886 6001
rect 10830 5935 10834 5995
rect 10915 5985 11115 6010
rect 11170 6001 11200 6189
rect 11144 5995 11200 6001
rect 10886 5935 11144 5955
rect 11196 5935 11200 5995
rect 10830 5925 11200 5935
rect 11230 6255 11600 6265
rect 11230 6195 11234 6255
rect 11286 6235 11544 6255
rect 11230 6189 11286 6195
rect 11230 6001 11260 6189
rect 11315 6180 11515 6205
rect 11596 6195 11600 6255
rect 11544 6189 11600 6195
rect 11315 6160 11385 6180
rect 11290 6120 11385 6160
rect 11445 6160 11515 6180
rect 11445 6120 11540 6160
rect 11290 6070 11540 6120
rect 11290 6030 11385 6070
rect 11315 6010 11385 6030
rect 11445 6030 11540 6070
rect 11445 6010 11515 6030
rect 11230 5995 11286 6001
rect 11230 5935 11234 5995
rect 11315 5985 11515 6010
rect 11570 6001 11600 6189
rect 11544 5995 11600 6001
rect 11286 5935 11544 5955
rect 11596 5935 11600 5995
rect 11230 5925 11600 5935
rect 11630 6255 12000 6265
rect 11630 6195 11634 6255
rect 11686 6235 11944 6255
rect 11630 6189 11686 6195
rect 11630 6001 11660 6189
rect 11715 6180 11915 6205
rect 11996 6195 12000 6255
rect 11944 6189 12000 6195
rect 11715 6160 11785 6180
rect 11690 6120 11785 6160
rect 11845 6160 11915 6180
rect 11845 6120 11940 6160
rect 11690 6070 11940 6120
rect 11690 6030 11785 6070
rect 11715 6010 11785 6030
rect 11845 6030 11940 6070
rect 11845 6010 11915 6030
rect 11630 5995 11686 6001
rect 11630 5935 11634 5995
rect 11715 5985 11915 6010
rect 11970 6001 12000 6189
rect 11944 5995 12000 6001
rect 11686 5935 11944 5955
rect 11996 5935 12000 5995
rect 11630 5925 12000 5935
rect 12030 6255 12400 6265
rect 12030 6195 12034 6255
rect 12086 6235 12344 6255
rect 12030 6189 12086 6195
rect 12030 6001 12060 6189
rect 12115 6180 12315 6205
rect 12396 6195 12400 6255
rect 12344 6189 12400 6195
rect 12115 6160 12185 6180
rect 12090 6120 12185 6160
rect 12245 6160 12315 6180
rect 12245 6120 12340 6160
rect 12090 6070 12340 6120
rect 12090 6030 12185 6070
rect 12115 6010 12185 6030
rect 12245 6030 12340 6070
rect 12245 6010 12315 6030
rect 12030 5995 12086 6001
rect 12030 5935 12034 5995
rect 12115 5985 12315 6010
rect 12370 6001 12400 6189
rect 12344 5995 12400 6001
rect 12086 5935 12344 5955
rect 12396 5935 12400 5995
rect 12030 5925 12400 5935
rect 12430 6255 12800 6265
rect 12430 6195 12434 6255
rect 12486 6235 12744 6255
rect 12430 6189 12486 6195
rect 12430 6001 12460 6189
rect 12515 6180 12715 6205
rect 12796 6195 12800 6255
rect 12744 6189 12800 6195
rect 12515 6160 12585 6180
rect 12490 6120 12585 6160
rect 12645 6160 12715 6180
rect 12645 6120 12740 6160
rect 12490 6070 12740 6120
rect 12490 6030 12585 6070
rect 12515 6010 12585 6030
rect 12645 6030 12740 6070
rect 12645 6010 12715 6030
rect 12430 5995 12486 6001
rect 12430 5935 12434 5995
rect 12515 5985 12715 6010
rect 12770 6001 12800 6189
rect 12744 5995 12800 6001
rect 12486 5935 12744 5955
rect 12796 5935 12800 5995
rect 12430 5925 12800 5935
rect 12830 6255 13200 6265
rect 12830 6195 12834 6255
rect 12886 6235 13144 6255
rect 12830 6189 12886 6195
rect 12830 6001 12860 6189
rect 12915 6180 13115 6205
rect 13196 6195 13200 6255
rect 13144 6189 13200 6195
rect 12915 6160 12985 6180
rect 12890 6120 12985 6160
rect 13045 6160 13115 6180
rect 13045 6120 13140 6160
rect 12890 6070 13140 6120
rect 12890 6030 12985 6070
rect 12915 6010 12985 6030
rect 13045 6030 13140 6070
rect 13045 6010 13115 6030
rect 12830 5995 12886 6001
rect 12830 5935 12834 5995
rect 12915 5985 13115 6010
rect 13170 6001 13200 6189
rect 13144 5995 13200 6001
rect 12886 5935 13144 5955
rect 13196 5935 13200 5995
rect 12830 5925 13200 5935
rect -370 5885 0 5895
rect -370 5825 -366 5885
rect -314 5865 -56 5885
rect -370 5819 -314 5825
rect -370 5631 -340 5819
rect -285 5810 -85 5835
rect -4 5825 0 5885
rect -56 5819 0 5825
rect -285 5790 -215 5810
rect -310 5750 -215 5790
rect -155 5790 -85 5810
rect -155 5750 -60 5790
rect -310 5700 -60 5750
rect -310 5660 -215 5700
rect -285 5640 -215 5660
rect -155 5660 -60 5700
rect -155 5640 -85 5660
rect -370 5625 -314 5631
rect -370 5565 -366 5625
rect -285 5615 -85 5640
rect -30 5631 0 5819
rect -56 5625 0 5631
rect -314 5565 -56 5585
rect -4 5565 0 5625
rect -370 5555 0 5565
rect 30 5885 400 5895
rect 30 5825 34 5885
rect 86 5865 344 5885
rect 30 5819 86 5825
rect 30 5631 60 5819
rect 115 5810 315 5835
rect 396 5825 400 5885
rect 344 5819 400 5825
rect 115 5790 185 5810
rect 90 5750 185 5790
rect 245 5790 315 5810
rect 245 5750 340 5790
rect 90 5700 340 5750
rect 90 5660 185 5700
rect 115 5640 185 5660
rect 245 5660 340 5700
rect 245 5640 315 5660
rect 30 5625 86 5631
rect 30 5565 34 5625
rect 115 5615 315 5640
rect 370 5631 400 5819
rect 344 5625 400 5631
rect 86 5565 344 5585
rect 396 5565 400 5625
rect 30 5555 400 5565
rect 430 5885 800 5895
rect 430 5825 434 5885
rect 486 5865 744 5885
rect 430 5819 486 5825
rect 430 5631 460 5819
rect 515 5810 715 5835
rect 796 5825 800 5885
rect 744 5819 800 5825
rect 515 5790 585 5810
rect 490 5750 585 5790
rect 645 5790 715 5810
rect 645 5750 740 5790
rect 490 5700 740 5750
rect 490 5660 585 5700
rect 515 5640 585 5660
rect 645 5660 740 5700
rect 645 5640 715 5660
rect 430 5625 486 5631
rect 430 5565 434 5625
rect 515 5615 715 5640
rect 770 5631 800 5819
rect 744 5625 800 5631
rect 486 5565 744 5585
rect 796 5565 800 5625
rect 430 5555 800 5565
rect 830 5885 1200 5895
rect 830 5825 834 5885
rect 886 5865 1144 5885
rect 830 5819 886 5825
rect 830 5631 860 5819
rect 915 5810 1115 5835
rect 1196 5825 1200 5885
rect 1144 5819 1200 5825
rect 915 5790 985 5810
rect 890 5750 985 5790
rect 1045 5790 1115 5810
rect 1045 5750 1140 5790
rect 890 5700 1140 5750
rect 890 5660 985 5700
rect 915 5640 985 5660
rect 1045 5660 1140 5700
rect 1045 5640 1115 5660
rect 830 5625 886 5631
rect 830 5565 834 5625
rect 915 5615 1115 5640
rect 1170 5631 1200 5819
rect 1144 5625 1200 5631
rect 886 5565 1144 5585
rect 1196 5565 1200 5625
rect 830 5555 1200 5565
rect 1230 5885 1600 5895
rect 1230 5825 1234 5885
rect 1286 5865 1544 5885
rect 1230 5819 1286 5825
rect 1230 5631 1260 5819
rect 1315 5810 1515 5835
rect 1596 5825 1600 5885
rect 1544 5819 1600 5825
rect 1315 5790 1385 5810
rect 1290 5750 1385 5790
rect 1445 5790 1515 5810
rect 1445 5750 1540 5790
rect 1290 5700 1540 5750
rect 1290 5660 1385 5700
rect 1315 5640 1385 5660
rect 1445 5660 1540 5700
rect 1445 5640 1515 5660
rect 1230 5625 1286 5631
rect 1230 5565 1234 5625
rect 1315 5615 1515 5640
rect 1570 5631 1600 5819
rect 1544 5625 1600 5631
rect 1286 5565 1544 5585
rect 1596 5565 1600 5625
rect 1230 5555 1600 5565
rect 1630 5885 2000 5895
rect 1630 5825 1634 5885
rect 1686 5865 1944 5885
rect 1630 5819 1686 5825
rect 1630 5631 1660 5819
rect 1715 5810 1915 5835
rect 1996 5825 2000 5885
rect 1944 5819 2000 5825
rect 1715 5790 1785 5810
rect 1690 5750 1785 5790
rect 1845 5790 1915 5810
rect 1845 5750 1940 5790
rect 1690 5700 1940 5750
rect 1690 5660 1785 5700
rect 1715 5640 1785 5660
rect 1845 5660 1940 5700
rect 1845 5640 1915 5660
rect 1630 5625 1686 5631
rect 1630 5565 1634 5625
rect 1715 5615 1915 5640
rect 1970 5631 2000 5819
rect 1944 5625 2000 5631
rect 1686 5565 1944 5585
rect 1996 5565 2000 5625
rect 1630 5555 2000 5565
rect 2030 5885 2400 5895
rect 2030 5825 2034 5885
rect 2086 5865 2344 5885
rect 2030 5819 2086 5825
rect 2030 5631 2060 5819
rect 2115 5810 2315 5835
rect 2396 5825 2400 5885
rect 2344 5819 2400 5825
rect 2115 5790 2185 5810
rect 2090 5750 2185 5790
rect 2245 5790 2315 5810
rect 2245 5750 2340 5790
rect 2090 5700 2340 5750
rect 2090 5660 2185 5700
rect 2115 5640 2185 5660
rect 2245 5660 2340 5700
rect 2245 5640 2315 5660
rect 2030 5625 2086 5631
rect 2030 5565 2034 5625
rect 2115 5615 2315 5640
rect 2370 5631 2400 5819
rect 2344 5625 2400 5631
rect 2086 5565 2344 5585
rect 2396 5565 2400 5625
rect 2030 5555 2400 5565
rect 2430 5885 2800 5895
rect 2430 5825 2434 5885
rect 2486 5865 2744 5885
rect 2430 5819 2486 5825
rect 2430 5631 2460 5819
rect 2515 5810 2715 5835
rect 2796 5825 2800 5885
rect 2744 5819 2800 5825
rect 2515 5790 2585 5810
rect 2490 5750 2585 5790
rect 2645 5790 2715 5810
rect 2645 5750 2740 5790
rect 2490 5700 2740 5750
rect 2490 5660 2585 5700
rect 2515 5640 2585 5660
rect 2645 5660 2740 5700
rect 2645 5640 2715 5660
rect 2430 5625 2486 5631
rect 2430 5565 2434 5625
rect 2515 5615 2715 5640
rect 2770 5631 2800 5819
rect 2744 5625 2800 5631
rect 2486 5565 2744 5585
rect 2796 5565 2800 5625
rect 2430 5555 2800 5565
rect 2830 5885 3200 5895
rect 2830 5825 2834 5885
rect 2886 5865 3144 5885
rect 2830 5819 2886 5825
rect 2830 5631 2860 5819
rect 2915 5810 3115 5835
rect 3196 5825 3200 5885
rect 3144 5819 3200 5825
rect 2915 5790 2985 5810
rect 2890 5750 2985 5790
rect 3045 5790 3115 5810
rect 3045 5750 3140 5790
rect 2890 5700 3140 5750
rect 2890 5660 2985 5700
rect 2915 5640 2985 5660
rect 3045 5660 3140 5700
rect 3045 5640 3115 5660
rect 2830 5625 2886 5631
rect 2830 5565 2834 5625
rect 2915 5615 3115 5640
rect 3170 5631 3200 5819
rect 3144 5625 3200 5631
rect 2886 5565 3144 5585
rect 3196 5565 3200 5625
rect 2830 5555 3200 5565
rect 3230 5885 3600 5895
rect 3230 5825 3234 5885
rect 3286 5865 3544 5885
rect 3230 5819 3286 5825
rect 3230 5631 3260 5819
rect 3315 5810 3515 5835
rect 3596 5825 3600 5885
rect 3544 5819 3600 5825
rect 3315 5790 3385 5810
rect 3290 5750 3385 5790
rect 3445 5790 3515 5810
rect 3445 5750 3540 5790
rect 3290 5700 3540 5750
rect 3290 5660 3385 5700
rect 3315 5640 3385 5660
rect 3445 5660 3540 5700
rect 3445 5640 3515 5660
rect 3230 5625 3286 5631
rect 3230 5565 3234 5625
rect 3315 5615 3515 5640
rect 3570 5631 3600 5819
rect 3544 5625 3600 5631
rect 3286 5565 3544 5585
rect 3596 5565 3600 5625
rect 3230 5555 3600 5565
rect 3630 5885 4000 5895
rect 3630 5825 3634 5885
rect 3686 5865 3944 5885
rect 3630 5819 3686 5825
rect 3630 5631 3660 5819
rect 3715 5810 3915 5835
rect 3996 5825 4000 5885
rect 3944 5819 4000 5825
rect 3715 5790 3785 5810
rect 3690 5750 3785 5790
rect 3845 5790 3915 5810
rect 3845 5750 3940 5790
rect 3690 5700 3940 5750
rect 3690 5660 3785 5700
rect 3715 5640 3785 5660
rect 3845 5660 3940 5700
rect 3845 5640 3915 5660
rect 3630 5625 3686 5631
rect 3630 5565 3634 5625
rect 3715 5615 3915 5640
rect 3970 5631 4000 5819
rect 3944 5625 4000 5631
rect 3686 5565 3944 5585
rect 3996 5565 4000 5625
rect 3630 5555 4000 5565
rect 4030 5885 4400 5895
rect 4030 5825 4034 5885
rect 4086 5865 4344 5885
rect 4030 5819 4086 5825
rect 4030 5631 4060 5819
rect 4115 5810 4315 5835
rect 4396 5825 4400 5885
rect 4344 5819 4400 5825
rect 4115 5790 4185 5810
rect 4090 5750 4185 5790
rect 4245 5790 4315 5810
rect 4245 5750 4340 5790
rect 4090 5700 4340 5750
rect 4090 5660 4185 5700
rect 4115 5640 4185 5660
rect 4245 5660 4340 5700
rect 4245 5640 4315 5660
rect 4030 5625 4086 5631
rect 4030 5565 4034 5625
rect 4115 5615 4315 5640
rect 4370 5631 4400 5819
rect 4344 5625 4400 5631
rect 4086 5565 4344 5585
rect 4396 5565 4400 5625
rect 4030 5555 4400 5565
rect 4430 5885 4800 5895
rect 4430 5825 4434 5885
rect 4486 5865 4744 5885
rect 4430 5819 4486 5825
rect 4430 5631 4460 5819
rect 4515 5810 4715 5835
rect 4796 5825 4800 5885
rect 4744 5819 4800 5825
rect 4515 5790 4585 5810
rect 4490 5750 4585 5790
rect 4645 5790 4715 5810
rect 4645 5750 4740 5790
rect 4490 5700 4740 5750
rect 4490 5660 4585 5700
rect 4515 5640 4585 5660
rect 4645 5660 4740 5700
rect 4645 5640 4715 5660
rect 4430 5625 4486 5631
rect 4430 5565 4434 5625
rect 4515 5615 4715 5640
rect 4770 5631 4800 5819
rect 4744 5625 4800 5631
rect 4486 5565 4744 5585
rect 4796 5565 4800 5625
rect 4430 5555 4800 5565
rect 4830 5885 5200 5895
rect 4830 5825 4834 5885
rect 4886 5865 5144 5885
rect 4830 5819 4886 5825
rect 4830 5631 4860 5819
rect 4915 5810 5115 5835
rect 5196 5825 5200 5885
rect 5144 5819 5200 5825
rect 4915 5790 4985 5810
rect 4890 5750 4985 5790
rect 5045 5790 5115 5810
rect 5045 5750 5140 5790
rect 4890 5700 5140 5750
rect 4890 5660 4985 5700
rect 4915 5640 4985 5660
rect 5045 5660 5140 5700
rect 5045 5640 5115 5660
rect 4830 5625 4886 5631
rect 4830 5565 4834 5625
rect 4915 5615 5115 5640
rect 5170 5631 5200 5819
rect 5144 5625 5200 5631
rect 4886 5565 5144 5585
rect 5196 5565 5200 5625
rect 4830 5555 5200 5565
rect 5230 5885 5600 5895
rect 5230 5825 5234 5885
rect 5286 5865 5544 5885
rect 5230 5819 5286 5825
rect 5230 5631 5260 5819
rect 5315 5810 5515 5835
rect 5596 5825 5600 5885
rect 5544 5819 5600 5825
rect 5315 5790 5385 5810
rect 5290 5750 5385 5790
rect 5445 5790 5515 5810
rect 5445 5750 5540 5790
rect 5290 5700 5540 5750
rect 5290 5660 5385 5700
rect 5315 5640 5385 5660
rect 5445 5660 5540 5700
rect 5445 5640 5515 5660
rect 5230 5625 5286 5631
rect 5230 5565 5234 5625
rect 5315 5615 5515 5640
rect 5570 5631 5600 5819
rect 5544 5625 5600 5631
rect 5286 5565 5544 5585
rect 5596 5565 5600 5625
rect 5230 5555 5600 5565
rect 5630 5885 6000 5895
rect 5630 5825 5634 5885
rect 5686 5865 5944 5885
rect 5630 5819 5686 5825
rect 5630 5631 5660 5819
rect 5715 5810 5915 5835
rect 5996 5825 6000 5885
rect 5944 5819 6000 5825
rect 5715 5790 5785 5810
rect 5690 5750 5785 5790
rect 5845 5790 5915 5810
rect 5845 5750 5940 5790
rect 5690 5700 5940 5750
rect 5690 5660 5785 5700
rect 5715 5640 5785 5660
rect 5845 5660 5940 5700
rect 5845 5640 5915 5660
rect 5630 5625 5686 5631
rect 5630 5565 5634 5625
rect 5715 5615 5915 5640
rect 5970 5631 6000 5819
rect 5944 5625 6000 5631
rect 5686 5565 5944 5585
rect 5996 5565 6000 5625
rect 5630 5555 6000 5565
rect 6030 5885 6400 5895
rect 6030 5825 6034 5885
rect 6086 5865 6344 5885
rect 6030 5819 6086 5825
rect 6030 5631 6060 5819
rect 6115 5810 6315 5835
rect 6396 5825 6400 5885
rect 6344 5819 6400 5825
rect 6115 5790 6185 5810
rect 6090 5750 6185 5790
rect 6245 5790 6315 5810
rect 6245 5750 6340 5790
rect 6090 5700 6340 5750
rect 6090 5660 6185 5700
rect 6115 5640 6185 5660
rect 6245 5660 6340 5700
rect 6245 5640 6315 5660
rect 6030 5625 6086 5631
rect 6030 5565 6034 5625
rect 6115 5615 6315 5640
rect 6370 5631 6400 5819
rect 6344 5625 6400 5631
rect 6086 5565 6344 5585
rect 6396 5565 6400 5625
rect 6030 5555 6400 5565
rect 6430 5885 6800 5895
rect 6430 5825 6434 5885
rect 6486 5865 6744 5885
rect 6430 5819 6486 5825
rect 6430 5631 6460 5819
rect 6515 5810 6715 5835
rect 6796 5825 6800 5885
rect 6744 5819 6800 5825
rect 6515 5790 6585 5810
rect 6490 5750 6585 5790
rect 6645 5790 6715 5810
rect 6645 5750 6740 5790
rect 6490 5700 6740 5750
rect 6490 5660 6585 5700
rect 6515 5640 6585 5660
rect 6645 5660 6740 5700
rect 6645 5640 6715 5660
rect 6430 5625 6486 5631
rect 6430 5565 6434 5625
rect 6515 5615 6715 5640
rect 6770 5631 6800 5819
rect 6744 5625 6800 5631
rect 6486 5565 6744 5585
rect 6796 5565 6800 5625
rect 6430 5555 6800 5565
rect 6830 5885 7200 5895
rect 6830 5825 6834 5885
rect 6886 5865 7144 5885
rect 6830 5819 6886 5825
rect 6830 5631 6860 5819
rect 6915 5810 7115 5835
rect 7196 5825 7200 5885
rect 7144 5819 7200 5825
rect 6915 5790 6985 5810
rect 6890 5750 6985 5790
rect 7045 5790 7115 5810
rect 7045 5750 7140 5790
rect 6890 5700 7140 5750
rect 6890 5660 6985 5700
rect 6915 5640 6985 5660
rect 7045 5660 7140 5700
rect 7045 5640 7115 5660
rect 6830 5625 6886 5631
rect 6830 5565 6834 5625
rect 6915 5615 7115 5640
rect 7170 5631 7200 5819
rect 7144 5625 7200 5631
rect 6886 5565 7144 5585
rect 7196 5565 7200 5625
rect 6830 5555 7200 5565
rect 7230 5885 7600 5895
rect 7230 5825 7234 5885
rect 7286 5865 7544 5885
rect 7230 5819 7286 5825
rect 7230 5631 7260 5819
rect 7315 5810 7515 5835
rect 7596 5825 7600 5885
rect 7544 5819 7600 5825
rect 7315 5790 7385 5810
rect 7290 5750 7385 5790
rect 7445 5790 7515 5810
rect 7445 5750 7540 5790
rect 7290 5700 7540 5750
rect 7290 5660 7385 5700
rect 7315 5640 7385 5660
rect 7445 5660 7540 5700
rect 7445 5640 7515 5660
rect 7230 5625 7286 5631
rect 7230 5565 7234 5625
rect 7315 5615 7515 5640
rect 7570 5631 7600 5819
rect 7544 5625 7600 5631
rect 7286 5565 7544 5585
rect 7596 5565 7600 5625
rect 7230 5555 7600 5565
rect 7630 5885 8000 5895
rect 7630 5825 7634 5885
rect 7686 5865 7944 5885
rect 7630 5819 7686 5825
rect 7630 5631 7660 5819
rect 7715 5810 7915 5835
rect 7996 5825 8000 5885
rect 7944 5819 8000 5825
rect 7715 5790 7785 5810
rect 7690 5750 7785 5790
rect 7845 5790 7915 5810
rect 7845 5750 7940 5790
rect 7690 5700 7940 5750
rect 7690 5660 7785 5700
rect 7715 5640 7785 5660
rect 7845 5660 7940 5700
rect 7845 5640 7915 5660
rect 7630 5625 7686 5631
rect 7630 5565 7634 5625
rect 7715 5615 7915 5640
rect 7970 5631 8000 5819
rect 7944 5625 8000 5631
rect 7686 5565 7944 5585
rect 7996 5565 8000 5625
rect 7630 5555 8000 5565
rect 8030 5885 8400 5895
rect 8030 5825 8034 5885
rect 8086 5865 8344 5885
rect 8030 5819 8086 5825
rect 8030 5631 8060 5819
rect 8115 5810 8315 5835
rect 8396 5825 8400 5885
rect 8344 5819 8400 5825
rect 8115 5790 8185 5810
rect 8090 5750 8185 5790
rect 8245 5790 8315 5810
rect 8245 5750 8340 5790
rect 8090 5700 8340 5750
rect 8090 5660 8185 5700
rect 8115 5640 8185 5660
rect 8245 5660 8340 5700
rect 8245 5640 8315 5660
rect 8030 5625 8086 5631
rect 8030 5565 8034 5625
rect 8115 5615 8315 5640
rect 8370 5631 8400 5819
rect 8344 5625 8400 5631
rect 8086 5565 8344 5585
rect 8396 5565 8400 5625
rect 8030 5555 8400 5565
rect 8430 5885 8800 5895
rect 8430 5825 8434 5885
rect 8486 5865 8744 5885
rect 8430 5819 8486 5825
rect 8430 5631 8460 5819
rect 8515 5810 8715 5835
rect 8796 5825 8800 5885
rect 8744 5819 8800 5825
rect 8515 5790 8585 5810
rect 8490 5750 8585 5790
rect 8645 5790 8715 5810
rect 8645 5750 8740 5790
rect 8490 5700 8740 5750
rect 8490 5660 8585 5700
rect 8515 5640 8585 5660
rect 8645 5660 8740 5700
rect 8645 5640 8715 5660
rect 8430 5625 8486 5631
rect 8430 5565 8434 5625
rect 8515 5615 8715 5640
rect 8770 5631 8800 5819
rect 8744 5625 8800 5631
rect 8486 5565 8744 5585
rect 8796 5565 8800 5625
rect 8430 5555 8800 5565
rect 8830 5885 9200 5895
rect 8830 5825 8834 5885
rect 8886 5865 9144 5885
rect 8830 5819 8886 5825
rect 8830 5631 8860 5819
rect 8915 5810 9115 5835
rect 9196 5825 9200 5885
rect 9144 5819 9200 5825
rect 8915 5790 8985 5810
rect 8890 5750 8985 5790
rect 9045 5790 9115 5810
rect 9045 5750 9140 5790
rect 8890 5700 9140 5750
rect 8890 5660 8985 5700
rect 8915 5640 8985 5660
rect 9045 5660 9140 5700
rect 9045 5640 9115 5660
rect 8830 5625 8886 5631
rect 8830 5565 8834 5625
rect 8915 5615 9115 5640
rect 9170 5631 9200 5819
rect 9144 5625 9200 5631
rect 8886 5565 9144 5585
rect 9196 5565 9200 5625
rect 8830 5555 9200 5565
rect 9230 5885 9600 5895
rect 9230 5825 9234 5885
rect 9286 5865 9544 5885
rect 9230 5819 9286 5825
rect 9230 5631 9260 5819
rect 9315 5810 9515 5835
rect 9596 5825 9600 5885
rect 9544 5819 9600 5825
rect 9315 5790 9385 5810
rect 9290 5750 9385 5790
rect 9445 5790 9515 5810
rect 9445 5750 9540 5790
rect 9290 5700 9540 5750
rect 9290 5660 9385 5700
rect 9315 5640 9385 5660
rect 9445 5660 9540 5700
rect 9445 5640 9515 5660
rect 9230 5625 9286 5631
rect 9230 5565 9234 5625
rect 9315 5615 9515 5640
rect 9570 5631 9600 5819
rect 9544 5625 9600 5631
rect 9286 5565 9544 5585
rect 9596 5565 9600 5625
rect 9230 5555 9600 5565
rect 9630 5885 10000 5895
rect 9630 5825 9634 5885
rect 9686 5865 9944 5885
rect 9630 5819 9686 5825
rect 9630 5631 9660 5819
rect 9715 5810 9915 5835
rect 9996 5825 10000 5885
rect 9944 5819 10000 5825
rect 9715 5790 9785 5810
rect 9690 5750 9785 5790
rect 9845 5790 9915 5810
rect 9845 5750 9940 5790
rect 9690 5700 9940 5750
rect 9690 5660 9785 5700
rect 9715 5640 9785 5660
rect 9845 5660 9940 5700
rect 9845 5640 9915 5660
rect 9630 5625 9686 5631
rect 9630 5565 9634 5625
rect 9715 5615 9915 5640
rect 9970 5631 10000 5819
rect 9944 5625 10000 5631
rect 9686 5565 9944 5585
rect 9996 5565 10000 5625
rect 9630 5555 10000 5565
rect 10030 5885 10400 5895
rect 10030 5825 10034 5885
rect 10086 5865 10344 5885
rect 10030 5819 10086 5825
rect 10030 5631 10060 5819
rect 10115 5810 10315 5835
rect 10396 5825 10400 5885
rect 10344 5819 10400 5825
rect 10115 5790 10185 5810
rect 10090 5750 10185 5790
rect 10245 5790 10315 5810
rect 10245 5750 10340 5790
rect 10090 5700 10340 5750
rect 10090 5660 10185 5700
rect 10115 5640 10185 5660
rect 10245 5660 10340 5700
rect 10245 5640 10315 5660
rect 10030 5625 10086 5631
rect 10030 5565 10034 5625
rect 10115 5615 10315 5640
rect 10370 5631 10400 5819
rect 10344 5625 10400 5631
rect 10086 5565 10344 5585
rect 10396 5565 10400 5625
rect 10030 5555 10400 5565
rect 10430 5885 10800 5895
rect 10430 5825 10434 5885
rect 10486 5865 10744 5885
rect 10430 5819 10486 5825
rect 10430 5631 10460 5819
rect 10515 5810 10715 5835
rect 10796 5825 10800 5885
rect 10744 5819 10800 5825
rect 10515 5790 10585 5810
rect 10490 5750 10585 5790
rect 10645 5790 10715 5810
rect 10645 5750 10740 5790
rect 10490 5700 10740 5750
rect 10490 5660 10585 5700
rect 10515 5640 10585 5660
rect 10645 5660 10740 5700
rect 10645 5640 10715 5660
rect 10430 5625 10486 5631
rect 10430 5565 10434 5625
rect 10515 5615 10715 5640
rect 10770 5631 10800 5819
rect 10744 5625 10800 5631
rect 10486 5565 10744 5585
rect 10796 5565 10800 5625
rect 10430 5555 10800 5565
rect 10830 5885 11200 5895
rect 10830 5825 10834 5885
rect 10886 5865 11144 5885
rect 10830 5819 10886 5825
rect 10830 5631 10860 5819
rect 10915 5810 11115 5835
rect 11196 5825 11200 5885
rect 11144 5819 11200 5825
rect 10915 5790 10985 5810
rect 10890 5750 10985 5790
rect 11045 5790 11115 5810
rect 11045 5750 11140 5790
rect 10890 5700 11140 5750
rect 10890 5660 10985 5700
rect 10915 5640 10985 5660
rect 11045 5660 11140 5700
rect 11045 5640 11115 5660
rect 10830 5625 10886 5631
rect 10830 5565 10834 5625
rect 10915 5615 11115 5640
rect 11170 5631 11200 5819
rect 11144 5625 11200 5631
rect 10886 5565 11144 5585
rect 11196 5565 11200 5625
rect 10830 5555 11200 5565
rect 11230 5885 11600 5895
rect 11230 5825 11234 5885
rect 11286 5865 11544 5885
rect 11230 5819 11286 5825
rect 11230 5631 11260 5819
rect 11315 5810 11515 5835
rect 11596 5825 11600 5885
rect 11544 5819 11600 5825
rect 11315 5790 11385 5810
rect 11290 5750 11385 5790
rect 11445 5790 11515 5810
rect 11445 5750 11540 5790
rect 11290 5700 11540 5750
rect 11290 5660 11385 5700
rect 11315 5640 11385 5660
rect 11445 5660 11540 5700
rect 11445 5640 11515 5660
rect 11230 5625 11286 5631
rect 11230 5565 11234 5625
rect 11315 5615 11515 5640
rect 11570 5631 11600 5819
rect 11544 5625 11600 5631
rect 11286 5565 11544 5585
rect 11596 5565 11600 5625
rect 11230 5555 11600 5565
rect 11630 5885 12000 5895
rect 11630 5825 11634 5885
rect 11686 5865 11944 5885
rect 11630 5819 11686 5825
rect 11630 5631 11660 5819
rect 11715 5810 11915 5835
rect 11996 5825 12000 5885
rect 11944 5819 12000 5825
rect 11715 5790 11785 5810
rect 11690 5750 11785 5790
rect 11845 5790 11915 5810
rect 11845 5750 11940 5790
rect 11690 5700 11940 5750
rect 11690 5660 11785 5700
rect 11715 5640 11785 5660
rect 11845 5660 11940 5700
rect 11845 5640 11915 5660
rect 11630 5625 11686 5631
rect 11630 5565 11634 5625
rect 11715 5615 11915 5640
rect 11970 5631 12000 5819
rect 11944 5625 12000 5631
rect 11686 5565 11944 5585
rect 11996 5565 12000 5625
rect 11630 5555 12000 5565
rect 12030 5885 12400 5895
rect 12030 5825 12034 5885
rect 12086 5865 12344 5885
rect 12030 5819 12086 5825
rect 12030 5631 12060 5819
rect 12115 5810 12315 5835
rect 12396 5825 12400 5885
rect 12344 5819 12400 5825
rect 12115 5790 12185 5810
rect 12090 5750 12185 5790
rect 12245 5790 12315 5810
rect 12245 5750 12340 5790
rect 12090 5700 12340 5750
rect 12090 5660 12185 5700
rect 12115 5640 12185 5660
rect 12245 5660 12340 5700
rect 12245 5640 12315 5660
rect 12030 5625 12086 5631
rect 12030 5565 12034 5625
rect 12115 5615 12315 5640
rect 12370 5631 12400 5819
rect 12344 5625 12400 5631
rect 12086 5565 12344 5585
rect 12396 5565 12400 5625
rect 12030 5555 12400 5565
rect 12430 5885 12800 5895
rect 12430 5825 12434 5885
rect 12486 5865 12744 5885
rect 12430 5819 12486 5825
rect 12430 5631 12460 5819
rect 12515 5810 12715 5835
rect 12796 5825 12800 5885
rect 12744 5819 12800 5825
rect 12515 5790 12585 5810
rect 12490 5750 12585 5790
rect 12645 5790 12715 5810
rect 12645 5750 12740 5790
rect 12490 5700 12740 5750
rect 12490 5660 12585 5700
rect 12515 5640 12585 5660
rect 12645 5660 12740 5700
rect 12645 5640 12715 5660
rect 12430 5625 12486 5631
rect 12430 5565 12434 5625
rect 12515 5615 12715 5640
rect 12770 5631 12800 5819
rect 12744 5625 12800 5631
rect 12486 5565 12744 5585
rect 12796 5565 12800 5625
rect 12430 5555 12800 5565
rect 12830 5885 13200 5895
rect 12830 5825 12834 5885
rect 12886 5865 13144 5885
rect 12830 5819 12886 5825
rect 12830 5631 12860 5819
rect 12915 5810 13115 5835
rect 13196 5825 13200 5885
rect 13144 5819 13200 5825
rect 12915 5790 12985 5810
rect 12890 5750 12985 5790
rect 13045 5790 13115 5810
rect 13045 5750 13140 5790
rect 12890 5700 13140 5750
rect 12890 5660 12985 5700
rect 12915 5640 12985 5660
rect 13045 5660 13140 5700
rect 13045 5640 13115 5660
rect 12830 5625 12886 5631
rect 12830 5565 12834 5625
rect 12915 5615 13115 5640
rect 13170 5631 13200 5819
rect 13144 5625 13200 5631
rect 12886 5565 13144 5585
rect 13196 5565 13200 5625
rect 12830 5555 13200 5565
rect -370 5515 0 5525
rect -370 5455 -366 5515
rect -314 5495 -56 5515
rect -370 5449 -314 5455
rect -370 5261 -340 5449
rect -285 5440 -85 5465
rect -4 5455 0 5515
rect -56 5449 0 5455
rect -285 5420 -215 5440
rect -310 5380 -215 5420
rect -155 5420 -85 5440
rect -155 5380 -60 5420
rect -310 5330 -60 5380
rect -310 5290 -215 5330
rect -285 5270 -215 5290
rect -155 5290 -60 5330
rect -155 5270 -85 5290
rect -370 5255 -314 5261
rect -370 5195 -366 5255
rect -285 5245 -85 5270
rect -30 5261 0 5449
rect -56 5255 0 5261
rect -314 5195 -56 5215
rect -4 5195 0 5255
rect -370 5185 0 5195
rect 30 5515 400 5525
rect 30 5455 34 5515
rect 86 5495 344 5515
rect 30 5449 86 5455
rect 30 5261 60 5449
rect 115 5440 315 5465
rect 396 5455 400 5515
rect 344 5449 400 5455
rect 115 5420 185 5440
rect 90 5380 185 5420
rect 245 5420 315 5440
rect 245 5380 340 5420
rect 90 5330 340 5380
rect 90 5290 185 5330
rect 115 5270 185 5290
rect 245 5290 340 5330
rect 245 5270 315 5290
rect 30 5255 86 5261
rect 30 5195 34 5255
rect 115 5245 315 5270
rect 370 5261 400 5449
rect 344 5255 400 5261
rect 86 5195 344 5215
rect 396 5195 400 5255
rect 30 5185 400 5195
rect 430 5515 800 5525
rect 430 5455 434 5515
rect 486 5495 744 5515
rect 430 5449 486 5455
rect 430 5261 460 5449
rect 515 5440 715 5465
rect 796 5455 800 5515
rect 744 5449 800 5455
rect 515 5420 585 5440
rect 490 5380 585 5420
rect 645 5420 715 5440
rect 645 5380 740 5420
rect 490 5330 740 5380
rect 490 5290 585 5330
rect 515 5270 585 5290
rect 645 5290 740 5330
rect 645 5270 715 5290
rect 430 5255 486 5261
rect 430 5195 434 5255
rect 515 5245 715 5270
rect 770 5261 800 5449
rect 744 5255 800 5261
rect 486 5195 744 5215
rect 796 5195 800 5255
rect 430 5185 800 5195
rect 830 5515 1200 5525
rect 830 5455 834 5515
rect 886 5495 1144 5515
rect 830 5449 886 5455
rect 830 5261 860 5449
rect 915 5440 1115 5465
rect 1196 5455 1200 5515
rect 1144 5449 1200 5455
rect 915 5420 985 5440
rect 890 5380 985 5420
rect 1045 5420 1115 5440
rect 1045 5380 1140 5420
rect 890 5330 1140 5380
rect 890 5290 985 5330
rect 915 5270 985 5290
rect 1045 5290 1140 5330
rect 1045 5270 1115 5290
rect 830 5255 886 5261
rect 830 5195 834 5255
rect 915 5245 1115 5270
rect 1170 5261 1200 5449
rect 1144 5255 1200 5261
rect 886 5195 1144 5215
rect 1196 5195 1200 5255
rect 830 5185 1200 5195
rect 1230 5515 1600 5525
rect 1230 5455 1234 5515
rect 1286 5495 1544 5515
rect 1230 5449 1286 5455
rect 1230 5261 1260 5449
rect 1315 5440 1515 5465
rect 1596 5455 1600 5515
rect 1544 5449 1600 5455
rect 1315 5420 1385 5440
rect 1290 5380 1385 5420
rect 1445 5420 1515 5440
rect 1445 5380 1540 5420
rect 1290 5330 1540 5380
rect 1290 5290 1385 5330
rect 1315 5270 1385 5290
rect 1445 5290 1540 5330
rect 1445 5270 1515 5290
rect 1230 5255 1286 5261
rect 1230 5195 1234 5255
rect 1315 5245 1515 5270
rect 1570 5261 1600 5449
rect 1544 5255 1600 5261
rect 1286 5195 1544 5215
rect 1596 5195 1600 5255
rect 1230 5185 1600 5195
rect 1630 5515 2000 5525
rect 1630 5455 1634 5515
rect 1686 5495 1944 5515
rect 1630 5449 1686 5455
rect 1630 5261 1660 5449
rect 1715 5440 1915 5465
rect 1996 5455 2000 5515
rect 1944 5449 2000 5455
rect 1715 5420 1785 5440
rect 1690 5380 1785 5420
rect 1845 5420 1915 5440
rect 1845 5380 1940 5420
rect 1690 5330 1940 5380
rect 1690 5290 1785 5330
rect 1715 5270 1785 5290
rect 1845 5290 1940 5330
rect 1845 5270 1915 5290
rect 1630 5255 1686 5261
rect 1630 5195 1634 5255
rect 1715 5245 1915 5270
rect 1970 5261 2000 5449
rect 1944 5255 2000 5261
rect 1686 5195 1944 5215
rect 1996 5195 2000 5255
rect 1630 5185 2000 5195
rect 2030 5515 2400 5525
rect 2030 5455 2034 5515
rect 2086 5495 2344 5515
rect 2030 5449 2086 5455
rect 2030 5261 2060 5449
rect 2115 5440 2315 5465
rect 2396 5455 2400 5515
rect 2344 5449 2400 5455
rect 2115 5420 2185 5440
rect 2090 5380 2185 5420
rect 2245 5420 2315 5440
rect 2245 5380 2340 5420
rect 2090 5330 2340 5380
rect 2090 5290 2185 5330
rect 2115 5270 2185 5290
rect 2245 5290 2340 5330
rect 2245 5270 2315 5290
rect 2030 5255 2086 5261
rect 2030 5195 2034 5255
rect 2115 5245 2315 5270
rect 2370 5261 2400 5449
rect 2344 5255 2400 5261
rect 2086 5195 2344 5215
rect 2396 5195 2400 5255
rect 2030 5185 2400 5195
rect 2430 5515 2800 5525
rect 2430 5455 2434 5515
rect 2486 5495 2744 5515
rect 2430 5449 2486 5455
rect 2430 5261 2460 5449
rect 2515 5440 2715 5465
rect 2796 5455 2800 5515
rect 2744 5449 2800 5455
rect 2515 5420 2585 5440
rect 2490 5380 2585 5420
rect 2645 5420 2715 5440
rect 2645 5380 2740 5420
rect 2490 5330 2740 5380
rect 2490 5290 2585 5330
rect 2515 5270 2585 5290
rect 2645 5290 2740 5330
rect 2645 5270 2715 5290
rect 2430 5255 2486 5261
rect 2430 5195 2434 5255
rect 2515 5245 2715 5270
rect 2770 5261 2800 5449
rect 2744 5255 2800 5261
rect 2486 5195 2744 5215
rect 2796 5195 2800 5255
rect 2430 5185 2800 5195
rect 2830 5515 3200 5525
rect 2830 5455 2834 5515
rect 2886 5495 3144 5515
rect 2830 5449 2886 5455
rect 2830 5261 2860 5449
rect 2915 5440 3115 5465
rect 3196 5455 3200 5515
rect 3144 5449 3200 5455
rect 2915 5420 2985 5440
rect 2890 5380 2985 5420
rect 3045 5420 3115 5440
rect 3045 5380 3140 5420
rect 2890 5330 3140 5380
rect 2890 5290 2985 5330
rect 2915 5270 2985 5290
rect 3045 5290 3140 5330
rect 3045 5270 3115 5290
rect 2830 5255 2886 5261
rect 2830 5195 2834 5255
rect 2915 5245 3115 5270
rect 3170 5261 3200 5449
rect 3144 5255 3200 5261
rect 2886 5195 3144 5215
rect 3196 5195 3200 5255
rect 2830 5185 3200 5195
rect 3230 5515 3600 5525
rect 3230 5455 3234 5515
rect 3286 5495 3544 5515
rect 3230 5449 3286 5455
rect 3230 5261 3260 5449
rect 3315 5440 3515 5465
rect 3596 5455 3600 5515
rect 3544 5449 3600 5455
rect 3315 5420 3385 5440
rect 3290 5380 3385 5420
rect 3445 5420 3515 5440
rect 3445 5380 3540 5420
rect 3290 5330 3540 5380
rect 3290 5290 3385 5330
rect 3315 5270 3385 5290
rect 3445 5290 3540 5330
rect 3445 5270 3515 5290
rect 3230 5255 3286 5261
rect 3230 5195 3234 5255
rect 3315 5245 3515 5270
rect 3570 5261 3600 5449
rect 3544 5255 3600 5261
rect 3286 5195 3544 5215
rect 3596 5195 3600 5255
rect 3230 5185 3600 5195
rect 3630 5515 4000 5525
rect 3630 5455 3634 5515
rect 3686 5495 3944 5515
rect 3630 5449 3686 5455
rect 3630 5261 3660 5449
rect 3715 5440 3915 5465
rect 3996 5455 4000 5515
rect 3944 5449 4000 5455
rect 3715 5420 3785 5440
rect 3690 5380 3785 5420
rect 3845 5420 3915 5440
rect 3845 5380 3940 5420
rect 3690 5330 3940 5380
rect 3690 5290 3785 5330
rect 3715 5270 3785 5290
rect 3845 5290 3940 5330
rect 3845 5270 3915 5290
rect 3630 5255 3686 5261
rect 3630 5195 3634 5255
rect 3715 5245 3915 5270
rect 3970 5261 4000 5449
rect 3944 5255 4000 5261
rect 3686 5195 3944 5215
rect 3996 5195 4000 5255
rect 3630 5185 4000 5195
rect 4030 5515 4400 5525
rect 4030 5455 4034 5515
rect 4086 5495 4344 5515
rect 4030 5449 4086 5455
rect 4030 5261 4060 5449
rect 4115 5440 4315 5465
rect 4396 5455 4400 5515
rect 4344 5449 4400 5455
rect 4115 5420 4185 5440
rect 4090 5380 4185 5420
rect 4245 5420 4315 5440
rect 4245 5380 4340 5420
rect 4090 5330 4340 5380
rect 4090 5290 4185 5330
rect 4115 5270 4185 5290
rect 4245 5290 4340 5330
rect 4245 5270 4315 5290
rect 4030 5255 4086 5261
rect 4030 5195 4034 5255
rect 4115 5245 4315 5270
rect 4370 5261 4400 5449
rect 4344 5255 4400 5261
rect 4086 5195 4344 5215
rect 4396 5195 4400 5255
rect 4030 5185 4400 5195
rect 4430 5515 4800 5525
rect 4430 5455 4434 5515
rect 4486 5495 4744 5515
rect 4430 5449 4486 5455
rect 4430 5261 4460 5449
rect 4515 5440 4715 5465
rect 4796 5455 4800 5515
rect 4744 5449 4800 5455
rect 4515 5420 4585 5440
rect 4490 5380 4585 5420
rect 4645 5420 4715 5440
rect 4645 5380 4740 5420
rect 4490 5330 4740 5380
rect 4490 5290 4585 5330
rect 4515 5270 4585 5290
rect 4645 5290 4740 5330
rect 4645 5270 4715 5290
rect 4430 5255 4486 5261
rect 4430 5195 4434 5255
rect 4515 5245 4715 5270
rect 4770 5261 4800 5449
rect 4744 5255 4800 5261
rect 4486 5195 4744 5215
rect 4796 5195 4800 5255
rect 4430 5185 4800 5195
rect 4830 5515 5200 5525
rect 4830 5455 4834 5515
rect 4886 5495 5144 5515
rect 4830 5449 4886 5455
rect 4830 5261 4860 5449
rect 4915 5440 5115 5465
rect 5196 5455 5200 5515
rect 5144 5449 5200 5455
rect 4915 5420 4985 5440
rect 4890 5380 4985 5420
rect 5045 5420 5115 5440
rect 5045 5380 5140 5420
rect 4890 5330 5140 5380
rect 4890 5290 4985 5330
rect 4915 5270 4985 5290
rect 5045 5290 5140 5330
rect 5045 5270 5115 5290
rect 4830 5255 4886 5261
rect 4830 5195 4834 5255
rect 4915 5245 5115 5270
rect 5170 5261 5200 5449
rect 5144 5255 5200 5261
rect 4886 5195 5144 5215
rect 5196 5195 5200 5255
rect 4830 5185 5200 5195
rect 5230 5515 5600 5525
rect 5230 5455 5234 5515
rect 5286 5495 5544 5515
rect 5230 5449 5286 5455
rect 5230 5261 5260 5449
rect 5315 5440 5515 5465
rect 5596 5455 5600 5515
rect 5544 5449 5600 5455
rect 5315 5420 5385 5440
rect 5290 5380 5385 5420
rect 5445 5420 5515 5440
rect 5445 5380 5540 5420
rect 5290 5330 5540 5380
rect 5290 5290 5385 5330
rect 5315 5270 5385 5290
rect 5445 5290 5540 5330
rect 5445 5270 5515 5290
rect 5230 5255 5286 5261
rect 5230 5195 5234 5255
rect 5315 5245 5515 5270
rect 5570 5261 5600 5449
rect 5544 5255 5600 5261
rect 5286 5195 5544 5215
rect 5596 5195 5600 5255
rect 5230 5185 5600 5195
rect 5630 5515 6000 5525
rect 5630 5455 5634 5515
rect 5686 5495 5944 5515
rect 5630 5449 5686 5455
rect 5630 5261 5660 5449
rect 5715 5440 5915 5465
rect 5996 5455 6000 5515
rect 5944 5449 6000 5455
rect 5715 5420 5785 5440
rect 5690 5380 5785 5420
rect 5845 5420 5915 5440
rect 5845 5380 5940 5420
rect 5690 5330 5940 5380
rect 5690 5290 5785 5330
rect 5715 5270 5785 5290
rect 5845 5290 5940 5330
rect 5845 5270 5915 5290
rect 5630 5255 5686 5261
rect 5630 5195 5634 5255
rect 5715 5245 5915 5270
rect 5970 5261 6000 5449
rect 5944 5255 6000 5261
rect 5686 5195 5944 5215
rect 5996 5195 6000 5255
rect 5630 5185 6000 5195
rect 6030 5515 6400 5525
rect 6030 5455 6034 5515
rect 6086 5495 6344 5515
rect 6030 5449 6086 5455
rect 6030 5261 6060 5449
rect 6115 5440 6315 5465
rect 6396 5455 6400 5515
rect 6344 5449 6400 5455
rect 6115 5420 6185 5440
rect 6090 5380 6185 5420
rect 6245 5420 6315 5440
rect 6245 5380 6340 5420
rect 6090 5330 6340 5380
rect 6090 5290 6185 5330
rect 6115 5270 6185 5290
rect 6245 5290 6340 5330
rect 6245 5270 6315 5290
rect 6030 5255 6086 5261
rect 6030 5195 6034 5255
rect 6115 5245 6315 5270
rect 6370 5261 6400 5449
rect 6344 5255 6400 5261
rect 6086 5195 6344 5215
rect 6396 5195 6400 5255
rect 6030 5185 6400 5195
rect 6430 5515 6800 5525
rect 6430 5455 6434 5515
rect 6486 5495 6744 5515
rect 6430 5449 6486 5455
rect 6430 5261 6460 5449
rect 6515 5440 6715 5465
rect 6796 5455 6800 5515
rect 6744 5449 6800 5455
rect 6515 5420 6585 5440
rect 6490 5380 6585 5420
rect 6645 5420 6715 5440
rect 6645 5380 6740 5420
rect 6490 5330 6740 5380
rect 6490 5290 6585 5330
rect 6515 5270 6585 5290
rect 6645 5290 6740 5330
rect 6645 5270 6715 5290
rect 6430 5255 6486 5261
rect 6430 5195 6434 5255
rect 6515 5245 6715 5270
rect 6770 5261 6800 5449
rect 6744 5255 6800 5261
rect 6486 5195 6744 5215
rect 6796 5195 6800 5255
rect 6430 5185 6800 5195
rect 6830 5515 7200 5525
rect 6830 5455 6834 5515
rect 6886 5495 7144 5515
rect 6830 5449 6886 5455
rect 6830 5261 6860 5449
rect 6915 5440 7115 5465
rect 7196 5455 7200 5515
rect 7144 5449 7200 5455
rect 6915 5420 6985 5440
rect 6890 5380 6985 5420
rect 7045 5420 7115 5440
rect 7045 5380 7140 5420
rect 6890 5330 7140 5380
rect 6890 5290 6985 5330
rect 6915 5270 6985 5290
rect 7045 5290 7140 5330
rect 7045 5270 7115 5290
rect 6830 5255 6886 5261
rect 6830 5195 6834 5255
rect 6915 5245 7115 5270
rect 7170 5261 7200 5449
rect 7144 5255 7200 5261
rect 6886 5195 7144 5215
rect 7196 5195 7200 5255
rect 6830 5185 7200 5195
rect 7230 5515 7600 5525
rect 7230 5455 7234 5515
rect 7286 5495 7544 5515
rect 7230 5449 7286 5455
rect 7230 5261 7260 5449
rect 7315 5440 7515 5465
rect 7596 5455 7600 5515
rect 7544 5449 7600 5455
rect 7315 5420 7385 5440
rect 7290 5380 7385 5420
rect 7445 5420 7515 5440
rect 7445 5380 7540 5420
rect 7290 5330 7540 5380
rect 7290 5290 7385 5330
rect 7315 5270 7385 5290
rect 7445 5290 7540 5330
rect 7445 5270 7515 5290
rect 7230 5255 7286 5261
rect 7230 5195 7234 5255
rect 7315 5245 7515 5270
rect 7570 5261 7600 5449
rect 7544 5255 7600 5261
rect 7286 5195 7544 5215
rect 7596 5195 7600 5255
rect 7230 5185 7600 5195
rect 7630 5515 8000 5525
rect 7630 5455 7634 5515
rect 7686 5495 7944 5515
rect 7630 5449 7686 5455
rect 7630 5261 7660 5449
rect 7715 5440 7915 5465
rect 7996 5455 8000 5515
rect 7944 5449 8000 5455
rect 7715 5420 7785 5440
rect 7690 5380 7785 5420
rect 7845 5420 7915 5440
rect 7845 5380 7940 5420
rect 7690 5330 7940 5380
rect 7690 5290 7785 5330
rect 7715 5270 7785 5290
rect 7845 5290 7940 5330
rect 7845 5270 7915 5290
rect 7630 5255 7686 5261
rect 7630 5195 7634 5255
rect 7715 5245 7915 5270
rect 7970 5261 8000 5449
rect 7944 5255 8000 5261
rect 7686 5195 7944 5215
rect 7996 5195 8000 5255
rect 7630 5185 8000 5195
rect 8030 5515 8400 5525
rect 8030 5455 8034 5515
rect 8086 5495 8344 5515
rect 8030 5449 8086 5455
rect 8030 5261 8060 5449
rect 8115 5440 8315 5465
rect 8396 5455 8400 5515
rect 8344 5449 8400 5455
rect 8115 5420 8185 5440
rect 8090 5380 8185 5420
rect 8245 5420 8315 5440
rect 8245 5380 8340 5420
rect 8090 5330 8340 5380
rect 8090 5290 8185 5330
rect 8115 5270 8185 5290
rect 8245 5290 8340 5330
rect 8245 5270 8315 5290
rect 8030 5255 8086 5261
rect 8030 5195 8034 5255
rect 8115 5245 8315 5270
rect 8370 5261 8400 5449
rect 8344 5255 8400 5261
rect 8086 5195 8344 5215
rect 8396 5195 8400 5255
rect 8030 5185 8400 5195
rect 8430 5515 8800 5525
rect 8430 5455 8434 5515
rect 8486 5495 8744 5515
rect 8430 5449 8486 5455
rect 8430 5261 8460 5449
rect 8515 5440 8715 5465
rect 8796 5455 8800 5515
rect 8744 5449 8800 5455
rect 8515 5420 8585 5440
rect 8490 5380 8585 5420
rect 8645 5420 8715 5440
rect 8645 5380 8740 5420
rect 8490 5330 8740 5380
rect 8490 5290 8585 5330
rect 8515 5270 8585 5290
rect 8645 5290 8740 5330
rect 8645 5270 8715 5290
rect 8430 5255 8486 5261
rect 8430 5195 8434 5255
rect 8515 5245 8715 5270
rect 8770 5261 8800 5449
rect 8744 5255 8800 5261
rect 8486 5195 8744 5215
rect 8796 5195 8800 5255
rect 8430 5185 8800 5195
rect 8830 5515 9200 5525
rect 8830 5455 8834 5515
rect 8886 5495 9144 5515
rect 8830 5449 8886 5455
rect 8830 5261 8860 5449
rect 8915 5440 9115 5465
rect 9196 5455 9200 5515
rect 9144 5449 9200 5455
rect 8915 5420 8985 5440
rect 8890 5380 8985 5420
rect 9045 5420 9115 5440
rect 9045 5380 9140 5420
rect 8890 5330 9140 5380
rect 8890 5290 8985 5330
rect 8915 5270 8985 5290
rect 9045 5290 9140 5330
rect 9045 5270 9115 5290
rect 8830 5255 8886 5261
rect 8830 5195 8834 5255
rect 8915 5245 9115 5270
rect 9170 5261 9200 5449
rect 9144 5255 9200 5261
rect 8886 5195 9144 5215
rect 9196 5195 9200 5255
rect 8830 5185 9200 5195
rect 9230 5515 9600 5525
rect 9230 5455 9234 5515
rect 9286 5495 9544 5515
rect 9230 5449 9286 5455
rect 9230 5261 9260 5449
rect 9315 5440 9515 5465
rect 9596 5455 9600 5515
rect 9544 5449 9600 5455
rect 9315 5420 9385 5440
rect 9290 5380 9385 5420
rect 9445 5420 9515 5440
rect 9445 5380 9540 5420
rect 9290 5330 9540 5380
rect 9290 5290 9385 5330
rect 9315 5270 9385 5290
rect 9445 5290 9540 5330
rect 9445 5270 9515 5290
rect 9230 5255 9286 5261
rect 9230 5195 9234 5255
rect 9315 5245 9515 5270
rect 9570 5261 9600 5449
rect 9544 5255 9600 5261
rect 9286 5195 9544 5215
rect 9596 5195 9600 5255
rect 9230 5185 9600 5195
rect 9630 5515 10000 5525
rect 9630 5455 9634 5515
rect 9686 5495 9944 5515
rect 9630 5449 9686 5455
rect 9630 5261 9660 5449
rect 9715 5440 9915 5465
rect 9996 5455 10000 5515
rect 9944 5449 10000 5455
rect 9715 5420 9785 5440
rect 9690 5380 9785 5420
rect 9845 5420 9915 5440
rect 9845 5380 9940 5420
rect 9690 5330 9940 5380
rect 9690 5290 9785 5330
rect 9715 5270 9785 5290
rect 9845 5290 9940 5330
rect 9845 5270 9915 5290
rect 9630 5255 9686 5261
rect 9630 5195 9634 5255
rect 9715 5245 9915 5270
rect 9970 5261 10000 5449
rect 9944 5255 10000 5261
rect 9686 5195 9944 5215
rect 9996 5195 10000 5255
rect 9630 5185 10000 5195
rect 10030 5515 10400 5525
rect 10030 5455 10034 5515
rect 10086 5495 10344 5515
rect 10030 5449 10086 5455
rect 10030 5261 10060 5449
rect 10115 5440 10315 5465
rect 10396 5455 10400 5515
rect 10344 5449 10400 5455
rect 10115 5420 10185 5440
rect 10090 5380 10185 5420
rect 10245 5420 10315 5440
rect 10245 5380 10340 5420
rect 10090 5330 10340 5380
rect 10090 5290 10185 5330
rect 10115 5270 10185 5290
rect 10245 5290 10340 5330
rect 10245 5270 10315 5290
rect 10030 5255 10086 5261
rect 10030 5195 10034 5255
rect 10115 5245 10315 5270
rect 10370 5261 10400 5449
rect 10344 5255 10400 5261
rect 10086 5195 10344 5215
rect 10396 5195 10400 5255
rect 10030 5185 10400 5195
rect 10430 5515 10800 5525
rect 10430 5455 10434 5515
rect 10486 5495 10744 5515
rect 10430 5449 10486 5455
rect 10430 5261 10460 5449
rect 10515 5440 10715 5465
rect 10796 5455 10800 5515
rect 10744 5449 10800 5455
rect 10515 5420 10585 5440
rect 10490 5380 10585 5420
rect 10645 5420 10715 5440
rect 10645 5380 10740 5420
rect 10490 5330 10740 5380
rect 10490 5290 10585 5330
rect 10515 5270 10585 5290
rect 10645 5290 10740 5330
rect 10645 5270 10715 5290
rect 10430 5255 10486 5261
rect 10430 5195 10434 5255
rect 10515 5245 10715 5270
rect 10770 5261 10800 5449
rect 10744 5255 10800 5261
rect 10486 5195 10744 5215
rect 10796 5195 10800 5255
rect 10430 5185 10800 5195
rect 10830 5515 11200 5525
rect 10830 5455 10834 5515
rect 10886 5495 11144 5515
rect 10830 5449 10886 5455
rect 10830 5261 10860 5449
rect 10915 5440 11115 5465
rect 11196 5455 11200 5515
rect 11144 5449 11200 5455
rect 10915 5420 10985 5440
rect 10890 5380 10985 5420
rect 11045 5420 11115 5440
rect 11045 5380 11140 5420
rect 10890 5330 11140 5380
rect 10890 5290 10985 5330
rect 10915 5270 10985 5290
rect 11045 5290 11140 5330
rect 11045 5270 11115 5290
rect 10830 5255 10886 5261
rect 10830 5195 10834 5255
rect 10915 5245 11115 5270
rect 11170 5261 11200 5449
rect 11144 5255 11200 5261
rect 10886 5195 11144 5215
rect 11196 5195 11200 5255
rect 10830 5185 11200 5195
rect 11230 5515 11600 5525
rect 11230 5455 11234 5515
rect 11286 5495 11544 5515
rect 11230 5449 11286 5455
rect 11230 5261 11260 5449
rect 11315 5440 11515 5465
rect 11596 5455 11600 5515
rect 11544 5449 11600 5455
rect 11315 5420 11385 5440
rect 11290 5380 11385 5420
rect 11445 5420 11515 5440
rect 11445 5380 11540 5420
rect 11290 5330 11540 5380
rect 11290 5290 11385 5330
rect 11315 5270 11385 5290
rect 11445 5290 11540 5330
rect 11445 5270 11515 5290
rect 11230 5255 11286 5261
rect 11230 5195 11234 5255
rect 11315 5245 11515 5270
rect 11570 5261 11600 5449
rect 11544 5255 11600 5261
rect 11286 5195 11544 5215
rect 11596 5195 11600 5255
rect 11230 5185 11600 5195
rect 11630 5515 12000 5525
rect 11630 5455 11634 5515
rect 11686 5495 11944 5515
rect 11630 5449 11686 5455
rect 11630 5261 11660 5449
rect 11715 5440 11915 5465
rect 11996 5455 12000 5515
rect 11944 5449 12000 5455
rect 11715 5420 11785 5440
rect 11690 5380 11785 5420
rect 11845 5420 11915 5440
rect 11845 5380 11940 5420
rect 11690 5330 11940 5380
rect 11690 5290 11785 5330
rect 11715 5270 11785 5290
rect 11845 5290 11940 5330
rect 11845 5270 11915 5290
rect 11630 5255 11686 5261
rect 11630 5195 11634 5255
rect 11715 5245 11915 5270
rect 11970 5261 12000 5449
rect 11944 5255 12000 5261
rect 11686 5195 11944 5215
rect 11996 5195 12000 5255
rect 11630 5185 12000 5195
rect 12030 5515 12400 5525
rect 12030 5455 12034 5515
rect 12086 5495 12344 5515
rect 12030 5449 12086 5455
rect 12030 5261 12060 5449
rect 12115 5440 12315 5465
rect 12396 5455 12400 5515
rect 12344 5449 12400 5455
rect 12115 5420 12185 5440
rect 12090 5380 12185 5420
rect 12245 5420 12315 5440
rect 12245 5380 12340 5420
rect 12090 5330 12340 5380
rect 12090 5290 12185 5330
rect 12115 5270 12185 5290
rect 12245 5290 12340 5330
rect 12245 5270 12315 5290
rect 12030 5255 12086 5261
rect 12030 5195 12034 5255
rect 12115 5245 12315 5270
rect 12370 5261 12400 5449
rect 12344 5255 12400 5261
rect 12086 5195 12344 5215
rect 12396 5195 12400 5255
rect 12030 5185 12400 5195
rect 12430 5515 12800 5525
rect 12430 5455 12434 5515
rect 12486 5495 12744 5515
rect 12430 5449 12486 5455
rect 12430 5261 12460 5449
rect 12515 5440 12715 5465
rect 12796 5455 12800 5515
rect 12744 5449 12800 5455
rect 12515 5420 12585 5440
rect 12490 5380 12585 5420
rect 12645 5420 12715 5440
rect 12645 5380 12740 5420
rect 12490 5330 12740 5380
rect 12490 5290 12585 5330
rect 12515 5270 12585 5290
rect 12645 5290 12740 5330
rect 12645 5270 12715 5290
rect 12430 5255 12486 5261
rect 12430 5195 12434 5255
rect 12515 5245 12715 5270
rect 12770 5261 12800 5449
rect 12744 5255 12800 5261
rect 12486 5195 12744 5215
rect 12796 5195 12800 5255
rect 12430 5185 12800 5195
rect 12830 5515 13200 5525
rect 12830 5455 12834 5515
rect 12886 5495 13144 5515
rect 12830 5449 12886 5455
rect 12830 5261 12860 5449
rect 12915 5440 13115 5465
rect 13196 5455 13200 5515
rect 13144 5449 13200 5455
rect 12915 5420 12985 5440
rect 12890 5380 12985 5420
rect 13045 5420 13115 5440
rect 13045 5380 13140 5420
rect 12890 5330 13140 5380
rect 12890 5290 12985 5330
rect 12915 5270 12985 5290
rect 13045 5290 13140 5330
rect 13045 5270 13115 5290
rect 12830 5255 12886 5261
rect 12830 5195 12834 5255
rect 12915 5245 13115 5270
rect 13170 5261 13200 5449
rect 13144 5255 13200 5261
rect 12886 5195 13144 5215
rect 13196 5195 13200 5255
rect 12830 5185 13200 5195
rect -370 5145 0 5155
rect -370 5085 -366 5145
rect -314 5125 -56 5145
rect -370 5079 -314 5085
rect -370 4891 -340 5079
rect -285 5070 -85 5095
rect -4 5085 0 5145
rect -56 5079 0 5085
rect -285 5050 -215 5070
rect -310 5010 -215 5050
rect -155 5050 -85 5070
rect -155 5010 -60 5050
rect -310 4960 -60 5010
rect -310 4920 -215 4960
rect -285 4900 -215 4920
rect -155 4920 -60 4960
rect -155 4900 -85 4920
rect -370 4885 -314 4891
rect -370 4825 -366 4885
rect -285 4875 -85 4900
rect -30 4891 0 5079
rect -56 4885 0 4891
rect -314 4825 -56 4845
rect -4 4825 0 4885
rect -370 4815 0 4825
rect 30 5145 400 5155
rect 30 5085 34 5145
rect 86 5125 344 5145
rect 30 5079 86 5085
rect 30 4891 60 5079
rect 115 5070 315 5095
rect 396 5085 400 5145
rect 344 5079 400 5085
rect 115 5050 185 5070
rect 90 5010 185 5050
rect 245 5050 315 5070
rect 245 5010 340 5050
rect 90 4960 340 5010
rect 90 4920 185 4960
rect 115 4900 185 4920
rect 245 4920 340 4960
rect 245 4900 315 4920
rect 30 4885 86 4891
rect 30 4825 34 4885
rect 115 4875 315 4900
rect 370 4891 400 5079
rect 344 4885 400 4891
rect 86 4825 344 4845
rect 396 4825 400 4885
rect 30 4815 400 4825
rect 430 5145 800 5155
rect 430 5085 434 5145
rect 486 5125 744 5145
rect 430 5079 486 5085
rect 430 4891 460 5079
rect 515 5070 715 5095
rect 796 5085 800 5145
rect 744 5079 800 5085
rect 515 5050 585 5070
rect 490 5010 585 5050
rect 645 5050 715 5070
rect 645 5010 740 5050
rect 490 4960 740 5010
rect 490 4920 585 4960
rect 515 4900 585 4920
rect 645 4920 740 4960
rect 645 4900 715 4920
rect 430 4885 486 4891
rect 430 4825 434 4885
rect 515 4875 715 4900
rect 770 4891 800 5079
rect 744 4885 800 4891
rect 486 4825 744 4845
rect 796 4825 800 4885
rect 430 4815 800 4825
rect 830 5145 1200 5155
rect 830 5085 834 5145
rect 886 5125 1144 5145
rect 830 5079 886 5085
rect 830 4891 860 5079
rect 915 5070 1115 5095
rect 1196 5085 1200 5145
rect 1144 5079 1200 5085
rect 915 5050 985 5070
rect 890 5010 985 5050
rect 1045 5050 1115 5070
rect 1045 5010 1140 5050
rect 890 4960 1140 5010
rect 890 4920 985 4960
rect 915 4900 985 4920
rect 1045 4920 1140 4960
rect 1045 4900 1115 4920
rect 830 4885 886 4891
rect 830 4825 834 4885
rect 915 4875 1115 4900
rect 1170 4891 1200 5079
rect 1144 4885 1200 4891
rect 886 4825 1144 4845
rect 1196 4825 1200 4885
rect 830 4815 1200 4825
rect 1230 5145 1600 5155
rect 1230 5085 1234 5145
rect 1286 5125 1544 5145
rect 1230 5079 1286 5085
rect 1230 4891 1260 5079
rect 1315 5070 1515 5095
rect 1596 5085 1600 5145
rect 1544 5079 1600 5085
rect 1315 5050 1385 5070
rect 1290 5010 1385 5050
rect 1445 5050 1515 5070
rect 1445 5010 1540 5050
rect 1290 4960 1540 5010
rect 1290 4920 1385 4960
rect 1315 4900 1385 4920
rect 1445 4920 1540 4960
rect 1445 4900 1515 4920
rect 1230 4885 1286 4891
rect 1230 4825 1234 4885
rect 1315 4875 1515 4900
rect 1570 4891 1600 5079
rect 1544 4885 1600 4891
rect 1286 4825 1544 4845
rect 1596 4825 1600 4885
rect 1230 4815 1600 4825
rect 1630 5145 2000 5155
rect 1630 5085 1634 5145
rect 1686 5125 1944 5145
rect 1630 5079 1686 5085
rect 1630 4891 1660 5079
rect 1715 5070 1915 5095
rect 1996 5085 2000 5145
rect 1944 5079 2000 5085
rect 1715 5050 1785 5070
rect 1690 5010 1785 5050
rect 1845 5050 1915 5070
rect 1845 5010 1940 5050
rect 1690 4960 1940 5010
rect 1690 4920 1785 4960
rect 1715 4900 1785 4920
rect 1845 4920 1940 4960
rect 1845 4900 1915 4920
rect 1630 4885 1686 4891
rect 1630 4825 1634 4885
rect 1715 4875 1915 4900
rect 1970 4891 2000 5079
rect 1944 4885 2000 4891
rect 1686 4825 1944 4845
rect 1996 4825 2000 4885
rect 1630 4815 2000 4825
rect 2030 5145 2400 5155
rect 2030 5085 2034 5145
rect 2086 5125 2344 5145
rect 2030 5079 2086 5085
rect 2030 4891 2060 5079
rect 2115 5070 2315 5095
rect 2396 5085 2400 5145
rect 2344 5079 2400 5085
rect 2115 5050 2185 5070
rect 2090 5010 2185 5050
rect 2245 5050 2315 5070
rect 2245 5010 2340 5050
rect 2090 4960 2340 5010
rect 2090 4920 2185 4960
rect 2115 4900 2185 4920
rect 2245 4920 2340 4960
rect 2245 4900 2315 4920
rect 2030 4885 2086 4891
rect 2030 4825 2034 4885
rect 2115 4875 2315 4900
rect 2370 4891 2400 5079
rect 2344 4885 2400 4891
rect 2086 4825 2344 4845
rect 2396 4825 2400 4885
rect 2030 4815 2400 4825
rect 2430 5145 2800 5155
rect 2430 5085 2434 5145
rect 2486 5125 2744 5145
rect 2430 5079 2486 5085
rect 2430 4891 2460 5079
rect 2515 5070 2715 5095
rect 2796 5085 2800 5145
rect 2744 5079 2800 5085
rect 2515 5050 2585 5070
rect 2490 5010 2585 5050
rect 2645 5050 2715 5070
rect 2645 5010 2740 5050
rect 2490 4960 2740 5010
rect 2490 4920 2585 4960
rect 2515 4900 2585 4920
rect 2645 4920 2740 4960
rect 2645 4900 2715 4920
rect 2430 4885 2486 4891
rect 2430 4825 2434 4885
rect 2515 4875 2715 4900
rect 2770 4891 2800 5079
rect 2744 4885 2800 4891
rect 2486 4825 2744 4845
rect 2796 4825 2800 4885
rect 2430 4815 2800 4825
rect 2830 5145 3200 5155
rect 2830 5085 2834 5145
rect 2886 5125 3144 5145
rect 2830 5079 2886 5085
rect 2830 4891 2860 5079
rect 2915 5070 3115 5095
rect 3196 5085 3200 5145
rect 3144 5079 3200 5085
rect 2915 5050 2985 5070
rect 2890 5010 2985 5050
rect 3045 5050 3115 5070
rect 3045 5010 3140 5050
rect 2890 4960 3140 5010
rect 2890 4920 2985 4960
rect 2915 4900 2985 4920
rect 3045 4920 3140 4960
rect 3045 4900 3115 4920
rect 2830 4885 2886 4891
rect 2830 4825 2834 4885
rect 2915 4875 3115 4900
rect 3170 4891 3200 5079
rect 3144 4885 3200 4891
rect 2886 4825 3144 4845
rect 3196 4825 3200 4885
rect 2830 4815 3200 4825
rect 3230 5145 3600 5155
rect 3230 5085 3234 5145
rect 3286 5125 3544 5145
rect 3230 5079 3286 5085
rect 3230 4891 3260 5079
rect 3315 5070 3515 5095
rect 3596 5085 3600 5145
rect 3544 5079 3600 5085
rect 3315 5050 3385 5070
rect 3290 5010 3385 5050
rect 3445 5050 3515 5070
rect 3445 5010 3540 5050
rect 3290 4960 3540 5010
rect 3290 4920 3385 4960
rect 3315 4900 3385 4920
rect 3445 4920 3540 4960
rect 3445 4900 3515 4920
rect 3230 4885 3286 4891
rect 3230 4825 3234 4885
rect 3315 4875 3515 4900
rect 3570 4891 3600 5079
rect 3544 4885 3600 4891
rect 3286 4825 3544 4845
rect 3596 4825 3600 4885
rect 3230 4815 3600 4825
rect 3630 5145 4000 5155
rect 3630 5085 3634 5145
rect 3686 5125 3944 5145
rect 3630 5079 3686 5085
rect 3630 4891 3660 5079
rect 3715 5070 3915 5095
rect 3996 5085 4000 5145
rect 3944 5079 4000 5085
rect 3715 5050 3785 5070
rect 3690 5010 3785 5050
rect 3845 5050 3915 5070
rect 3845 5010 3940 5050
rect 3690 4960 3940 5010
rect 3690 4920 3785 4960
rect 3715 4900 3785 4920
rect 3845 4920 3940 4960
rect 3845 4900 3915 4920
rect 3630 4885 3686 4891
rect 3630 4825 3634 4885
rect 3715 4875 3915 4900
rect 3970 4891 4000 5079
rect 3944 4885 4000 4891
rect 3686 4825 3944 4845
rect 3996 4825 4000 4885
rect 3630 4815 4000 4825
rect 4030 5145 4400 5155
rect 4030 5085 4034 5145
rect 4086 5125 4344 5145
rect 4030 5079 4086 5085
rect 4030 4891 4060 5079
rect 4115 5070 4315 5095
rect 4396 5085 4400 5145
rect 4344 5079 4400 5085
rect 4115 5050 4185 5070
rect 4090 5010 4185 5050
rect 4245 5050 4315 5070
rect 4245 5010 4340 5050
rect 4090 4960 4340 5010
rect 4090 4920 4185 4960
rect 4115 4900 4185 4920
rect 4245 4920 4340 4960
rect 4245 4900 4315 4920
rect 4030 4885 4086 4891
rect 4030 4825 4034 4885
rect 4115 4875 4315 4900
rect 4370 4891 4400 5079
rect 4344 4885 4400 4891
rect 4086 4825 4344 4845
rect 4396 4825 4400 4885
rect 4030 4815 4400 4825
rect 4430 5145 4800 5155
rect 4430 5085 4434 5145
rect 4486 5125 4744 5145
rect 4430 5079 4486 5085
rect 4430 4891 4460 5079
rect 4515 5070 4715 5095
rect 4796 5085 4800 5145
rect 4744 5079 4800 5085
rect 4515 5050 4585 5070
rect 4490 5010 4585 5050
rect 4645 5050 4715 5070
rect 4645 5010 4740 5050
rect 4490 4960 4740 5010
rect 4490 4920 4585 4960
rect 4515 4900 4585 4920
rect 4645 4920 4740 4960
rect 4645 4900 4715 4920
rect 4430 4885 4486 4891
rect 4430 4825 4434 4885
rect 4515 4875 4715 4900
rect 4770 4891 4800 5079
rect 4744 4885 4800 4891
rect 4486 4825 4744 4845
rect 4796 4825 4800 4885
rect 4430 4815 4800 4825
rect 4830 5145 5200 5155
rect 4830 5085 4834 5145
rect 4886 5125 5144 5145
rect 4830 5079 4886 5085
rect 4830 4891 4860 5079
rect 4915 5070 5115 5095
rect 5196 5085 5200 5145
rect 5144 5079 5200 5085
rect 4915 5050 4985 5070
rect 4890 5010 4985 5050
rect 5045 5050 5115 5070
rect 5045 5010 5140 5050
rect 4890 4960 5140 5010
rect 4890 4920 4985 4960
rect 4915 4900 4985 4920
rect 5045 4920 5140 4960
rect 5045 4900 5115 4920
rect 4830 4885 4886 4891
rect 4830 4825 4834 4885
rect 4915 4875 5115 4900
rect 5170 4891 5200 5079
rect 5144 4885 5200 4891
rect 4886 4825 5144 4845
rect 5196 4825 5200 4885
rect 4830 4815 5200 4825
rect 5230 5145 5600 5155
rect 5230 5085 5234 5145
rect 5286 5125 5544 5145
rect 5230 5079 5286 5085
rect 5230 4891 5260 5079
rect 5315 5070 5515 5095
rect 5596 5085 5600 5145
rect 5544 5079 5600 5085
rect 5315 5050 5385 5070
rect 5290 5010 5385 5050
rect 5445 5050 5515 5070
rect 5445 5010 5540 5050
rect 5290 4960 5540 5010
rect 5290 4920 5385 4960
rect 5315 4900 5385 4920
rect 5445 4920 5540 4960
rect 5445 4900 5515 4920
rect 5230 4885 5286 4891
rect 5230 4825 5234 4885
rect 5315 4875 5515 4900
rect 5570 4891 5600 5079
rect 5544 4885 5600 4891
rect 5286 4825 5544 4845
rect 5596 4825 5600 4885
rect 5230 4815 5600 4825
rect 5630 5145 6000 5155
rect 5630 5085 5634 5145
rect 5686 5125 5944 5145
rect 5630 5079 5686 5085
rect 5630 4891 5660 5079
rect 5715 5070 5915 5095
rect 5996 5085 6000 5145
rect 5944 5079 6000 5085
rect 5715 5050 5785 5070
rect 5690 5010 5785 5050
rect 5845 5050 5915 5070
rect 5845 5010 5940 5050
rect 5690 4960 5940 5010
rect 5690 4920 5785 4960
rect 5715 4900 5785 4920
rect 5845 4920 5940 4960
rect 5845 4900 5915 4920
rect 5630 4885 5686 4891
rect 5630 4825 5634 4885
rect 5715 4875 5915 4900
rect 5970 4891 6000 5079
rect 5944 4885 6000 4891
rect 5686 4825 5944 4845
rect 5996 4825 6000 4885
rect 5630 4815 6000 4825
rect 6030 5145 6400 5155
rect 6030 5085 6034 5145
rect 6086 5125 6344 5145
rect 6030 5079 6086 5085
rect 6030 4891 6060 5079
rect 6115 5070 6315 5095
rect 6396 5085 6400 5145
rect 6344 5079 6400 5085
rect 6115 5050 6185 5070
rect 6090 5010 6185 5050
rect 6245 5050 6315 5070
rect 6245 5010 6340 5050
rect 6090 4960 6340 5010
rect 6090 4920 6185 4960
rect 6115 4900 6185 4920
rect 6245 4920 6340 4960
rect 6245 4900 6315 4920
rect 6030 4885 6086 4891
rect 6030 4825 6034 4885
rect 6115 4875 6315 4900
rect 6370 4891 6400 5079
rect 6344 4885 6400 4891
rect 6086 4825 6344 4845
rect 6396 4825 6400 4885
rect 6030 4815 6400 4825
rect 6430 5145 6800 5155
rect 6430 5085 6434 5145
rect 6486 5125 6744 5145
rect 6430 5079 6486 5085
rect 6430 4891 6460 5079
rect 6515 5070 6715 5095
rect 6796 5085 6800 5145
rect 6744 5079 6800 5085
rect 6515 5050 6585 5070
rect 6490 5010 6585 5050
rect 6645 5050 6715 5070
rect 6645 5010 6740 5050
rect 6490 4960 6740 5010
rect 6490 4920 6585 4960
rect 6515 4900 6585 4920
rect 6645 4920 6740 4960
rect 6645 4900 6715 4920
rect 6430 4885 6486 4891
rect 6430 4825 6434 4885
rect 6515 4875 6715 4900
rect 6770 4891 6800 5079
rect 6744 4885 6800 4891
rect 6486 4825 6744 4845
rect 6796 4825 6800 4885
rect 6430 4815 6800 4825
rect 6830 5145 7200 5155
rect 6830 5085 6834 5145
rect 6886 5125 7144 5145
rect 6830 5079 6886 5085
rect 6830 4891 6860 5079
rect 6915 5070 7115 5095
rect 7196 5085 7200 5145
rect 7144 5079 7200 5085
rect 6915 5050 6985 5070
rect 6890 5010 6985 5050
rect 7045 5050 7115 5070
rect 7045 5010 7140 5050
rect 6890 4960 7140 5010
rect 6890 4920 6985 4960
rect 6915 4900 6985 4920
rect 7045 4920 7140 4960
rect 7045 4900 7115 4920
rect 6830 4885 6886 4891
rect 6830 4825 6834 4885
rect 6915 4875 7115 4900
rect 7170 4891 7200 5079
rect 7144 4885 7200 4891
rect 6886 4825 7144 4845
rect 7196 4825 7200 4885
rect 6830 4815 7200 4825
rect 7230 5145 7600 5155
rect 7230 5085 7234 5145
rect 7286 5125 7544 5145
rect 7230 5079 7286 5085
rect 7230 4891 7260 5079
rect 7315 5070 7515 5095
rect 7596 5085 7600 5145
rect 7544 5079 7600 5085
rect 7315 5050 7385 5070
rect 7290 5010 7385 5050
rect 7445 5050 7515 5070
rect 7445 5010 7540 5050
rect 7290 4960 7540 5010
rect 7290 4920 7385 4960
rect 7315 4900 7385 4920
rect 7445 4920 7540 4960
rect 7445 4900 7515 4920
rect 7230 4885 7286 4891
rect 7230 4825 7234 4885
rect 7315 4875 7515 4900
rect 7570 4891 7600 5079
rect 7544 4885 7600 4891
rect 7286 4825 7544 4845
rect 7596 4825 7600 4885
rect 7230 4815 7600 4825
rect 7630 5145 8000 5155
rect 7630 5085 7634 5145
rect 7686 5125 7944 5145
rect 7630 5079 7686 5085
rect 7630 4891 7660 5079
rect 7715 5070 7915 5095
rect 7996 5085 8000 5145
rect 7944 5079 8000 5085
rect 7715 5050 7785 5070
rect 7690 5010 7785 5050
rect 7845 5050 7915 5070
rect 7845 5010 7940 5050
rect 7690 4960 7940 5010
rect 7690 4920 7785 4960
rect 7715 4900 7785 4920
rect 7845 4920 7940 4960
rect 7845 4900 7915 4920
rect 7630 4885 7686 4891
rect 7630 4825 7634 4885
rect 7715 4875 7915 4900
rect 7970 4891 8000 5079
rect 7944 4885 8000 4891
rect 7686 4825 7944 4845
rect 7996 4825 8000 4885
rect 7630 4815 8000 4825
rect 8030 5145 8400 5155
rect 8030 5085 8034 5145
rect 8086 5125 8344 5145
rect 8030 5079 8086 5085
rect 8030 4891 8060 5079
rect 8115 5070 8315 5095
rect 8396 5085 8400 5145
rect 8344 5079 8400 5085
rect 8115 5050 8185 5070
rect 8090 5010 8185 5050
rect 8245 5050 8315 5070
rect 8245 5010 8340 5050
rect 8090 4960 8340 5010
rect 8090 4920 8185 4960
rect 8115 4900 8185 4920
rect 8245 4920 8340 4960
rect 8245 4900 8315 4920
rect 8030 4885 8086 4891
rect 8030 4825 8034 4885
rect 8115 4875 8315 4900
rect 8370 4891 8400 5079
rect 8344 4885 8400 4891
rect 8086 4825 8344 4845
rect 8396 4825 8400 4885
rect 8030 4815 8400 4825
rect 8430 5145 8800 5155
rect 8430 5085 8434 5145
rect 8486 5125 8744 5145
rect 8430 5079 8486 5085
rect 8430 4891 8460 5079
rect 8515 5070 8715 5095
rect 8796 5085 8800 5145
rect 8744 5079 8800 5085
rect 8515 5050 8585 5070
rect 8490 5010 8585 5050
rect 8645 5050 8715 5070
rect 8645 5010 8740 5050
rect 8490 4960 8740 5010
rect 8490 4920 8585 4960
rect 8515 4900 8585 4920
rect 8645 4920 8740 4960
rect 8645 4900 8715 4920
rect 8430 4885 8486 4891
rect 8430 4825 8434 4885
rect 8515 4875 8715 4900
rect 8770 4891 8800 5079
rect 8744 4885 8800 4891
rect 8486 4825 8744 4845
rect 8796 4825 8800 4885
rect 8430 4815 8800 4825
rect 8830 5145 9200 5155
rect 8830 5085 8834 5145
rect 8886 5125 9144 5145
rect 8830 5079 8886 5085
rect 8830 4891 8860 5079
rect 8915 5070 9115 5095
rect 9196 5085 9200 5145
rect 9144 5079 9200 5085
rect 8915 5050 8985 5070
rect 8890 5010 8985 5050
rect 9045 5050 9115 5070
rect 9045 5010 9140 5050
rect 8890 4960 9140 5010
rect 8890 4920 8985 4960
rect 8915 4900 8985 4920
rect 9045 4920 9140 4960
rect 9045 4900 9115 4920
rect 8830 4885 8886 4891
rect 8830 4825 8834 4885
rect 8915 4875 9115 4900
rect 9170 4891 9200 5079
rect 9144 4885 9200 4891
rect 8886 4825 9144 4845
rect 9196 4825 9200 4885
rect 8830 4815 9200 4825
rect 9230 5145 9600 5155
rect 9230 5085 9234 5145
rect 9286 5125 9544 5145
rect 9230 5079 9286 5085
rect 9230 4891 9260 5079
rect 9315 5070 9515 5095
rect 9596 5085 9600 5145
rect 9544 5079 9600 5085
rect 9315 5050 9385 5070
rect 9290 5010 9385 5050
rect 9445 5050 9515 5070
rect 9445 5010 9540 5050
rect 9290 4960 9540 5010
rect 9290 4920 9385 4960
rect 9315 4900 9385 4920
rect 9445 4920 9540 4960
rect 9445 4900 9515 4920
rect 9230 4885 9286 4891
rect 9230 4825 9234 4885
rect 9315 4875 9515 4900
rect 9570 4891 9600 5079
rect 9544 4885 9600 4891
rect 9286 4825 9544 4845
rect 9596 4825 9600 4885
rect 9230 4815 9600 4825
rect 9630 5145 10000 5155
rect 9630 5085 9634 5145
rect 9686 5125 9944 5145
rect 9630 5079 9686 5085
rect 9630 4891 9660 5079
rect 9715 5070 9915 5095
rect 9996 5085 10000 5145
rect 9944 5079 10000 5085
rect 9715 5050 9785 5070
rect 9690 5010 9785 5050
rect 9845 5050 9915 5070
rect 9845 5010 9940 5050
rect 9690 4960 9940 5010
rect 9690 4920 9785 4960
rect 9715 4900 9785 4920
rect 9845 4920 9940 4960
rect 9845 4900 9915 4920
rect 9630 4885 9686 4891
rect 9630 4825 9634 4885
rect 9715 4875 9915 4900
rect 9970 4891 10000 5079
rect 9944 4885 10000 4891
rect 9686 4825 9944 4845
rect 9996 4825 10000 4885
rect 9630 4815 10000 4825
rect 10030 5145 10400 5155
rect 10030 5085 10034 5145
rect 10086 5125 10344 5145
rect 10030 5079 10086 5085
rect 10030 4891 10060 5079
rect 10115 5070 10315 5095
rect 10396 5085 10400 5145
rect 10344 5079 10400 5085
rect 10115 5050 10185 5070
rect 10090 5010 10185 5050
rect 10245 5050 10315 5070
rect 10245 5010 10340 5050
rect 10090 4960 10340 5010
rect 10090 4920 10185 4960
rect 10115 4900 10185 4920
rect 10245 4920 10340 4960
rect 10245 4900 10315 4920
rect 10030 4885 10086 4891
rect 10030 4825 10034 4885
rect 10115 4875 10315 4900
rect 10370 4891 10400 5079
rect 10344 4885 10400 4891
rect 10086 4825 10344 4845
rect 10396 4825 10400 4885
rect 10030 4815 10400 4825
rect 10430 5145 10800 5155
rect 10430 5085 10434 5145
rect 10486 5125 10744 5145
rect 10430 5079 10486 5085
rect 10430 4891 10460 5079
rect 10515 5070 10715 5095
rect 10796 5085 10800 5145
rect 10744 5079 10800 5085
rect 10515 5050 10585 5070
rect 10490 5010 10585 5050
rect 10645 5050 10715 5070
rect 10645 5010 10740 5050
rect 10490 4960 10740 5010
rect 10490 4920 10585 4960
rect 10515 4900 10585 4920
rect 10645 4920 10740 4960
rect 10645 4900 10715 4920
rect 10430 4885 10486 4891
rect 10430 4825 10434 4885
rect 10515 4875 10715 4900
rect 10770 4891 10800 5079
rect 10744 4885 10800 4891
rect 10486 4825 10744 4845
rect 10796 4825 10800 4885
rect 10430 4815 10800 4825
rect 10830 5145 11200 5155
rect 10830 5085 10834 5145
rect 10886 5125 11144 5145
rect 10830 5079 10886 5085
rect 10830 4891 10860 5079
rect 10915 5070 11115 5095
rect 11196 5085 11200 5145
rect 11144 5079 11200 5085
rect 10915 5050 10985 5070
rect 10890 5010 10985 5050
rect 11045 5050 11115 5070
rect 11045 5010 11140 5050
rect 10890 4960 11140 5010
rect 10890 4920 10985 4960
rect 10915 4900 10985 4920
rect 11045 4920 11140 4960
rect 11045 4900 11115 4920
rect 10830 4885 10886 4891
rect 10830 4825 10834 4885
rect 10915 4875 11115 4900
rect 11170 4891 11200 5079
rect 11144 4885 11200 4891
rect 10886 4825 11144 4845
rect 11196 4825 11200 4885
rect 10830 4815 11200 4825
rect 11230 5145 11600 5155
rect 11230 5085 11234 5145
rect 11286 5125 11544 5145
rect 11230 5079 11286 5085
rect 11230 4891 11260 5079
rect 11315 5070 11515 5095
rect 11596 5085 11600 5145
rect 11544 5079 11600 5085
rect 11315 5050 11385 5070
rect 11290 5010 11385 5050
rect 11445 5050 11515 5070
rect 11445 5010 11540 5050
rect 11290 4960 11540 5010
rect 11290 4920 11385 4960
rect 11315 4900 11385 4920
rect 11445 4920 11540 4960
rect 11445 4900 11515 4920
rect 11230 4885 11286 4891
rect 11230 4825 11234 4885
rect 11315 4875 11515 4900
rect 11570 4891 11600 5079
rect 11544 4885 11600 4891
rect 11286 4825 11544 4845
rect 11596 4825 11600 4885
rect 11230 4815 11600 4825
rect 11630 5145 12000 5155
rect 11630 5085 11634 5145
rect 11686 5125 11944 5145
rect 11630 5079 11686 5085
rect 11630 4891 11660 5079
rect 11715 5070 11915 5095
rect 11996 5085 12000 5145
rect 11944 5079 12000 5085
rect 11715 5050 11785 5070
rect 11690 5010 11785 5050
rect 11845 5050 11915 5070
rect 11845 5010 11940 5050
rect 11690 4960 11940 5010
rect 11690 4920 11785 4960
rect 11715 4900 11785 4920
rect 11845 4920 11940 4960
rect 11845 4900 11915 4920
rect 11630 4885 11686 4891
rect 11630 4825 11634 4885
rect 11715 4875 11915 4900
rect 11970 4891 12000 5079
rect 11944 4885 12000 4891
rect 11686 4825 11944 4845
rect 11996 4825 12000 4885
rect 11630 4815 12000 4825
rect 12030 5145 12400 5155
rect 12030 5085 12034 5145
rect 12086 5125 12344 5145
rect 12030 5079 12086 5085
rect 12030 4891 12060 5079
rect 12115 5070 12315 5095
rect 12396 5085 12400 5145
rect 12344 5079 12400 5085
rect 12115 5050 12185 5070
rect 12090 5010 12185 5050
rect 12245 5050 12315 5070
rect 12245 5010 12340 5050
rect 12090 4960 12340 5010
rect 12090 4920 12185 4960
rect 12115 4900 12185 4920
rect 12245 4920 12340 4960
rect 12245 4900 12315 4920
rect 12030 4885 12086 4891
rect 12030 4825 12034 4885
rect 12115 4875 12315 4900
rect 12370 4891 12400 5079
rect 12344 4885 12400 4891
rect 12086 4825 12344 4845
rect 12396 4825 12400 4885
rect 12030 4815 12400 4825
rect 12430 5145 12800 5155
rect 12430 5085 12434 5145
rect 12486 5125 12744 5145
rect 12430 5079 12486 5085
rect 12430 4891 12460 5079
rect 12515 5070 12715 5095
rect 12796 5085 12800 5145
rect 12744 5079 12800 5085
rect 12515 5050 12585 5070
rect 12490 5010 12585 5050
rect 12645 5050 12715 5070
rect 12645 5010 12740 5050
rect 12490 4960 12740 5010
rect 12490 4920 12585 4960
rect 12515 4900 12585 4920
rect 12645 4920 12740 4960
rect 12645 4900 12715 4920
rect 12430 4885 12486 4891
rect 12430 4825 12434 4885
rect 12515 4875 12715 4900
rect 12770 4891 12800 5079
rect 12744 4885 12800 4891
rect 12486 4825 12744 4845
rect 12796 4825 12800 4885
rect 12430 4815 12800 4825
rect 12830 5145 13200 5155
rect 12830 5085 12834 5145
rect 12886 5125 13144 5145
rect 12830 5079 12886 5085
rect 12830 4891 12860 5079
rect 12915 5070 13115 5095
rect 13196 5085 13200 5145
rect 13144 5079 13200 5085
rect 12915 5050 12985 5070
rect 12890 5010 12985 5050
rect 13045 5050 13115 5070
rect 13045 5010 13140 5050
rect 12890 4960 13140 5010
rect 12890 4920 12985 4960
rect 12915 4900 12985 4920
rect 13045 4920 13140 4960
rect 13045 4900 13115 4920
rect 12830 4885 12886 4891
rect 12830 4825 12834 4885
rect 12915 4875 13115 4900
rect 13170 4891 13200 5079
rect 13144 4885 13200 4891
rect 12886 4825 13144 4845
rect 13196 4825 13200 4885
rect 12830 4815 13200 4825
rect -370 4775 0 4785
rect -370 4715 -366 4775
rect -314 4755 -56 4775
rect -370 4709 -314 4715
rect -370 4521 -340 4709
rect -285 4700 -85 4725
rect -4 4715 0 4775
rect -56 4709 0 4715
rect -285 4680 -215 4700
rect -310 4640 -215 4680
rect -155 4680 -85 4700
rect -155 4640 -60 4680
rect -310 4590 -60 4640
rect -310 4550 -215 4590
rect -285 4530 -215 4550
rect -155 4550 -60 4590
rect -155 4530 -85 4550
rect -370 4515 -314 4521
rect -370 4455 -366 4515
rect -285 4505 -85 4530
rect -30 4521 0 4709
rect -56 4515 0 4521
rect -314 4455 -56 4475
rect -4 4455 0 4515
rect -370 4445 0 4455
rect 30 4775 400 4785
rect 30 4715 34 4775
rect 86 4755 344 4775
rect 30 4709 86 4715
rect 30 4521 60 4709
rect 115 4700 315 4725
rect 396 4715 400 4775
rect 344 4709 400 4715
rect 115 4680 185 4700
rect 90 4640 185 4680
rect 245 4680 315 4700
rect 245 4640 340 4680
rect 90 4590 340 4640
rect 90 4550 185 4590
rect 115 4530 185 4550
rect 245 4550 340 4590
rect 245 4530 315 4550
rect 30 4515 86 4521
rect 30 4455 34 4515
rect 115 4505 315 4530
rect 370 4521 400 4709
rect 344 4515 400 4521
rect 86 4455 344 4475
rect 396 4455 400 4515
rect 30 4445 400 4455
rect 430 4775 800 4785
rect 430 4715 434 4775
rect 486 4755 744 4775
rect 430 4709 486 4715
rect 430 4521 460 4709
rect 515 4700 715 4725
rect 796 4715 800 4775
rect 744 4709 800 4715
rect 515 4680 585 4700
rect 490 4640 585 4680
rect 645 4680 715 4700
rect 645 4640 740 4680
rect 490 4590 740 4640
rect 490 4550 585 4590
rect 515 4530 585 4550
rect 645 4550 740 4590
rect 645 4530 715 4550
rect 430 4515 486 4521
rect 430 4455 434 4515
rect 515 4505 715 4530
rect 770 4521 800 4709
rect 744 4515 800 4521
rect 486 4455 744 4475
rect 796 4455 800 4515
rect 430 4445 800 4455
rect 830 4775 1200 4785
rect 830 4715 834 4775
rect 886 4755 1144 4775
rect 830 4709 886 4715
rect 830 4521 860 4709
rect 915 4700 1115 4725
rect 1196 4715 1200 4775
rect 1144 4709 1200 4715
rect 915 4680 985 4700
rect 890 4640 985 4680
rect 1045 4680 1115 4700
rect 1045 4640 1140 4680
rect 890 4590 1140 4640
rect 890 4550 985 4590
rect 915 4530 985 4550
rect 1045 4550 1140 4590
rect 1045 4530 1115 4550
rect 830 4515 886 4521
rect 830 4455 834 4515
rect 915 4505 1115 4530
rect 1170 4521 1200 4709
rect 1144 4515 1200 4521
rect 886 4455 1144 4475
rect 1196 4455 1200 4515
rect 830 4445 1200 4455
rect 1230 4775 1600 4785
rect 1230 4715 1234 4775
rect 1286 4755 1544 4775
rect 1230 4709 1286 4715
rect 1230 4521 1260 4709
rect 1315 4700 1515 4725
rect 1596 4715 1600 4775
rect 1544 4709 1600 4715
rect 1315 4680 1385 4700
rect 1290 4640 1385 4680
rect 1445 4680 1515 4700
rect 1445 4640 1540 4680
rect 1290 4590 1540 4640
rect 1290 4550 1385 4590
rect 1315 4530 1385 4550
rect 1445 4550 1540 4590
rect 1445 4530 1515 4550
rect 1230 4515 1286 4521
rect 1230 4455 1234 4515
rect 1315 4505 1515 4530
rect 1570 4521 1600 4709
rect 1544 4515 1600 4521
rect 1286 4455 1544 4475
rect 1596 4455 1600 4515
rect 1230 4445 1600 4455
rect 1630 4775 2000 4785
rect 1630 4715 1634 4775
rect 1686 4755 1944 4775
rect 1630 4709 1686 4715
rect 1630 4521 1660 4709
rect 1715 4700 1915 4725
rect 1996 4715 2000 4775
rect 1944 4709 2000 4715
rect 1715 4680 1785 4700
rect 1690 4640 1785 4680
rect 1845 4680 1915 4700
rect 1845 4640 1940 4680
rect 1690 4590 1940 4640
rect 1690 4550 1785 4590
rect 1715 4530 1785 4550
rect 1845 4550 1940 4590
rect 1845 4530 1915 4550
rect 1630 4515 1686 4521
rect 1630 4455 1634 4515
rect 1715 4505 1915 4530
rect 1970 4521 2000 4709
rect 1944 4515 2000 4521
rect 1686 4455 1944 4475
rect 1996 4455 2000 4515
rect 1630 4445 2000 4455
rect 2030 4775 2400 4785
rect 2030 4715 2034 4775
rect 2086 4755 2344 4775
rect 2030 4709 2086 4715
rect 2030 4521 2060 4709
rect 2115 4700 2315 4725
rect 2396 4715 2400 4775
rect 2344 4709 2400 4715
rect 2115 4680 2185 4700
rect 2090 4640 2185 4680
rect 2245 4680 2315 4700
rect 2245 4640 2340 4680
rect 2090 4590 2340 4640
rect 2090 4550 2185 4590
rect 2115 4530 2185 4550
rect 2245 4550 2340 4590
rect 2245 4530 2315 4550
rect 2030 4515 2086 4521
rect 2030 4455 2034 4515
rect 2115 4505 2315 4530
rect 2370 4521 2400 4709
rect 2344 4515 2400 4521
rect 2086 4455 2344 4475
rect 2396 4455 2400 4515
rect 2030 4445 2400 4455
rect 2430 4775 2800 4785
rect 2430 4715 2434 4775
rect 2486 4755 2744 4775
rect 2430 4709 2486 4715
rect 2430 4521 2460 4709
rect 2515 4700 2715 4725
rect 2796 4715 2800 4775
rect 2744 4709 2800 4715
rect 2515 4680 2585 4700
rect 2490 4640 2585 4680
rect 2645 4680 2715 4700
rect 2645 4640 2740 4680
rect 2490 4590 2740 4640
rect 2490 4550 2585 4590
rect 2515 4530 2585 4550
rect 2645 4550 2740 4590
rect 2645 4530 2715 4550
rect 2430 4515 2486 4521
rect 2430 4455 2434 4515
rect 2515 4505 2715 4530
rect 2770 4521 2800 4709
rect 2744 4515 2800 4521
rect 2486 4455 2744 4475
rect 2796 4455 2800 4515
rect 2430 4445 2800 4455
rect 2830 4775 3200 4785
rect 2830 4715 2834 4775
rect 2886 4755 3144 4775
rect 2830 4709 2886 4715
rect 2830 4521 2860 4709
rect 2915 4700 3115 4725
rect 3196 4715 3200 4775
rect 3144 4709 3200 4715
rect 2915 4680 2985 4700
rect 2890 4640 2985 4680
rect 3045 4680 3115 4700
rect 3045 4640 3140 4680
rect 2890 4590 3140 4640
rect 2890 4550 2985 4590
rect 2915 4530 2985 4550
rect 3045 4550 3140 4590
rect 3045 4530 3115 4550
rect 2830 4515 2886 4521
rect 2830 4455 2834 4515
rect 2915 4505 3115 4530
rect 3170 4521 3200 4709
rect 3144 4515 3200 4521
rect 2886 4455 3144 4475
rect 3196 4455 3200 4515
rect 2830 4445 3200 4455
rect 3230 4775 3600 4785
rect 3230 4715 3234 4775
rect 3286 4755 3544 4775
rect 3230 4709 3286 4715
rect 3230 4521 3260 4709
rect 3315 4700 3515 4725
rect 3596 4715 3600 4775
rect 3544 4709 3600 4715
rect 3315 4680 3385 4700
rect 3290 4640 3385 4680
rect 3445 4680 3515 4700
rect 3445 4640 3540 4680
rect 3290 4590 3540 4640
rect 3290 4550 3385 4590
rect 3315 4530 3385 4550
rect 3445 4550 3540 4590
rect 3445 4530 3515 4550
rect 3230 4515 3286 4521
rect 3230 4455 3234 4515
rect 3315 4505 3515 4530
rect 3570 4521 3600 4709
rect 3544 4515 3600 4521
rect 3286 4455 3544 4475
rect 3596 4455 3600 4515
rect 3230 4445 3600 4455
rect 3630 4775 4000 4785
rect 3630 4715 3634 4775
rect 3686 4755 3944 4775
rect 3630 4709 3686 4715
rect 3630 4521 3660 4709
rect 3715 4700 3915 4725
rect 3996 4715 4000 4775
rect 3944 4709 4000 4715
rect 3715 4680 3785 4700
rect 3690 4640 3785 4680
rect 3845 4680 3915 4700
rect 3845 4640 3940 4680
rect 3690 4590 3940 4640
rect 3690 4550 3785 4590
rect 3715 4530 3785 4550
rect 3845 4550 3940 4590
rect 3845 4530 3915 4550
rect 3630 4515 3686 4521
rect 3630 4455 3634 4515
rect 3715 4505 3915 4530
rect 3970 4521 4000 4709
rect 3944 4515 4000 4521
rect 3686 4455 3944 4475
rect 3996 4455 4000 4515
rect 3630 4445 4000 4455
rect 4030 4775 4400 4785
rect 4030 4715 4034 4775
rect 4086 4755 4344 4775
rect 4030 4709 4086 4715
rect 4030 4521 4060 4709
rect 4115 4700 4315 4725
rect 4396 4715 4400 4775
rect 4344 4709 4400 4715
rect 4115 4680 4185 4700
rect 4090 4640 4185 4680
rect 4245 4680 4315 4700
rect 4245 4640 4340 4680
rect 4090 4590 4340 4640
rect 4090 4550 4185 4590
rect 4115 4530 4185 4550
rect 4245 4550 4340 4590
rect 4245 4530 4315 4550
rect 4030 4515 4086 4521
rect 4030 4455 4034 4515
rect 4115 4505 4315 4530
rect 4370 4521 4400 4709
rect 4344 4515 4400 4521
rect 4086 4455 4344 4475
rect 4396 4455 4400 4515
rect 4030 4445 4400 4455
rect 4430 4775 4800 4785
rect 4430 4715 4434 4775
rect 4486 4755 4744 4775
rect 4430 4709 4486 4715
rect 4430 4521 4460 4709
rect 4515 4700 4715 4725
rect 4796 4715 4800 4775
rect 4744 4709 4800 4715
rect 4515 4680 4585 4700
rect 4490 4640 4585 4680
rect 4645 4680 4715 4700
rect 4645 4640 4740 4680
rect 4490 4590 4740 4640
rect 4490 4550 4585 4590
rect 4515 4530 4585 4550
rect 4645 4550 4740 4590
rect 4645 4530 4715 4550
rect 4430 4515 4486 4521
rect 4430 4455 4434 4515
rect 4515 4505 4715 4530
rect 4770 4521 4800 4709
rect 4744 4515 4800 4521
rect 4486 4455 4744 4475
rect 4796 4455 4800 4515
rect 4430 4445 4800 4455
rect 4830 4775 5200 4785
rect 4830 4715 4834 4775
rect 4886 4755 5144 4775
rect 4830 4709 4886 4715
rect 4830 4521 4860 4709
rect 4915 4700 5115 4725
rect 5196 4715 5200 4775
rect 5144 4709 5200 4715
rect 4915 4680 4985 4700
rect 4890 4640 4985 4680
rect 5045 4680 5115 4700
rect 5045 4640 5140 4680
rect 4890 4590 5140 4640
rect 4890 4550 4985 4590
rect 4915 4530 4985 4550
rect 5045 4550 5140 4590
rect 5045 4530 5115 4550
rect 4830 4515 4886 4521
rect 4830 4455 4834 4515
rect 4915 4505 5115 4530
rect 5170 4521 5200 4709
rect 5144 4515 5200 4521
rect 4886 4455 5144 4475
rect 5196 4455 5200 4515
rect 4830 4445 5200 4455
rect 5230 4775 5600 4785
rect 5230 4715 5234 4775
rect 5286 4755 5544 4775
rect 5230 4709 5286 4715
rect 5230 4521 5260 4709
rect 5315 4700 5515 4725
rect 5596 4715 5600 4775
rect 5544 4709 5600 4715
rect 5315 4680 5385 4700
rect 5290 4640 5385 4680
rect 5445 4680 5515 4700
rect 5445 4640 5540 4680
rect 5290 4590 5540 4640
rect 5290 4550 5385 4590
rect 5315 4530 5385 4550
rect 5445 4550 5540 4590
rect 5445 4530 5515 4550
rect 5230 4515 5286 4521
rect 5230 4455 5234 4515
rect 5315 4505 5515 4530
rect 5570 4521 5600 4709
rect 5544 4515 5600 4521
rect 5286 4455 5544 4475
rect 5596 4455 5600 4515
rect 5230 4445 5600 4455
rect 5630 4775 6000 4785
rect 5630 4715 5634 4775
rect 5686 4755 5944 4775
rect 5630 4709 5686 4715
rect 5630 4521 5660 4709
rect 5715 4700 5915 4725
rect 5996 4715 6000 4775
rect 5944 4709 6000 4715
rect 5715 4680 5785 4700
rect 5690 4640 5785 4680
rect 5845 4680 5915 4700
rect 5845 4640 5940 4680
rect 5690 4590 5940 4640
rect 5690 4550 5785 4590
rect 5715 4530 5785 4550
rect 5845 4550 5940 4590
rect 5845 4530 5915 4550
rect 5630 4515 5686 4521
rect 5630 4455 5634 4515
rect 5715 4505 5915 4530
rect 5970 4521 6000 4709
rect 5944 4515 6000 4521
rect 5686 4455 5944 4475
rect 5996 4455 6000 4515
rect 5630 4445 6000 4455
rect 6030 4775 6400 4785
rect 6030 4715 6034 4775
rect 6086 4755 6344 4775
rect 6030 4709 6086 4715
rect 6030 4521 6060 4709
rect 6115 4700 6315 4725
rect 6396 4715 6400 4775
rect 6344 4709 6400 4715
rect 6115 4680 6185 4700
rect 6090 4640 6185 4680
rect 6245 4680 6315 4700
rect 6245 4640 6340 4680
rect 6090 4590 6340 4640
rect 6090 4550 6185 4590
rect 6115 4530 6185 4550
rect 6245 4550 6340 4590
rect 6245 4530 6315 4550
rect 6030 4515 6086 4521
rect 6030 4455 6034 4515
rect 6115 4505 6315 4530
rect 6370 4521 6400 4709
rect 6344 4515 6400 4521
rect 6086 4455 6344 4475
rect 6396 4455 6400 4515
rect 6030 4445 6400 4455
rect 6430 4775 6800 4785
rect 6430 4715 6434 4775
rect 6486 4755 6744 4775
rect 6430 4709 6486 4715
rect 6430 4521 6460 4709
rect 6515 4700 6715 4725
rect 6796 4715 6800 4775
rect 6744 4709 6800 4715
rect 6515 4680 6585 4700
rect 6490 4640 6585 4680
rect 6645 4680 6715 4700
rect 6645 4640 6740 4680
rect 6490 4590 6740 4640
rect 6490 4550 6585 4590
rect 6515 4530 6585 4550
rect 6645 4550 6740 4590
rect 6645 4530 6715 4550
rect 6430 4515 6486 4521
rect 6430 4455 6434 4515
rect 6515 4505 6715 4530
rect 6770 4521 6800 4709
rect 6744 4515 6800 4521
rect 6486 4455 6744 4475
rect 6796 4455 6800 4515
rect 6430 4445 6800 4455
rect 6830 4775 7200 4785
rect 6830 4715 6834 4775
rect 6886 4755 7144 4775
rect 6830 4709 6886 4715
rect 6830 4521 6860 4709
rect 6915 4700 7115 4725
rect 7196 4715 7200 4775
rect 7144 4709 7200 4715
rect 6915 4680 6985 4700
rect 6890 4640 6985 4680
rect 7045 4680 7115 4700
rect 7045 4640 7140 4680
rect 6890 4590 7140 4640
rect 6890 4550 6985 4590
rect 6915 4530 6985 4550
rect 7045 4550 7140 4590
rect 7045 4530 7115 4550
rect 6830 4515 6886 4521
rect 6830 4455 6834 4515
rect 6915 4505 7115 4530
rect 7170 4521 7200 4709
rect 7144 4515 7200 4521
rect 6886 4455 7144 4475
rect 7196 4455 7200 4515
rect 6830 4445 7200 4455
rect 7230 4775 7600 4785
rect 7230 4715 7234 4775
rect 7286 4755 7544 4775
rect 7230 4709 7286 4715
rect 7230 4521 7260 4709
rect 7315 4700 7515 4725
rect 7596 4715 7600 4775
rect 7544 4709 7600 4715
rect 7315 4680 7385 4700
rect 7290 4640 7385 4680
rect 7445 4680 7515 4700
rect 7445 4640 7540 4680
rect 7290 4590 7540 4640
rect 7290 4550 7385 4590
rect 7315 4530 7385 4550
rect 7445 4550 7540 4590
rect 7445 4530 7515 4550
rect 7230 4515 7286 4521
rect 7230 4455 7234 4515
rect 7315 4505 7515 4530
rect 7570 4521 7600 4709
rect 7544 4515 7600 4521
rect 7286 4455 7544 4475
rect 7596 4455 7600 4515
rect 7230 4445 7600 4455
rect 7630 4775 8000 4785
rect 7630 4715 7634 4775
rect 7686 4755 7944 4775
rect 7630 4709 7686 4715
rect 7630 4521 7660 4709
rect 7715 4700 7915 4725
rect 7996 4715 8000 4775
rect 7944 4709 8000 4715
rect 7715 4680 7785 4700
rect 7690 4640 7785 4680
rect 7845 4680 7915 4700
rect 7845 4640 7940 4680
rect 7690 4590 7940 4640
rect 7690 4550 7785 4590
rect 7715 4530 7785 4550
rect 7845 4550 7940 4590
rect 7845 4530 7915 4550
rect 7630 4515 7686 4521
rect 7630 4455 7634 4515
rect 7715 4505 7915 4530
rect 7970 4521 8000 4709
rect 7944 4515 8000 4521
rect 7686 4455 7944 4475
rect 7996 4455 8000 4515
rect 7630 4445 8000 4455
rect 8030 4775 8400 4785
rect 8030 4715 8034 4775
rect 8086 4755 8344 4775
rect 8030 4709 8086 4715
rect 8030 4521 8060 4709
rect 8115 4700 8315 4725
rect 8396 4715 8400 4775
rect 8344 4709 8400 4715
rect 8115 4680 8185 4700
rect 8090 4640 8185 4680
rect 8245 4680 8315 4700
rect 8245 4640 8340 4680
rect 8090 4590 8340 4640
rect 8090 4550 8185 4590
rect 8115 4530 8185 4550
rect 8245 4550 8340 4590
rect 8245 4530 8315 4550
rect 8030 4515 8086 4521
rect 8030 4455 8034 4515
rect 8115 4505 8315 4530
rect 8370 4521 8400 4709
rect 8344 4515 8400 4521
rect 8086 4455 8344 4475
rect 8396 4455 8400 4515
rect 8030 4445 8400 4455
rect 8430 4775 8800 4785
rect 8430 4715 8434 4775
rect 8486 4755 8744 4775
rect 8430 4709 8486 4715
rect 8430 4521 8460 4709
rect 8515 4700 8715 4725
rect 8796 4715 8800 4775
rect 8744 4709 8800 4715
rect 8515 4680 8585 4700
rect 8490 4640 8585 4680
rect 8645 4680 8715 4700
rect 8645 4640 8740 4680
rect 8490 4590 8740 4640
rect 8490 4550 8585 4590
rect 8515 4530 8585 4550
rect 8645 4550 8740 4590
rect 8645 4530 8715 4550
rect 8430 4515 8486 4521
rect 8430 4455 8434 4515
rect 8515 4505 8715 4530
rect 8770 4521 8800 4709
rect 8744 4515 8800 4521
rect 8486 4455 8744 4475
rect 8796 4455 8800 4515
rect 8430 4445 8800 4455
rect 8830 4775 9200 4785
rect 8830 4715 8834 4775
rect 8886 4755 9144 4775
rect 8830 4709 8886 4715
rect 8830 4521 8860 4709
rect 8915 4700 9115 4725
rect 9196 4715 9200 4775
rect 9144 4709 9200 4715
rect 8915 4680 8985 4700
rect 8890 4640 8985 4680
rect 9045 4680 9115 4700
rect 9045 4640 9140 4680
rect 8890 4590 9140 4640
rect 8890 4550 8985 4590
rect 8915 4530 8985 4550
rect 9045 4550 9140 4590
rect 9045 4530 9115 4550
rect 8830 4515 8886 4521
rect 8830 4455 8834 4515
rect 8915 4505 9115 4530
rect 9170 4521 9200 4709
rect 9144 4515 9200 4521
rect 8886 4455 9144 4475
rect 9196 4455 9200 4515
rect 8830 4445 9200 4455
rect 9230 4775 9600 4785
rect 9230 4715 9234 4775
rect 9286 4755 9544 4775
rect 9230 4709 9286 4715
rect 9230 4521 9260 4709
rect 9315 4700 9515 4725
rect 9596 4715 9600 4775
rect 9544 4709 9600 4715
rect 9315 4680 9385 4700
rect 9290 4640 9385 4680
rect 9445 4680 9515 4700
rect 9445 4640 9540 4680
rect 9290 4590 9540 4640
rect 9290 4550 9385 4590
rect 9315 4530 9385 4550
rect 9445 4550 9540 4590
rect 9445 4530 9515 4550
rect 9230 4515 9286 4521
rect 9230 4455 9234 4515
rect 9315 4505 9515 4530
rect 9570 4521 9600 4709
rect 9544 4515 9600 4521
rect 9286 4455 9544 4475
rect 9596 4455 9600 4515
rect 9230 4445 9600 4455
rect 9630 4775 10000 4785
rect 9630 4715 9634 4775
rect 9686 4755 9944 4775
rect 9630 4709 9686 4715
rect 9630 4521 9660 4709
rect 9715 4700 9915 4725
rect 9996 4715 10000 4775
rect 9944 4709 10000 4715
rect 9715 4680 9785 4700
rect 9690 4640 9785 4680
rect 9845 4680 9915 4700
rect 9845 4640 9940 4680
rect 9690 4590 9940 4640
rect 9690 4550 9785 4590
rect 9715 4530 9785 4550
rect 9845 4550 9940 4590
rect 9845 4530 9915 4550
rect 9630 4515 9686 4521
rect 9630 4455 9634 4515
rect 9715 4505 9915 4530
rect 9970 4521 10000 4709
rect 9944 4515 10000 4521
rect 9686 4455 9944 4475
rect 9996 4455 10000 4515
rect 9630 4445 10000 4455
rect 10030 4775 10400 4785
rect 10030 4715 10034 4775
rect 10086 4755 10344 4775
rect 10030 4709 10086 4715
rect 10030 4521 10060 4709
rect 10115 4700 10315 4725
rect 10396 4715 10400 4775
rect 10344 4709 10400 4715
rect 10115 4680 10185 4700
rect 10090 4640 10185 4680
rect 10245 4680 10315 4700
rect 10245 4640 10340 4680
rect 10090 4590 10340 4640
rect 10090 4550 10185 4590
rect 10115 4530 10185 4550
rect 10245 4550 10340 4590
rect 10245 4530 10315 4550
rect 10030 4515 10086 4521
rect 10030 4455 10034 4515
rect 10115 4505 10315 4530
rect 10370 4521 10400 4709
rect 10344 4515 10400 4521
rect 10086 4455 10344 4475
rect 10396 4455 10400 4515
rect 10030 4445 10400 4455
rect 10430 4775 10800 4785
rect 10430 4715 10434 4775
rect 10486 4755 10744 4775
rect 10430 4709 10486 4715
rect 10430 4521 10460 4709
rect 10515 4700 10715 4725
rect 10796 4715 10800 4775
rect 10744 4709 10800 4715
rect 10515 4680 10585 4700
rect 10490 4640 10585 4680
rect 10645 4680 10715 4700
rect 10645 4640 10740 4680
rect 10490 4590 10740 4640
rect 10490 4550 10585 4590
rect 10515 4530 10585 4550
rect 10645 4550 10740 4590
rect 10645 4530 10715 4550
rect 10430 4515 10486 4521
rect 10430 4455 10434 4515
rect 10515 4505 10715 4530
rect 10770 4521 10800 4709
rect 10744 4515 10800 4521
rect 10486 4455 10744 4475
rect 10796 4455 10800 4515
rect 10430 4445 10800 4455
rect 10830 4775 11200 4785
rect 10830 4715 10834 4775
rect 10886 4755 11144 4775
rect 10830 4709 10886 4715
rect 10830 4521 10860 4709
rect 10915 4700 11115 4725
rect 11196 4715 11200 4775
rect 11144 4709 11200 4715
rect 10915 4680 10985 4700
rect 10890 4640 10985 4680
rect 11045 4680 11115 4700
rect 11045 4640 11140 4680
rect 10890 4590 11140 4640
rect 10890 4550 10985 4590
rect 10915 4530 10985 4550
rect 11045 4550 11140 4590
rect 11045 4530 11115 4550
rect 10830 4515 10886 4521
rect 10830 4455 10834 4515
rect 10915 4505 11115 4530
rect 11170 4521 11200 4709
rect 11144 4515 11200 4521
rect 10886 4455 11144 4475
rect 11196 4455 11200 4515
rect 10830 4445 11200 4455
rect 11230 4775 11600 4785
rect 11230 4715 11234 4775
rect 11286 4755 11544 4775
rect 11230 4709 11286 4715
rect 11230 4521 11260 4709
rect 11315 4700 11515 4725
rect 11596 4715 11600 4775
rect 11544 4709 11600 4715
rect 11315 4680 11385 4700
rect 11290 4640 11385 4680
rect 11445 4680 11515 4700
rect 11445 4640 11540 4680
rect 11290 4590 11540 4640
rect 11290 4550 11385 4590
rect 11315 4530 11385 4550
rect 11445 4550 11540 4590
rect 11445 4530 11515 4550
rect 11230 4515 11286 4521
rect 11230 4455 11234 4515
rect 11315 4505 11515 4530
rect 11570 4521 11600 4709
rect 11544 4515 11600 4521
rect 11286 4455 11544 4475
rect 11596 4455 11600 4515
rect 11230 4445 11600 4455
rect 11630 4775 12000 4785
rect 11630 4715 11634 4775
rect 11686 4755 11944 4775
rect 11630 4709 11686 4715
rect 11630 4521 11660 4709
rect 11715 4700 11915 4725
rect 11996 4715 12000 4775
rect 11944 4709 12000 4715
rect 11715 4680 11785 4700
rect 11690 4640 11785 4680
rect 11845 4680 11915 4700
rect 11845 4640 11940 4680
rect 11690 4590 11940 4640
rect 11690 4550 11785 4590
rect 11715 4530 11785 4550
rect 11845 4550 11940 4590
rect 11845 4530 11915 4550
rect 11630 4515 11686 4521
rect 11630 4455 11634 4515
rect 11715 4505 11915 4530
rect 11970 4521 12000 4709
rect 11944 4515 12000 4521
rect 11686 4455 11944 4475
rect 11996 4455 12000 4515
rect 11630 4445 12000 4455
rect 12030 4775 12400 4785
rect 12030 4715 12034 4775
rect 12086 4755 12344 4775
rect 12030 4709 12086 4715
rect 12030 4521 12060 4709
rect 12115 4700 12315 4725
rect 12396 4715 12400 4775
rect 12344 4709 12400 4715
rect 12115 4680 12185 4700
rect 12090 4640 12185 4680
rect 12245 4680 12315 4700
rect 12245 4640 12340 4680
rect 12090 4590 12340 4640
rect 12090 4550 12185 4590
rect 12115 4530 12185 4550
rect 12245 4550 12340 4590
rect 12245 4530 12315 4550
rect 12030 4515 12086 4521
rect 12030 4455 12034 4515
rect 12115 4505 12315 4530
rect 12370 4521 12400 4709
rect 12344 4515 12400 4521
rect 12086 4455 12344 4475
rect 12396 4455 12400 4515
rect 12030 4445 12400 4455
rect 12430 4775 12800 4785
rect 12430 4715 12434 4775
rect 12486 4755 12744 4775
rect 12430 4709 12486 4715
rect 12430 4521 12460 4709
rect 12515 4700 12715 4725
rect 12796 4715 12800 4775
rect 12744 4709 12800 4715
rect 12515 4680 12585 4700
rect 12490 4640 12585 4680
rect 12645 4680 12715 4700
rect 12645 4640 12740 4680
rect 12490 4590 12740 4640
rect 12490 4550 12585 4590
rect 12515 4530 12585 4550
rect 12645 4550 12740 4590
rect 12645 4530 12715 4550
rect 12430 4515 12486 4521
rect 12430 4455 12434 4515
rect 12515 4505 12715 4530
rect 12770 4521 12800 4709
rect 12744 4515 12800 4521
rect 12486 4455 12744 4475
rect 12796 4455 12800 4515
rect 12430 4445 12800 4455
rect 12830 4775 13200 4785
rect 12830 4715 12834 4775
rect 12886 4755 13144 4775
rect 12830 4709 12886 4715
rect 12830 4521 12860 4709
rect 12915 4700 13115 4725
rect 13196 4715 13200 4775
rect 13144 4709 13200 4715
rect 12915 4680 12985 4700
rect 12890 4640 12985 4680
rect 13045 4680 13115 4700
rect 13045 4640 13140 4680
rect 12890 4590 13140 4640
rect 12890 4550 12985 4590
rect 12915 4530 12985 4550
rect 13045 4550 13140 4590
rect 13045 4530 13115 4550
rect 12830 4515 12886 4521
rect 12830 4455 12834 4515
rect 12915 4505 13115 4530
rect 13170 4521 13200 4709
rect 13144 4515 13200 4521
rect 12886 4455 13144 4475
rect 13196 4455 13200 4515
rect 12830 4445 13200 4455
rect -370 4405 0 4415
rect -370 4345 -366 4405
rect -314 4385 -56 4405
rect -370 4339 -314 4345
rect -370 4151 -340 4339
rect -285 4330 -85 4355
rect -4 4345 0 4405
rect -56 4339 0 4345
rect -285 4310 -215 4330
rect -310 4270 -215 4310
rect -155 4310 -85 4330
rect -155 4270 -60 4310
rect -310 4220 -60 4270
rect -310 4180 -215 4220
rect -285 4160 -215 4180
rect -155 4180 -60 4220
rect -155 4160 -85 4180
rect -370 4145 -314 4151
rect -370 4085 -366 4145
rect -285 4135 -85 4160
rect -30 4151 0 4339
rect -56 4145 0 4151
rect -314 4085 -56 4105
rect -4 4085 0 4145
rect -370 4075 0 4085
rect 30 4405 400 4415
rect 30 4345 34 4405
rect 86 4385 344 4405
rect 30 4339 86 4345
rect 30 4151 60 4339
rect 115 4330 315 4355
rect 396 4345 400 4405
rect 344 4339 400 4345
rect 115 4310 185 4330
rect 90 4270 185 4310
rect 245 4310 315 4330
rect 245 4270 340 4310
rect 90 4220 340 4270
rect 90 4180 185 4220
rect 115 4160 185 4180
rect 245 4180 340 4220
rect 245 4160 315 4180
rect 30 4145 86 4151
rect 30 4085 34 4145
rect 115 4135 315 4160
rect 370 4151 400 4339
rect 344 4145 400 4151
rect 86 4085 344 4105
rect 396 4085 400 4145
rect 30 4075 400 4085
rect 430 4405 800 4415
rect 430 4345 434 4405
rect 486 4385 744 4405
rect 430 4339 486 4345
rect 430 4151 460 4339
rect 515 4330 715 4355
rect 796 4345 800 4405
rect 744 4339 800 4345
rect 515 4310 585 4330
rect 490 4270 585 4310
rect 645 4310 715 4330
rect 645 4270 740 4310
rect 490 4220 740 4270
rect 490 4180 585 4220
rect 515 4160 585 4180
rect 645 4180 740 4220
rect 645 4160 715 4180
rect 430 4145 486 4151
rect 430 4085 434 4145
rect 515 4135 715 4160
rect 770 4151 800 4339
rect 744 4145 800 4151
rect 486 4085 744 4105
rect 796 4085 800 4145
rect 430 4075 800 4085
rect 830 4405 1200 4415
rect 830 4345 834 4405
rect 886 4385 1144 4405
rect 830 4339 886 4345
rect 830 4151 860 4339
rect 915 4330 1115 4355
rect 1196 4345 1200 4405
rect 1144 4339 1200 4345
rect 915 4310 985 4330
rect 890 4270 985 4310
rect 1045 4310 1115 4330
rect 1045 4270 1140 4310
rect 890 4220 1140 4270
rect 890 4180 985 4220
rect 915 4160 985 4180
rect 1045 4180 1140 4220
rect 1045 4160 1115 4180
rect 830 4145 886 4151
rect 830 4085 834 4145
rect 915 4135 1115 4160
rect 1170 4151 1200 4339
rect 1144 4145 1200 4151
rect 886 4085 1144 4105
rect 1196 4085 1200 4145
rect 830 4075 1200 4085
rect 1230 4405 1600 4415
rect 1230 4345 1234 4405
rect 1286 4385 1544 4405
rect 1230 4339 1286 4345
rect 1230 4151 1260 4339
rect 1315 4330 1515 4355
rect 1596 4345 1600 4405
rect 1544 4339 1600 4345
rect 1315 4310 1385 4330
rect 1290 4270 1385 4310
rect 1445 4310 1515 4330
rect 1445 4270 1540 4310
rect 1290 4220 1540 4270
rect 1290 4180 1385 4220
rect 1315 4160 1385 4180
rect 1445 4180 1540 4220
rect 1445 4160 1515 4180
rect 1230 4145 1286 4151
rect 1230 4085 1234 4145
rect 1315 4135 1515 4160
rect 1570 4151 1600 4339
rect 1544 4145 1600 4151
rect 1286 4085 1544 4105
rect 1596 4085 1600 4145
rect 1230 4075 1600 4085
rect 1630 4405 2000 4415
rect 1630 4345 1634 4405
rect 1686 4385 1944 4405
rect 1630 4339 1686 4345
rect 1630 4151 1660 4339
rect 1715 4330 1915 4355
rect 1996 4345 2000 4405
rect 1944 4339 2000 4345
rect 1715 4310 1785 4330
rect 1690 4270 1785 4310
rect 1845 4310 1915 4330
rect 1845 4270 1940 4310
rect 1690 4220 1940 4270
rect 1690 4180 1785 4220
rect 1715 4160 1785 4180
rect 1845 4180 1940 4220
rect 1845 4160 1915 4180
rect 1630 4145 1686 4151
rect 1630 4085 1634 4145
rect 1715 4135 1915 4160
rect 1970 4151 2000 4339
rect 1944 4145 2000 4151
rect 1686 4085 1944 4105
rect 1996 4085 2000 4145
rect 1630 4075 2000 4085
rect 2030 4405 2400 4415
rect 2030 4345 2034 4405
rect 2086 4385 2344 4405
rect 2030 4339 2086 4345
rect 2030 4151 2060 4339
rect 2115 4330 2315 4355
rect 2396 4345 2400 4405
rect 2344 4339 2400 4345
rect 2115 4310 2185 4330
rect 2090 4270 2185 4310
rect 2245 4310 2315 4330
rect 2245 4270 2340 4310
rect 2090 4220 2340 4270
rect 2090 4180 2185 4220
rect 2115 4160 2185 4180
rect 2245 4180 2340 4220
rect 2245 4160 2315 4180
rect 2030 4145 2086 4151
rect 2030 4085 2034 4145
rect 2115 4135 2315 4160
rect 2370 4151 2400 4339
rect 2344 4145 2400 4151
rect 2086 4085 2344 4105
rect 2396 4085 2400 4145
rect 2030 4075 2400 4085
rect 2430 4405 2800 4415
rect 2430 4345 2434 4405
rect 2486 4385 2744 4405
rect 2430 4339 2486 4345
rect 2430 4151 2460 4339
rect 2515 4330 2715 4355
rect 2796 4345 2800 4405
rect 2744 4339 2800 4345
rect 2515 4310 2585 4330
rect 2490 4270 2585 4310
rect 2645 4310 2715 4330
rect 2645 4270 2740 4310
rect 2490 4220 2740 4270
rect 2490 4180 2585 4220
rect 2515 4160 2585 4180
rect 2645 4180 2740 4220
rect 2645 4160 2715 4180
rect 2430 4145 2486 4151
rect 2430 4085 2434 4145
rect 2515 4135 2715 4160
rect 2770 4151 2800 4339
rect 2744 4145 2800 4151
rect 2486 4085 2744 4105
rect 2796 4085 2800 4145
rect 2430 4075 2800 4085
rect 2830 4405 3200 4415
rect 2830 4345 2834 4405
rect 2886 4385 3144 4405
rect 2830 4339 2886 4345
rect 2830 4151 2860 4339
rect 2915 4330 3115 4355
rect 3196 4345 3200 4405
rect 3144 4339 3200 4345
rect 2915 4310 2985 4330
rect 2890 4270 2985 4310
rect 3045 4310 3115 4330
rect 3045 4270 3140 4310
rect 2890 4220 3140 4270
rect 2890 4180 2985 4220
rect 2915 4160 2985 4180
rect 3045 4180 3140 4220
rect 3045 4160 3115 4180
rect 2830 4145 2886 4151
rect 2830 4085 2834 4145
rect 2915 4135 3115 4160
rect 3170 4151 3200 4339
rect 3144 4145 3200 4151
rect 2886 4085 3144 4105
rect 3196 4085 3200 4145
rect 2830 4075 3200 4085
rect 3230 4405 3600 4415
rect 3230 4345 3234 4405
rect 3286 4385 3544 4405
rect 3230 4339 3286 4345
rect 3230 4151 3260 4339
rect 3315 4330 3515 4355
rect 3596 4345 3600 4405
rect 3544 4339 3600 4345
rect 3315 4310 3385 4330
rect 3290 4270 3385 4310
rect 3445 4310 3515 4330
rect 3445 4270 3540 4310
rect 3290 4220 3540 4270
rect 3290 4180 3385 4220
rect 3315 4160 3385 4180
rect 3445 4180 3540 4220
rect 3445 4160 3515 4180
rect 3230 4145 3286 4151
rect 3230 4085 3234 4145
rect 3315 4135 3515 4160
rect 3570 4151 3600 4339
rect 3544 4145 3600 4151
rect 3286 4085 3544 4105
rect 3596 4085 3600 4145
rect 3230 4075 3600 4085
rect 3630 4405 4000 4415
rect 3630 4345 3634 4405
rect 3686 4385 3944 4405
rect 3630 4339 3686 4345
rect 3630 4151 3660 4339
rect 3715 4330 3915 4355
rect 3996 4345 4000 4405
rect 3944 4339 4000 4345
rect 3715 4310 3785 4330
rect 3690 4270 3785 4310
rect 3845 4310 3915 4330
rect 3845 4270 3940 4310
rect 3690 4220 3940 4270
rect 3690 4180 3785 4220
rect 3715 4160 3785 4180
rect 3845 4180 3940 4220
rect 3845 4160 3915 4180
rect 3630 4145 3686 4151
rect 3630 4085 3634 4145
rect 3715 4135 3915 4160
rect 3970 4151 4000 4339
rect 3944 4145 4000 4151
rect 3686 4085 3944 4105
rect 3996 4085 4000 4145
rect 3630 4075 4000 4085
rect 4030 4405 4400 4415
rect 4030 4345 4034 4405
rect 4086 4385 4344 4405
rect 4030 4339 4086 4345
rect 4030 4151 4060 4339
rect 4115 4330 4315 4355
rect 4396 4345 4400 4405
rect 4344 4339 4400 4345
rect 4115 4310 4185 4330
rect 4090 4270 4185 4310
rect 4245 4310 4315 4330
rect 4245 4270 4340 4310
rect 4090 4220 4340 4270
rect 4090 4180 4185 4220
rect 4115 4160 4185 4180
rect 4245 4180 4340 4220
rect 4245 4160 4315 4180
rect 4030 4145 4086 4151
rect 4030 4085 4034 4145
rect 4115 4135 4315 4160
rect 4370 4151 4400 4339
rect 4344 4145 4400 4151
rect 4086 4085 4344 4105
rect 4396 4085 4400 4145
rect 4030 4075 4400 4085
rect 4430 4405 4800 4415
rect 4430 4345 4434 4405
rect 4486 4385 4744 4405
rect 4430 4339 4486 4345
rect 4430 4151 4460 4339
rect 4515 4330 4715 4355
rect 4796 4345 4800 4405
rect 4744 4339 4800 4345
rect 4515 4310 4585 4330
rect 4490 4270 4585 4310
rect 4645 4310 4715 4330
rect 4645 4270 4740 4310
rect 4490 4220 4740 4270
rect 4490 4180 4585 4220
rect 4515 4160 4585 4180
rect 4645 4180 4740 4220
rect 4645 4160 4715 4180
rect 4430 4145 4486 4151
rect 4430 4085 4434 4145
rect 4515 4135 4715 4160
rect 4770 4151 4800 4339
rect 4744 4145 4800 4151
rect 4486 4085 4744 4105
rect 4796 4085 4800 4145
rect 4430 4075 4800 4085
rect 4830 4405 5200 4415
rect 4830 4345 4834 4405
rect 4886 4385 5144 4405
rect 4830 4339 4886 4345
rect 4830 4151 4860 4339
rect 4915 4330 5115 4355
rect 5196 4345 5200 4405
rect 5144 4339 5200 4345
rect 4915 4310 4985 4330
rect 4890 4270 4985 4310
rect 5045 4310 5115 4330
rect 5045 4270 5140 4310
rect 4890 4220 5140 4270
rect 4890 4180 4985 4220
rect 4915 4160 4985 4180
rect 5045 4180 5140 4220
rect 5045 4160 5115 4180
rect 4830 4145 4886 4151
rect 4830 4085 4834 4145
rect 4915 4135 5115 4160
rect 5170 4151 5200 4339
rect 5144 4145 5200 4151
rect 4886 4085 5144 4105
rect 5196 4085 5200 4145
rect 4830 4075 5200 4085
rect 5230 4405 5600 4415
rect 5230 4345 5234 4405
rect 5286 4385 5544 4405
rect 5230 4339 5286 4345
rect 5230 4151 5260 4339
rect 5315 4330 5515 4355
rect 5596 4345 5600 4405
rect 5544 4339 5600 4345
rect 5315 4310 5385 4330
rect 5290 4270 5385 4310
rect 5445 4310 5515 4330
rect 5445 4270 5540 4310
rect 5290 4220 5540 4270
rect 5290 4180 5385 4220
rect 5315 4160 5385 4180
rect 5445 4180 5540 4220
rect 5445 4160 5515 4180
rect 5230 4145 5286 4151
rect 5230 4085 5234 4145
rect 5315 4135 5515 4160
rect 5570 4151 5600 4339
rect 5544 4145 5600 4151
rect 5286 4085 5544 4105
rect 5596 4085 5600 4145
rect 5230 4075 5600 4085
rect 5630 4405 6000 4415
rect 5630 4345 5634 4405
rect 5686 4385 5944 4405
rect 5630 4339 5686 4345
rect 5630 4151 5660 4339
rect 5715 4330 5915 4355
rect 5996 4345 6000 4405
rect 5944 4339 6000 4345
rect 5715 4310 5785 4330
rect 5690 4270 5785 4310
rect 5845 4310 5915 4330
rect 5845 4270 5940 4310
rect 5690 4220 5940 4270
rect 5690 4180 5785 4220
rect 5715 4160 5785 4180
rect 5845 4180 5940 4220
rect 5845 4160 5915 4180
rect 5630 4145 5686 4151
rect 5630 4085 5634 4145
rect 5715 4135 5915 4160
rect 5970 4151 6000 4339
rect 5944 4145 6000 4151
rect 5686 4085 5944 4105
rect 5996 4085 6000 4145
rect 5630 4075 6000 4085
rect 6030 4405 6400 4415
rect 6030 4345 6034 4405
rect 6086 4385 6344 4405
rect 6030 4339 6086 4345
rect 6030 4151 6060 4339
rect 6115 4330 6315 4355
rect 6396 4345 6400 4405
rect 6344 4339 6400 4345
rect 6115 4310 6185 4330
rect 6090 4270 6185 4310
rect 6245 4310 6315 4330
rect 6245 4270 6340 4310
rect 6090 4220 6340 4270
rect 6090 4180 6185 4220
rect 6115 4160 6185 4180
rect 6245 4180 6340 4220
rect 6245 4160 6315 4180
rect 6030 4145 6086 4151
rect 6030 4085 6034 4145
rect 6115 4135 6315 4160
rect 6370 4151 6400 4339
rect 6344 4145 6400 4151
rect 6086 4085 6344 4105
rect 6396 4085 6400 4145
rect 6030 4075 6400 4085
rect 6430 4405 6800 4415
rect 6430 4345 6434 4405
rect 6486 4385 6744 4405
rect 6430 4339 6486 4345
rect 6430 4151 6460 4339
rect 6515 4330 6715 4355
rect 6796 4345 6800 4405
rect 6744 4339 6800 4345
rect 6515 4310 6585 4330
rect 6490 4270 6585 4310
rect 6645 4310 6715 4330
rect 6645 4270 6740 4310
rect 6490 4220 6740 4270
rect 6490 4180 6585 4220
rect 6515 4160 6585 4180
rect 6645 4180 6740 4220
rect 6645 4160 6715 4180
rect 6430 4145 6486 4151
rect 6430 4085 6434 4145
rect 6515 4135 6715 4160
rect 6770 4151 6800 4339
rect 6744 4145 6800 4151
rect 6486 4085 6744 4105
rect 6796 4085 6800 4145
rect 6430 4075 6800 4085
rect 6830 4405 7200 4415
rect 6830 4345 6834 4405
rect 6886 4385 7144 4405
rect 6830 4339 6886 4345
rect 6830 4151 6860 4339
rect 6915 4330 7115 4355
rect 7196 4345 7200 4405
rect 7144 4339 7200 4345
rect 6915 4310 6985 4330
rect 6890 4270 6985 4310
rect 7045 4310 7115 4330
rect 7045 4270 7140 4310
rect 6890 4220 7140 4270
rect 6890 4180 6985 4220
rect 6915 4160 6985 4180
rect 7045 4180 7140 4220
rect 7045 4160 7115 4180
rect 6830 4145 6886 4151
rect 6830 4085 6834 4145
rect 6915 4135 7115 4160
rect 7170 4151 7200 4339
rect 7144 4145 7200 4151
rect 6886 4085 7144 4105
rect 7196 4085 7200 4145
rect 6830 4075 7200 4085
rect 7230 4405 7600 4415
rect 7230 4345 7234 4405
rect 7286 4385 7544 4405
rect 7230 4339 7286 4345
rect 7230 4151 7260 4339
rect 7315 4330 7515 4355
rect 7596 4345 7600 4405
rect 7544 4339 7600 4345
rect 7315 4310 7385 4330
rect 7290 4270 7385 4310
rect 7445 4310 7515 4330
rect 7445 4270 7540 4310
rect 7290 4220 7540 4270
rect 7290 4180 7385 4220
rect 7315 4160 7385 4180
rect 7445 4180 7540 4220
rect 7445 4160 7515 4180
rect 7230 4145 7286 4151
rect 7230 4085 7234 4145
rect 7315 4135 7515 4160
rect 7570 4151 7600 4339
rect 7544 4145 7600 4151
rect 7286 4085 7544 4105
rect 7596 4085 7600 4145
rect 7230 4075 7600 4085
rect 7630 4405 8000 4415
rect 7630 4345 7634 4405
rect 7686 4385 7944 4405
rect 7630 4339 7686 4345
rect 7630 4151 7660 4339
rect 7715 4330 7915 4355
rect 7996 4345 8000 4405
rect 7944 4339 8000 4345
rect 7715 4310 7785 4330
rect 7690 4270 7785 4310
rect 7845 4310 7915 4330
rect 7845 4270 7940 4310
rect 7690 4220 7940 4270
rect 7690 4180 7785 4220
rect 7715 4160 7785 4180
rect 7845 4180 7940 4220
rect 7845 4160 7915 4180
rect 7630 4145 7686 4151
rect 7630 4085 7634 4145
rect 7715 4135 7915 4160
rect 7970 4151 8000 4339
rect 7944 4145 8000 4151
rect 7686 4085 7944 4105
rect 7996 4085 8000 4145
rect 7630 4075 8000 4085
rect 8030 4405 8400 4415
rect 8030 4345 8034 4405
rect 8086 4385 8344 4405
rect 8030 4339 8086 4345
rect 8030 4151 8060 4339
rect 8115 4330 8315 4355
rect 8396 4345 8400 4405
rect 8344 4339 8400 4345
rect 8115 4310 8185 4330
rect 8090 4270 8185 4310
rect 8245 4310 8315 4330
rect 8245 4270 8340 4310
rect 8090 4220 8340 4270
rect 8090 4180 8185 4220
rect 8115 4160 8185 4180
rect 8245 4180 8340 4220
rect 8245 4160 8315 4180
rect 8030 4145 8086 4151
rect 8030 4085 8034 4145
rect 8115 4135 8315 4160
rect 8370 4151 8400 4339
rect 8344 4145 8400 4151
rect 8086 4085 8344 4105
rect 8396 4085 8400 4145
rect 8030 4075 8400 4085
rect 8430 4405 8800 4415
rect 8430 4345 8434 4405
rect 8486 4385 8744 4405
rect 8430 4339 8486 4345
rect 8430 4151 8460 4339
rect 8515 4330 8715 4355
rect 8796 4345 8800 4405
rect 8744 4339 8800 4345
rect 8515 4310 8585 4330
rect 8490 4270 8585 4310
rect 8645 4310 8715 4330
rect 8645 4270 8740 4310
rect 8490 4220 8740 4270
rect 8490 4180 8585 4220
rect 8515 4160 8585 4180
rect 8645 4180 8740 4220
rect 8645 4160 8715 4180
rect 8430 4145 8486 4151
rect 8430 4085 8434 4145
rect 8515 4135 8715 4160
rect 8770 4151 8800 4339
rect 8744 4145 8800 4151
rect 8486 4085 8744 4105
rect 8796 4085 8800 4145
rect 8430 4075 8800 4085
rect 8830 4405 9200 4415
rect 8830 4345 8834 4405
rect 8886 4385 9144 4405
rect 8830 4339 8886 4345
rect 8830 4151 8860 4339
rect 8915 4330 9115 4355
rect 9196 4345 9200 4405
rect 9144 4339 9200 4345
rect 8915 4310 8985 4330
rect 8890 4270 8985 4310
rect 9045 4310 9115 4330
rect 9045 4270 9140 4310
rect 8890 4220 9140 4270
rect 8890 4180 8985 4220
rect 8915 4160 8985 4180
rect 9045 4180 9140 4220
rect 9045 4160 9115 4180
rect 8830 4145 8886 4151
rect 8830 4085 8834 4145
rect 8915 4135 9115 4160
rect 9170 4151 9200 4339
rect 9144 4145 9200 4151
rect 8886 4085 9144 4105
rect 9196 4085 9200 4145
rect 8830 4075 9200 4085
rect 9230 4405 9600 4415
rect 9230 4345 9234 4405
rect 9286 4385 9544 4405
rect 9230 4339 9286 4345
rect 9230 4151 9260 4339
rect 9315 4330 9515 4355
rect 9596 4345 9600 4405
rect 9544 4339 9600 4345
rect 9315 4310 9385 4330
rect 9290 4270 9385 4310
rect 9445 4310 9515 4330
rect 9445 4270 9540 4310
rect 9290 4220 9540 4270
rect 9290 4180 9385 4220
rect 9315 4160 9385 4180
rect 9445 4180 9540 4220
rect 9445 4160 9515 4180
rect 9230 4145 9286 4151
rect 9230 4085 9234 4145
rect 9315 4135 9515 4160
rect 9570 4151 9600 4339
rect 9544 4145 9600 4151
rect 9286 4085 9544 4105
rect 9596 4085 9600 4145
rect 9230 4075 9600 4085
rect 9630 4405 10000 4415
rect 9630 4345 9634 4405
rect 9686 4385 9944 4405
rect 9630 4339 9686 4345
rect 9630 4151 9660 4339
rect 9715 4330 9915 4355
rect 9996 4345 10000 4405
rect 9944 4339 10000 4345
rect 9715 4310 9785 4330
rect 9690 4270 9785 4310
rect 9845 4310 9915 4330
rect 9845 4270 9940 4310
rect 9690 4220 9940 4270
rect 9690 4180 9785 4220
rect 9715 4160 9785 4180
rect 9845 4180 9940 4220
rect 9845 4160 9915 4180
rect 9630 4145 9686 4151
rect 9630 4085 9634 4145
rect 9715 4135 9915 4160
rect 9970 4151 10000 4339
rect 9944 4145 10000 4151
rect 9686 4085 9944 4105
rect 9996 4085 10000 4145
rect 9630 4075 10000 4085
rect 10030 4405 10400 4415
rect 10030 4345 10034 4405
rect 10086 4385 10344 4405
rect 10030 4339 10086 4345
rect 10030 4151 10060 4339
rect 10115 4330 10315 4355
rect 10396 4345 10400 4405
rect 10344 4339 10400 4345
rect 10115 4310 10185 4330
rect 10090 4270 10185 4310
rect 10245 4310 10315 4330
rect 10245 4270 10340 4310
rect 10090 4220 10340 4270
rect 10090 4180 10185 4220
rect 10115 4160 10185 4180
rect 10245 4180 10340 4220
rect 10245 4160 10315 4180
rect 10030 4145 10086 4151
rect 10030 4085 10034 4145
rect 10115 4135 10315 4160
rect 10370 4151 10400 4339
rect 10344 4145 10400 4151
rect 10086 4085 10344 4105
rect 10396 4085 10400 4145
rect 10030 4075 10400 4085
rect 10430 4405 10800 4415
rect 10430 4345 10434 4405
rect 10486 4385 10744 4405
rect 10430 4339 10486 4345
rect 10430 4151 10460 4339
rect 10515 4330 10715 4355
rect 10796 4345 10800 4405
rect 10744 4339 10800 4345
rect 10515 4310 10585 4330
rect 10490 4270 10585 4310
rect 10645 4310 10715 4330
rect 10645 4270 10740 4310
rect 10490 4220 10740 4270
rect 10490 4180 10585 4220
rect 10515 4160 10585 4180
rect 10645 4180 10740 4220
rect 10645 4160 10715 4180
rect 10430 4145 10486 4151
rect 10430 4085 10434 4145
rect 10515 4135 10715 4160
rect 10770 4151 10800 4339
rect 10744 4145 10800 4151
rect 10486 4085 10744 4105
rect 10796 4085 10800 4145
rect 10430 4075 10800 4085
rect 10830 4405 11200 4415
rect 10830 4345 10834 4405
rect 10886 4385 11144 4405
rect 10830 4339 10886 4345
rect 10830 4151 10860 4339
rect 10915 4330 11115 4355
rect 11196 4345 11200 4405
rect 11144 4339 11200 4345
rect 10915 4310 10985 4330
rect 10890 4270 10985 4310
rect 11045 4310 11115 4330
rect 11045 4270 11140 4310
rect 10890 4220 11140 4270
rect 10890 4180 10985 4220
rect 10915 4160 10985 4180
rect 11045 4180 11140 4220
rect 11045 4160 11115 4180
rect 10830 4145 10886 4151
rect 10830 4085 10834 4145
rect 10915 4135 11115 4160
rect 11170 4151 11200 4339
rect 11144 4145 11200 4151
rect 10886 4085 11144 4105
rect 11196 4085 11200 4145
rect 10830 4075 11200 4085
rect 11230 4405 11600 4415
rect 11230 4345 11234 4405
rect 11286 4385 11544 4405
rect 11230 4339 11286 4345
rect 11230 4151 11260 4339
rect 11315 4330 11515 4355
rect 11596 4345 11600 4405
rect 11544 4339 11600 4345
rect 11315 4310 11385 4330
rect 11290 4270 11385 4310
rect 11445 4310 11515 4330
rect 11445 4270 11540 4310
rect 11290 4220 11540 4270
rect 11290 4180 11385 4220
rect 11315 4160 11385 4180
rect 11445 4180 11540 4220
rect 11445 4160 11515 4180
rect 11230 4145 11286 4151
rect 11230 4085 11234 4145
rect 11315 4135 11515 4160
rect 11570 4151 11600 4339
rect 11544 4145 11600 4151
rect 11286 4085 11544 4105
rect 11596 4085 11600 4145
rect 11230 4075 11600 4085
rect 11630 4405 12000 4415
rect 11630 4345 11634 4405
rect 11686 4385 11944 4405
rect 11630 4339 11686 4345
rect 11630 4151 11660 4339
rect 11715 4330 11915 4355
rect 11996 4345 12000 4405
rect 11944 4339 12000 4345
rect 11715 4310 11785 4330
rect 11690 4270 11785 4310
rect 11845 4310 11915 4330
rect 11845 4270 11940 4310
rect 11690 4220 11940 4270
rect 11690 4180 11785 4220
rect 11715 4160 11785 4180
rect 11845 4180 11940 4220
rect 11845 4160 11915 4180
rect 11630 4145 11686 4151
rect 11630 4085 11634 4145
rect 11715 4135 11915 4160
rect 11970 4151 12000 4339
rect 11944 4145 12000 4151
rect 11686 4085 11944 4105
rect 11996 4085 12000 4145
rect 11630 4075 12000 4085
rect 12030 4405 12400 4415
rect 12030 4345 12034 4405
rect 12086 4385 12344 4405
rect 12030 4339 12086 4345
rect 12030 4151 12060 4339
rect 12115 4330 12315 4355
rect 12396 4345 12400 4405
rect 12344 4339 12400 4345
rect 12115 4310 12185 4330
rect 12090 4270 12185 4310
rect 12245 4310 12315 4330
rect 12245 4270 12340 4310
rect 12090 4220 12340 4270
rect 12090 4180 12185 4220
rect 12115 4160 12185 4180
rect 12245 4180 12340 4220
rect 12245 4160 12315 4180
rect 12030 4145 12086 4151
rect 12030 4085 12034 4145
rect 12115 4135 12315 4160
rect 12370 4151 12400 4339
rect 12344 4145 12400 4151
rect 12086 4085 12344 4105
rect 12396 4085 12400 4145
rect 12030 4075 12400 4085
rect 12430 4405 12800 4415
rect 12430 4345 12434 4405
rect 12486 4385 12744 4405
rect 12430 4339 12486 4345
rect 12430 4151 12460 4339
rect 12515 4330 12715 4355
rect 12796 4345 12800 4405
rect 12744 4339 12800 4345
rect 12515 4310 12585 4330
rect 12490 4270 12585 4310
rect 12645 4310 12715 4330
rect 12645 4270 12740 4310
rect 12490 4220 12740 4270
rect 12490 4180 12585 4220
rect 12515 4160 12585 4180
rect 12645 4180 12740 4220
rect 12645 4160 12715 4180
rect 12430 4145 12486 4151
rect 12430 4085 12434 4145
rect 12515 4135 12715 4160
rect 12770 4151 12800 4339
rect 12744 4145 12800 4151
rect 12486 4085 12744 4105
rect 12796 4085 12800 4145
rect 12430 4075 12800 4085
rect 12830 4405 13200 4415
rect 12830 4345 12834 4405
rect 12886 4385 13144 4405
rect 12830 4339 12886 4345
rect 12830 4151 12860 4339
rect 12915 4330 13115 4355
rect 13196 4345 13200 4405
rect 13144 4339 13200 4345
rect 12915 4310 12985 4330
rect 12890 4270 12985 4310
rect 13045 4310 13115 4330
rect 13045 4270 13140 4310
rect 12890 4220 13140 4270
rect 12890 4180 12985 4220
rect 12915 4160 12985 4180
rect 13045 4180 13140 4220
rect 13045 4160 13115 4180
rect 12830 4145 12886 4151
rect 12830 4085 12834 4145
rect 12915 4135 13115 4160
rect 13170 4151 13200 4339
rect 13144 4145 13200 4151
rect 12886 4085 13144 4105
rect 13196 4085 13200 4145
rect 12830 4075 13200 4085
rect -370 4035 0 4045
rect -370 3975 -366 4035
rect -314 4015 -56 4035
rect -370 3969 -314 3975
rect -370 3781 -340 3969
rect -285 3960 -85 3985
rect -4 3975 0 4035
rect -56 3969 0 3975
rect -285 3940 -215 3960
rect -310 3900 -215 3940
rect -155 3940 -85 3960
rect -155 3900 -60 3940
rect -310 3850 -60 3900
rect -310 3810 -215 3850
rect -285 3790 -215 3810
rect -155 3810 -60 3850
rect -155 3790 -85 3810
rect -370 3775 -314 3781
rect -370 3715 -366 3775
rect -285 3765 -85 3790
rect -30 3781 0 3969
rect -56 3775 0 3781
rect -314 3715 -56 3735
rect -4 3715 0 3775
rect -370 3705 0 3715
rect 30 4035 400 4045
rect 30 3975 34 4035
rect 86 4015 344 4035
rect 30 3969 86 3975
rect 30 3781 60 3969
rect 115 3960 315 3985
rect 396 3975 400 4035
rect 344 3969 400 3975
rect 115 3940 185 3960
rect 90 3900 185 3940
rect 245 3940 315 3960
rect 245 3900 340 3940
rect 90 3850 340 3900
rect 90 3810 185 3850
rect 115 3790 185 3810
rect 245 3810 340 3850
rect 245 3790 315 3810
rect 30 3775 86 3781
rect 30 3715 34 3775
rect 115 3765 315 3790
rect 370 3781 400 3969
rect 344 3775 400 3781
rect 86 3715 344 3735
rect 396 3715 400 3775
rect 30 3705 400 3715
rect 430 4035 800 4045
rect 430 3975 434 4035
rect 486 4015 744 4035
rect 430 3969 486 3975
rect 430 3781 460 3969
rect 515 3960 715 3985
rect 796 3975 800 4035
rect 744 3969 800 3975
rect 515 3940 585 3960
rect 490 3900 585 3940
rect 645 3940 715 3960
rect 645 3900 740 3940
rect 490 3850 740 3900
rect 490 3810 585 3850
rect 515 3790 585 3810
rect 645 3810 740 3850
rect 645 3790 715 3810
rect 430 3775 486 3781
rect 430 3715 434 3775
rect 515 3765 715 3790
rect 770 3781 800 3969
rect 744 3775 800 3781
rect 486 3715 744 3735
rect 796 3715 800 3775
rect 430 3705 800 3715
rect 830 4035 1200 4045
rect 830 3975 834 4035
rect 886 4015 1144 4035
rect 830 3969 886 3975
rect 830 3781 860 3969
rect 915 3960 1115 3985
rect 1196 3975 1200 4035
rect 1144 3969 1200 3975
rect 915 3940 985 3960
rect 890 3900 985 3940
rect 1045 3940 1115 3960
rect 1045 3900 1140 3940
rect 890 3850 1140 3900
rect 890 3810 985 3850
rect 915 3790 985 3810
rect 1045 3810 1140 3850
rect 1045 3790 1115 3810
rect 830 3775 886 3781
rect 830 3715 834 3775
rect 915 3765 1115 3790
rect 1170 3781 1200 3969
rect 1144 3775 1200 3781
rect 886 3715 1144 3735
rect 1196 3715 1200 3775
rect 830 3705 1200 3715
rect 1230 4035 1600 4045
rect 1230 3975 1234 4035
rect 1286 4015 1544 4035
rect 1230 3969 1286 3975
rect 1230 3781 1260 3969
rect 1315 3960 1515 3985
rect 1596 3975 1600 4035
rect 1544 3969 1600 3975
rect 1315 3940 1385 3960
rect 1290 3900 1385 3940
rect 1445 3940 1515 3960
rect 1445 3900 1540 3940
rect 1290 3850 1540 3900
rect 1290 3810 1385 3850
rect 1315 3790 1385 3810
rect 1445 3810 1540 3850
rect 1445 3790 1515 3810
rect 1230 3775 1286 3781
rect 1230 3715 1234 3775
rect 1315 3765 1515 3790
rect 1570 3781 1600 3969
rect 1544 3775 1600 3781
rect 1286 3715 1544 3735
rect 1596 3715 1600 3775
rect 1230 3705 1600 3715
rect 1630 4035 2000 4045
rect 1630 3975 1634 4035
rect 1686 4015 1944 4035
rect 1630 3969 1686 3975
rect 1630 3781 1660 3969
rect 1715 3960 1915 3985
rect 1996 3975 2000 4035
rect 1944 3969 2000 3975
rect 1715 3940 1785 3960
rect 1690 3900 1785 3940
rect 1845 3940 1915 3960
rect 1845 3900 1940 3940
rect 1690 3850 1940 3900
rect 1690 3810 1785 3850
rect 1715 3790 1785 3810
rect 1845 3810 1940 3850
rect 1845 3790 1915 3810
rect 1630 3775 1686 3781
rect 1630 3715 1634 3775
rect 1715 3765 1915 3790
rect 1970 3781 2000 3969
rect 1944 3775 2000 3781
rect 1686 3715 1944 3735
rect 1996 3715 2000 3775
rect 1630 3705 2000 3715
rect 2030 4035 2400 4045
rect 2030 3975 2034 4035
rect 2086 4015 2344 4035
rect 2030 3969 2086 3975
rect 2030 3781 2060 3969
rect 2115 3960 2315 3985
rect 2396 3975 2400 4035
rect 2344 3969 2400 3975
rect 2115 3940 2185 3960
rect 2090 3900 2185 3940
rect 2245 3940 2315 3960
rect 2245 3900 2340 3940
rect 2090 3850 2340 3900
rect 2090 3810 2185 3850
rect 2115 3790 2185 3810
rect 2245 3810 2340 3850
rect 2245 3790 2315 3810
rect 2030 3775 2086 3781
rect 2030 3715 2034 3775
rect 2115 3765 2315 3790
rect 2370 3781 2400 3969
rect 2344 3775 2400 3781
rect 2086 3715 2344 3735
rect 2396 3715 2400 3775
rect 2030 3705 2400 3715
rect 2430 4035 2800 4045
rect 2430 3975 2434 4035
rect 2486 4015 2744 4035
rect 2430 3969 2486 3975
rect 2430 3781 2460 3969
rect 2515 3960 2715 3985
rect 2796 3975 2800 4035
rect 2744 3969 2800 3975
rect 2515 3940 2585 3960
rect 2490 3900 2585 3940
rect 2645 3940 2715 3960
rect 2645 3900 2740 3940
rect 2490 3850 2740 3900
rect 2490 3810 2585 3850
rect 2515 3790 2585 3810
rect 2645 3810 2740 3850
rect 2645 3790 2715 3810
rect 2430 3775 2486 3781
rect 2430 3715 2434 3775
rect 2515 3765 2715 3790
rect 2770 3781 2800 3969
rect 2744 3775 2800 3781
rect 2486 3715 2744 3735
rect 2796 3715 2800 3775
rect 2430 3705 2800 3715
rect 2830 4035 3200 4045
rect 2830 3975 2834 4035
rect 2886 4015 3144 4035
rect 2830 3969 2886 3975
rect 2830 3781 2860 3969
rect 2915 3960 3115 3985
rect 3196 3975 3200 4035
rect 3144 3969 3200 3975
rect 2915 3940 2985 3960
rect 2890 3900 2985 3940
rect 3045 3940 3115 3960
rect 3045 3900 3140 3940
rect 2890 3850 3140 3900
rect 2890 3810 2985 3850
rect 2915 3790 2985 3810
rect 3045 3810 3140 3850
rect 3045 3790 3115 3810
rect 2830 3775 2886 3781
rect 2830 3715 2834 3775
rect 2915 3765 3115 3790
rect 3170 3781 3200 3969
rect 3144 3775 3200 3781
rect 2886 3715 3144 3735
rect 3196 3715 3200 3775
rect 2830 3705 3200 3715
rect 3230 4035 3600 4045
rect 3230 3975 3234 4035
rect 3286 4015 3544 4035
rect 3230 3969 3286 3975
rect 3230 3781 3260 3969
rect 3315 3960 3515 3985
rect 3596 3975 3600 4035
rect 3544 3969 3600 3975
rect 3315 3940 3385 3960
rect 3290 3900 3385 3940
rect 3445 3940 3515 3960
rect 3445 3900 3540 3940
rect 3290 3850 3540 3900
rect 3290 3810 3385 3850
rect 3315 3790 3385 3810
rect 3445 3810 3540 3850
rect 3445 3790 3515 3810
rect 3230 3775 3286 3781
rect 3230 3715 3234 3775
rect 3315 3765 3515 3790
rect 3570 3781 3600 3969
rect 3544 3775 3600 3781
rect 3286 3715 3544 3735
rect 3596 3715 3600 3775
rect 3230 3705 3600 3715
rect 3630 4035 4000 4045
rect 3630 3975 3634 4035
rect 3686 4015 3944 4035
rect 3630 3969 3686 3975
rect 3630 3781 3660 3969
rect 3715 3960 3915 3985
rect 3996 3975 4000 4035
rect 3944 3969 4000 3975
rect 3715 3940 3785 3960
rect 3690 3900 3785 3940
rect 3845 3940 3915 3960
rect 3845 3900 3940 3940
rect 3690 3850 3940 3900
rect 3690 3810 3785 3850
rect 3715 3790 3785 3810
rect 3845 3810 3940 3850
rect 3845 3790 3915 3810
rect 3630 3775 3686 3781
rect 3630 3715 3634 3775
rect 3715 3765 3915 3790
rect 3970 3781 4000 3969
rect 3944 3775 4000 3781
rect 3686 3715 3944 3735
rect 3996 3715 4000 3775
rect 3630 3705 4000 3715
rect 4030 4035 4400 4045
rect 4030 3975 4034 4035
rect 4086 4015 4344 4035
rect 4030 3969 4086 3975
rect 4030 3781 4060 3969
rect 4115 3960 4315 3985
rect 4396 3975 4400 4035
rect 4344 3969 4400 3975
rect 4115 3940 4185 3960
rect 4090 3900 4185 3940
rect 4245 3940 4315 3960
rect 4245 3900 4340 3940
rect 4090 3850 4340 3900
rect 4090 3810 4185 3850
rect 4115 3790 4185 3810
rect 4245 3810 4340 3850
rect 4245 3790 4315 3810
rect 4030 3775 4086 3781
rect 4030 3715 4034 3775
rect 4115 3765 4315 3790
rect 4370 3781 4400 3969
rect 4344 3775 4400 3781
rect 4086 3715 4344 3735
rect 4396 3715 4400 3775
rect 4030 3705 4400 3715
rect 4430 4035 4800 4045
rect 4430 3975 4434 4035
rect 4486 4015 4744 4035
rect 4430 3969 4486 3975
rect 4430 3781 4460 3969
rect 4515 3960 4715 3985
rect 4796 3975 4800 4035
rect 4744 3969 4800 3975
rect 4515 3940 4585 3960
rect 4490 3900 4585 3940
rect 4645 3940 4715 3960
rect 4645 3900 4740 3940
rect 4490 3850 4740 3900
rect 4490 3810 4585 3850
rect 4515 3790 4585 3810
rect 4645 3810 4740 3850
rect 4645 3790 4715 3810
rect 4430 3775 4486 3781
rect 4430 3715 4434 3775
rect 4515 3765 4715 3790
rect 4770 3781 4800 3969
rect 4744 3775 4800 3781
rect 4486 3715 4744 3735
rect 4796 3715 4800 3775
rect 4430 3705 4800 3715
rect 4830 4035 5200 4045
rect 4830 3975 4834 4035
rect 4886 4015 5144 4035
rect 4830 3969 4886 3975
rect 4830 3781 4860 3969
rect 4915 3960 5115 3985
rect 5196 3975 5200 4035
rect 5144 3969 5200 3975
rect 4915 3940 4985 3960
rect 4890 3900 4985 3940
rect 5045 3940 5115 3960
rect 5045 3900 5140 3940
rect 4890 3850 5140 3900
rect 4890 3810 4985 3850
rect 4915 3790 4985 3810
rect 5045 3810 5140 3850
rect 5045 3790 5115 3810
rect 4830 3775 4886 3781
rect 4830 3715 4834 3775
rect 4915 3765 5115 3790
rect 5170 3781 5200 3969
rect 5144 3775 5200 3781
rect 4886 3715 5144 3735
rect 5196 3715 5200 3775
rect 4830 3705 5200 3715
rect 5230 4035 5600 4045
rect 5230 3975 5234 4035
rect 5286 4015 5544 4035
rect 5230 3969 5286 3975
rect 5230 3781 5260 3969
rect 5315 3960 5515 3985
rect 5596 3975 5600 4035
rect 5544 3969 5600 3975
rect 5315 3940 5385 3960
rect 5290 3900 5385 3940
rect 5445 3940 5515 3960
rect 5445 3900 5540 3940
rect 5290 3850 5540 3900
rect 5290 3810 5385 3850
rect 5315 3790 5385 3810
rect 5445 3810 5540 3850
rect 5445 3790 5515 3810
rect 5230 3775 5286 3781
rect 5230 3715 5234 3775
rect 5315 3765 5515 3790
rect 5570 3781 5600 3969
rect 5544 3775 5600 3781
rect 5286 3715 5544 3735
rect 5596 3715 5600 3775
rect 5230 3705 5600 3715
rect 5630 4035 6000 4045
rect 5630 3975 5634 4035
rect 5686 4015 5944 4035
rect 5630 3969 5686 3975
rect 5630 3781 5660 3969
rect 5715 3960 5915 3985
rect 5996 3975 6000 4035
rect 5944 3969 6000 3975
rect 5715 3940 5785 3960
rect 5690 3900 5785 3940
rect 5845 3940 5915 3960
rect 5845 3900 5940 3940
rect 5690 3850 5940 3900
rect 5690 3810 5785 3850
rect 5715 3790 5785 3810
rect 5845 3810 5940 3850
rect 5845 3790 5915 3810
rect 5630 3775 5686 3781
rect 5630 3715 5634 3775
rect 5715 3765 5915 3790
rect 5970 3781 6000 3969
rect 5944 3775 6000 3781
rect 5686 3715 5944 3735
rect 5996 3715 6000 3775
rect 5630 3705 6000 3715
rect 6030 4035 6400 4045
rect 6030 3975 6034 4035
rect 6086 4015 6344 4035
rect 6030 3969 6086 3975
rect 6030 3781 6060 3969
rect 6115 3960 6315 3985
rect 6396 3975 6400 4035
rect 6344 3969 6400 3975
rect 6115 3940 6185 3960
rect 6090 3900 6185 3940
rect 6245 3940 6315 3960
rect 6245 3900 6340 3940
rect 6090 3850 6340 3900
rect 6090 3810 6185 3850
rect 6115 3790 6185 3810
rect 6245 3810 6340 3850
rect 6245 3790 6315 3810
rect 6030 3775 6086 3781
rect 6030 3715 6034 3775
rect 6115 3765 6315 3790
rect 6370 3781 6400 3969
rect 6344 3775 6400 3781
rect 6086 3715 6344 3735
rect 6396 3715 6400 3775
rect 6030 3705 6400 3715
rect 6430 4035 6800 4045
rect 6430 3975 6434 4035
rect 6486 4015 6744 4035
rect 6430 3969 6486 3975
rect 6430 3781 6460 3969
rect 6515 3960 6715 3985
rect 6796 3975 6800 4035
rect 6744 3969 6800 3975
rect 6515 3940 6585 3960
rect 6490 3900 6585 3940
rect 6645 3940 6715 3960
rect 6645 3900 6740 3940
rect 6490 3850 6740 3900
rect 6490 3810 6585 3850
rect 6515 3790 6585 3810
rect 6645 3810 6740 3850
rect 6645 3790 6715 3810
rect 6430 3775 6486 3781
rect 6430 3715 6434 3775
rect 6515 3765 6715 3790
rect 6770 3781 6800 3969
rect 6744 3775 6800 3781
rect 6486 3715 6744 3735
rect 6796 3715 6800 3775
rect 6430 3705 6800 3715
rect 6830 4035 7200 4045
rect 6830 3975 6834 4035
rect 6886 4015 7144 4035
rect 6830 3969 6886 3975
rect 6830 3781 6860 3969
rect 6915 3960 7115 3985
rect 7196 3975 7200 4035
rect 7144 3969 7200 3975
rect 6915 3940 6985 3960
rect 6890 3900 6985 3940
rect 7045 3940 7115 3960
rect 7045 3900 7140 3940
rect 6890 3850 7140 3900
rect 6890 3810 6985 3850
rect 6915 3790 6985 3810
rect 7045 3810 7140 3850
rect 7045 3790 7115 3810
rect 6830 3775 6886 3781
rect 6830 3715 6834 3775
rect 6915 3765 7115 3790
rect 7170 3781 7200 3969
rect 7144 3775 7200 3781
rect 6886 3715 7144 3735
rect 7196 3715 7200 3775
rect 6830 3705 7200 3715
rect 7230 4035 7600 4045
rect 7230 3975 7234 4035
rect 7286 4015 7544 4035
rect 7230 3969 7286 3975
rect 7230 3781 7260 3969
rect 7315 3960 7515 3985
rect 7596 3975 7600 4035
rect 7544 3969 7600 3975
rect 7315 3940 7385 3960
rect 7290 3900 7385 3940
rect 7445 3940 7515 3960
rect 7445 3900 7540 3940
rect 7290 3850 7540 3900
rect 7290 3810 7385 3850
rect 7315 3790 7385 3810
rect 7445 3810 7540 3850
rect 7445 3790 7515 3810
rect 7230 3775 7286 3781
rect 7230 3715 7234 3775
rect 7315 3765 7515 3790
rect 7570 3781 7600 3969
rect 7544 3775 7600 3781
rect 7286 3715 7544 3735
rect 7596 3715 7600 3775
rect 7230 3705 7600 3715
rect 7630 4035 8000 4045
rect 7630 3975 7634 4035
rect 7686 4015 7944 4035
rect 7630 3969 7686 3975
rect 7630 3781 7660 3969
rect 7715 3960 7915 3985
rect 7996 3975 8000 4035
rect 7944 3969 8000 3975
rect 7715 3940 7785 3960
rect 7690 3900 7785 3940
rect 7845 3940 7915 3960
rect 7845 3900 7940 3940
rect 7690 3850 7940 3900
rect 7690 3810 7785 3850
rect 7715 3790 7785 3810
rect 7845 3810 7940 3850
rect 7845 3790 7915 3810
rect 7630 3775 7686 3781
rect 7630 3715 7634 3775
rect 7715 3765 7915 3790
rect 7970 3781 8000 3969
rect 7944 3775 8000 3781
rect 7686 3715 7944 3735
rect 7996 3715 8000 3775
rect 7630 3705 8000 3715
rect 8030 4035 8400 4045
rect 8030 3975 8034 4035
rect 8086 4015 8344 4035
rect 8030 3969 8086 3975
rect 8030 3781 8060 3969
rect 8115 3960 8315 3985
rect 8396 3975 8400 4035
rect 8344 3969 8400 3975
rect 8115 3940 8185 3960
rect 8090 3900 8185 3940
rect 8245 3940 8315 3960
rect 8245 3900 8340 3940
rect 8090 3850 8340 3900
rect 8090 3810 8185 3850
rect 8115 3790 8185 3810
rect 8245 3810 8340 3850
rect 8245 3790 8315 3810
rect 8030 3775 8086 3781
rect 8030 3715 8034 3775
rect 8115 3765 8315 3790
rect 8370 3781 8400 3969
rect 8344 3775 8400 3781
rect 8086 3715 8344 3735
rect 8396 3715 8400 3775
rect 8030 3705 8400 3715
rect 8430 4035 8800 4045
rect 8430 3975 8434 4035
rect 8486 4015 8744 4035
rect 8430 3969 8486 3975
rect 8430 3781 8460 3969
rect 8515 3960 8715 3985
rect 8796 3975 8800 4035
rect 8744 3969 8800 3975
rect 8515 3940 8585 3960
rect 8490 3900 8585 3940
rect 8645 3940 8715 3960
rect 8645 3900 8740 3940
rect 8490 3850 8740 3900
rect 8490 3810 8585 3850
rect 8515 3790 8585 3810
rect 8645 3810 8740 3850
rect 8645 3790 8715 3810
rect 8430 3775 8486 3781
rect 8430 3715 8434 3775
rect 8515 3765 8715 3790
rect 8770 3781 8800 3969
rect 8744 3775 8800 3781
rect 8486 3715 8744 3735
rect 8796 3715 8800 3775
rect 8430 3705 8800 3715
rect 8830 4035 9200 4045
rect 8830 3975 8834 4035
rect 8886 4015 9144 4035
rect 8830 3969 8886 3975
rect 8830 3781 8860 3969
rect 8915 3960 9115 3985
rect 9196 3975 9200 4035
rect 9144 3969 9200 3975
rect 8915 3940 8985 3960
rect 8890 3900 8985 3940
rect 9045 3940 9115 3960
rect 9045 3900 9140 3940
rect 8890 3850 9140 3900
rect 8890 3810 8985 3850
rect 8915 3790 8985 3810
rect 9045 3810 9140 3850
rect 9045 3790 9115 3810
rect 8830 3775 8886 3781
rect 8830 3715 8834 3775
rect 8915 3765 9115 3790
rect 9170 3781 9200 3969
rect 9144 3775 9200 3781
rect 8886 3715 9144 3735
rect 9196 3715 9200 3775
rect 8830 3705 9200 3715
rect 9230 4035 9600 4045
rect 9230 3975 9234 4035
rect 9286 4015 9544 4035
rect 9230 3969 9286 3975
rect 9230 3781 9260 3969
rect 9315 3960 9515 3985
rect 9596 3975 9600 4035
rect 9544 3969 9600 3975
rect 9315 3940 9385 3960
rect 9290 3900 9385 3940
rect 9445 3940 9515 3960
rect 9445 3900 9540 3940
rect 9290 3850 9540 3900
rect 9290 3810 9385 3850
rect 9315 3790 9385 3810
rect 9445 3810 9540 3850
rect 9445 3790 9515 3810
rect 9230 3775 9286 3781
rect 9230 3715 9234 3775
rect 9315 3765 9515 3790
rect 9570 3781 9600 3969
rect 9544 3775 9600 3781
rect 9286 3715 9544 3735
rect 9596 3715 9600 3775
rect 9230 3705 9600 3715
rect 9630 4035 10000 4045
rect 9630 3975 9634 4035
rect 9686 4015 9944 4035
rect 9630 3969 9686 3975
rect 9630 3781 9660 3969
rect 9715 3960 9915 3985
rect 9996 3975 10000 4035
rect 9944 3969 10000 3975
rect 9715 3940 9785 3960
rect 9690 3900 9785 3940
rect 9845 3940 9915 3960
rect 9845 3900 9940 3940
rect 9690 3850 9940 3900
rect 9690 3810 9785 3850
rect 9715 3790 9785 3810
rect 9845 3810 9940 3850
rect 9845 3790 9915 3810
rect 9630 3775 9686 3781
rect 9630 3715 9634 3775
rect 9715 3765 9915 3790
rect 9970 3781 10000 3969
rect 9944 3775 10000 3781
rect 9686 3715 9944 3735
rect 9996 3715 10000 3775
rect 9630 3705 10000 3715
rect 10030 4035 10400 4045
rect 10030 3975 10034 4035
rect 10086 4015 10344 4035
rect 10030 3969 10086 3975
rect 10030 3781 10060 3969
rect 10115 3960 10315 3985
rect 10396 3975 10400 4035
rect 10344 3969 10400 3975
rect 10115 3940 10185 3960
rect 10090 3900 10185 3940
rect 10245 3940 10315 3960
rect 10245 3900 10340 3940
rect 10090 3850 10340 3900
rect 10090 3810 10185 3850
rect 10115 3790 10185 3810
rect 10245 3810 10340 3850
rect 10245 3790 10315 3810
rect 10030 3775 10086 3781
rect 10030 3715 10034 3775
rect 10115 3765 10315 3790
rect 10370 3781 10400 3969
rect 10344 3775 10400 3781
rect 10086 3715 10344 3735
rect 10396 3715 10400 3775
rect 10030 3705 10400 3715
rect 10430 4035 10800 4045
rect 10430 3975 10434 4035
rect 10486 4015 10744 4035
rect 10430 3969 10486 3975
rect 10430 3781 10460 3969
rect 10515 3960 10715 3985
rect 10796 3975 10800 4035
rect 10744 3969 10800 3975
rect 10515 3940 10585 3960
rect 10490 3900 10585 3940
rect 10645 3940 10715 3960
rect 10645 3900 10740 3940
rect 10490 3850 10740 3900
rect 10490 3810 10585 3850
rect 10515 3790 10585 3810
rect 10645 3810 10740 3850
rect 10645 3790 10715 3810
rect 10430 3775 10486 3781
rect 10430 3715 10434 3775
rect 10515 3765 10715 3790
rect 10770 3781 10800 3969
rect 10744 3775 10800 3781
rect 10486 3715 10744 3735
rect 10796 3715 10800 3775
rect 10430 3705 10800 3715
rect 10830 4035 11200 4045
rect 10830 3975 10834 4035
rect 10886 4015 11144 4035
rect 10830 3969 10886 3975
rect 10830 3781 10860 3969
rect 10915 3960 11115 3985
rect 11196 3975 11200 4035
rect 11144 3969 11200 3975
rect 10915 3940 10985 3960
rect 10890 3900 10985 3940
rect 11045 3940 11115 3960
rect 11045 3900 11140 3940
rect 10890 3850 11140 3900
rect 10890 3810 10985 3850
rect 10915 3790 10985 3810
rect 11045 3810 11140 3850
rect 11045 3790 11115 3810
rect 10830 3775 10886 3781
rect 10830 3715 10834 3775
rect 10915 3765 11115 3790
rect 11170 3781 11200 3969
rect 11144 3775 11200 3781
rect 10886 3715 11144 3735
rect 11196 3715 11200 3775
rect 10830 3705 11200 3715
rect 11230 4035 11600 4045
rect 11230 3975 11234 4035
rect 11286 4015 11544 4035
rect 11230 3969 11286 3975
rect 11230 3781 11260 3969
rect 11315 3960 11515 3985
rect 11596 3975 11600 4035
rect 11544 3969 11600 3975
rect 11315 3940 11385 3960
rect 11290 3900 11385 3940
rect 11445 3940 11515 3960
rect 11445 3900 11540 3940
rect 11290 3850 11540 3900
rect 11290 3810 11385 3850
rect 11315 3790 11385 3810
rect 11445 3810 11540 3850
rect 11445 3790 11515 3810
rect 11230 3775 11286 3781
rect 11230 3715 11234 3775
rect 11315 3765 11515 3790
rect 11570 3781 11600 3969
rect 11544 3775 11600 3781
rect 11286 3715 11544 3735
rect 11596 3715 11600 3775
rect 11230 3705 11600 3715
rect 11630 4035 12000 4045
rect 11630 3975 11634 4035
rect 11686 4015 11944 4035
rect 11630 3969 11686 3975
rect 11630 3781 11660 3969
rect 11715 3960 11915 3985
rect 11996 3975 12000 4035
rect 11944 3969 12000 3975
rect 11715 3940 11785 3960
rect 11690 3900 11785 3940
rect 11845 3940 11915 3960
rect 11845 3900 11940 3940
rect 11690 3850 11940 3900
rect 11690 3810 11785 3850
rect 11715 3790 11785 3810
rect 11845 3810 11940 3850
rect 11845 3790 11915 3810
rect 11630 3775 11686 3781
rect 11630 3715 11634 3775
rect 11715 3765 11915 3790
rect 11970 3781 12000 3969
rect 11944 3775 12000 3781
rect 11686 3715 11944 3735
rect 11996 3715 12000 3775
rect 11630 3705 12000 3715
rect 12030 4035 12400 4045
rect 12030 3975 12034 4035
rect 12086 4015 12344 4035
rect 12030 3969 12086 3975
rect 12030 3781 12060 3969
rect 12115 3960 12315 3985
rect 12396 3975 12400 4035
rect 12344 3969 12400 3975
rect 12115 3940 12185 3960
rect 12090 3900 12185 3940
rect 12245 3940 12315 3960
rect 12245 3900 12340 3940
rect 12090 3850 12340 3900
rect 12090 3810 12185 3850
rect 12115 3790 12185 3810
rect 12245 3810 12340 3850
rect 12245 3790 12315 3810
rect 12030 3775 12086 3781
rect 12030 3715 12034 3775
rect 12115 3765 12315 3790
rect 12370 3781 12400 3969
rect 12344 3775 12400 3781
rect 12086 3715 12344 3735
rect 12396 3715 12400 3775
rect 12030 3705 12400 3715
rect 12430 4035 12800 4045
rect 12430 3975 12434 4035
rect 12486 4015 12744 4035
rect 12430 3969 12486 3975
rect 12430 3781 12460 3969
rect 12515 3960 12715 3985
rect 12796 3975 12800 4035
rect 12744 3969 12800 3975
rect 12515 3940 12585 3960
rect 12490 3900 12585 3940
rect 12645 3940 12715 3960
rect 12645 3900 12740 3940
rect 12490 3850 12740 3900
rect 12490 3810 12585 3850
rect 12515 3790 12585 3810
rect 12645 3810 12740 3850
rect 12645 3790 12715 3810
rect 12430 3775 12486 3781
rect 12430 3715 12434 3775
rect 12515 3765 12715 3790
rect 12770 3781 12800 3969
rect 12744 3775 12800 3781
rect 12486 3715 12744 3735
rect 12796 3715 12800 3775
rect 12430 3705 12800 3715
rect 12830 4035 13200 4045
rect 12830 3975 12834 4035
rect 12886 4015 13144 4035
rect 12830 3969 12886 3975
rect 12830 3781 12860 3969
rect 12915 3960 13115 3985
rect 13196 3975 13200 4035
rect 13144 3969 13200 3975
rect 12915 3940 12985 3960
rect 12890 3900 12985 3940
rect 13045 3940 13115 3960
rect 13045 3900 13140 3940
rect 12890 3850 13140 3900
rect 12890 3810 12985 3850
rect 12915 3790 12985 3810
rect 13045 3810 13140 3850
rect 13045 3790 13115 3810
rect 12830 3775 12886 3781
rect 12830 3715 12834 3775
rect 12915 3765 13115 3790
rect 13170 3781 13200 3969
rect 13144 3775 13200 3781
rect 12886 3715 13144 3735
rect 13196 3715 13200 3775
rect 12830 3705 13200 3715
rect -370 3665 0 3675
rect -370 3605 -366 3665
rect -314 3645 -56 3665
rect -370 3599 -314 3605
rect -370 3411 -340 3599
rect -285 3590 -85 3615
rect -4 3605 0 3665
rect -56 3599 0 3605
rect -285 3570 -215 3590
rect -310 3530 -215 3570
rect -155 3570 -85 3590
rect -155 3530 -60 3570
rect -310 3480 -60 3530
rect -310 3440 -215 3480
rect -285 3420 -215 3440
rect -155 3440 -60 3480
rect -155 3420 -85 3440
rect -370 3405 -314 3411
rect -370 3345 -366 3405
rect -285 3395 -85 3420
rect -30 3411 0 3599
rect -56 3405 0 3411
rect -314 3345 -56 3365
rect -4 3345 0 3405
rect -370 3335 0 3345
rect 30 3665 400 3675
rect 30 3605 34 3665
rect 86 3645 344 3665
rect 30 3599 86 3605
rect 30 3411 60 3599
rect 115 3590 315 3615
rect 396 3605 400 3665
rect 344 3599 400 3605
rect 115 3570 185 3590
rect 90 3530 185 3570
rect 245 3570 315 3590
rect 245 3530 340 3570
rect 90 3480 340 3530
rect 90 3440 185 3480
rect 115 3420 185 3440
rect 245 3440 340 3480
rect 245 3420 315 3440
rect 30 3405 86 3411
rect 30 3345 34 3405
rect 115 3395 315 3420
rect 370 3411 400 3599
rect 344 3405 400 3411
rect 86 3345 344 3365
rect 396 3345 400 3405
rect 30 3335 400 3345
rect 430 3665 800 3675
rect 430 3605 434 3665
rect 486 3645 744 3665
rect 430 3599 486 3605
rect 430 3411 460 3599
rect 515 3590 715 3615
rect 796 3605 800 3665
rect 744 3599 800 3605
rect 515 3570 585 3590
rect 490 3530 585 3570
rect 645 3570 715 3590
rect 645 3530 740 3570
rect 490 3480 740 3530
rect 490 3440 585 3480
rect 515 3420 585 3440
rect 645 3440 740 3480
rect 645 3420 715 3440
rect 430 3405 486 3411
rect 430 3345 434 3405
rect 515 3395 715 3420
rect 770 3411 800 3599
rect 744 3405 800 3411
rect 486 3345 744 3365
rect 796 3345 800 3405
rect 430 3335 800 3345
rect 830 3665 1200 3675
rect 830 3605 834 3665
rect 886 3645 1144 3665
rect 830 3599 886 3605
rect 830 3411 860 3599
rect 915 3590 1115 3615
rect 1196 3605 1200 3665
rect 1144 3599 1200 3605
rect 915 3570 985 3590
rect 890 3530 985 3570
rect 1045 3570 1115 3590
rect 1045 3530 1140 3570
rect 890 3480 1140 3530
rect 890 3440 985 3480
rect 915 3420 985 3440
rect 1045 3440 1140 3480
rect 1045 3420 1115 3440
rect 830 3405 886 3411
rect 830 3345 834 3405
rect 915 3395 1115 3420
rect 1170 3411 1200 3599
rect 1144 3405 1200 3411
rect 886 3345 1144 3365
rect 1196 3345 1200 3405
rect 830 3335 1200 3345
rect 1230 3665 1600 3675
rect 1230 3605 1234 3665
rect 1286 3645 1544 3665
rect 1230 3599 1286 3605
rect 1230 3411 1260 3599
rect 1315 3590 1515 3615
rect 1596 3605 1600 3665
rect 1544 3599 1600 3605
rect 1315 3570 1385 3590
rect 1290 3530 1385 3570
rect 1445 3570 1515 3590
rect 1445 3530 1540 3570
rect 1290 3480 1540 3530
rect 1290 3440 1385 3480
rect 1315 3420 1385 3440
rect 1445 3440 1540 3480
rect 1445 3420 1515 3440
rect 1230 3405 1286 3411
rect 1230 3345 1234 3405
rect 1315 3395 1515 3420
rect 1570 3411 1600 3599
rect 1544 3405 1600 3411
rect 1286 3345 1544 3365
rect 1596 3345 1600 3405
rect 1230 3335 1600 3345
rect 1630 3665 2000 3675
rect 1630 3605 1634 3665
rect 1686 3645 1944 3665
rect 1630 3599 1686 3605
rect 1630 3411 1660 3599
rect 1715 3590 1915 3615
rect 1996 3605 2000 3665
rect 1944 3599 2000 3605
rect 1715 3570 1785 3590
rect 1690 3530 1785 3570
rect 1845 3570 1915 3590
rect 1845 3530 1940 3570
rect 1690 3480 1940 3530
rect 1690 3440 1785 3480
rect 1715 3420 1785 3440
rect 1845 3440 1940 3480
rect 1845 3420 1915 3440
rect 1630 3405 1686 3411
rect 1630 3345 1634 3405
rect 1715 3395 1915 3420
rect 1970 3411 2000 3599
rect 1944 3405 2000 3411
rect 1686 3345 1944 3365
rect 1996 3345 2000 3405
rect 1630 3335 2000 3345
rect 2030 3665 2400 3675
rect 2030 3605 2034 3665
rect 2086 3645 2344 3665
rect 2030 3599 2086 3605
rect 2030 3411 2060 3599
rect 2115 3590 2315 3615
rect 2396 3605 2400 3665
rect 2344 3599 2400 3605
rect 2115 3570 2185 3590
rect 2090 3530 2185 3570
rect 2245 3570 2315 3590
rect 2245 3530 2340 3570
rect 2090 3480 2340 3530
rect 2090 3440 2185 3480
rect 2115 3420 2185 3440
rect 2245 3440 2340 3480
rect 2245 3420 2315 3440
rect 2030 3405 2086 3411
rect 2030 3345 2034 3405
rect 2115 3395 2315 3420
rect 2370 3411 2400 3599
rect 2344 3405 2400 3411
rect 2086 3345 2344 3365
rect 2396 3345 2400 3405
rect 2030 3335 2400 3345
rect 2430 3665 2800 3675
rect 2430 3605 2434 3665
rect 2486 3645 2744 3665
rect 2430 3599 2486 3605
rect 2430 3411 2460 3599
rect 2515 3590 2715 3615
rect 2796 3605 2800 3665
rect 2744 3599 2800 3605
rect 2515 3570 2585 3590
rect 2490 3530 2585 3570
rect 2645 3570 2715 3590
rect 2645 3530 2740 3570
rect 2490 3480 2740 3530
rect 2490 3440 2585 3480
rect 2515 3420 2585 3440
rect 2645 3440 2740 3480
rect 2645 3420 2715 3440
rect 2430 3405 2486 3411
rect 2430 3345 2434 3405
rect 2515 3395 2715 3420
rect 2770 3411 2800 3599
rect 2744 3405 2800 3411
rect 2486 3345 2744 3365
rect 2796 3345 2800 3405
rect 2430 3335 2800 3345
rect 2830 3665 3200 3675
rect 2830 3605 2834 3665
rect 2886 3645 3144 3665
rect 2830 3599 2886 3605
rect 2830 3411 2860 3599
rect 2915 3590 3115 3615
rect 3196 3605 3200 3665
rect 3144 3599 3200 3605
rect 2915 3570 2985 3590
rect 2890 3530 2985 3570
rect 3045 3570 3115 3590
rect 3045 3530 3140 3570
rect 2890 3480 3140 3530
rect 2890 3440 2985 3480
rect 2915 3420 2985 3440
rect 3045 3440 3140 3480
rect 3045 3420 3115 3440
rect 2830 3405 2886 3411
rect 2830 3345 2834 3405
rect 2915 3395 3115 3420
rect 3170 3411 3200 3599
rect 3144 3405 3200 3411
rect 2886 3345 3144 3365
rect 3196 3345 3200 3405
rect 2830 3335 3200 3345
rect 3230 3665 3600 3675
rect 3230 3605 3234 3665
rect 3286 3645 3544 3665
rect 3230 3599 3286 3605
rect 3230 3411 3260 3599
rect 3315 3590 3515 3615
rect 3596 3605 3600 3665
rect 3544 3599 3600 3605
rect 3315 3570 3385 3590
rect 3290 3530 3385 3570
rect 3445 3570 3515 3590
rect 3445 3530 3540 3570
rect 3290 3480 3540 3530
rect 3290 3440 3385 3480
rect 3315 3420 3385 3440
rect 3445 3440 3540 3480
rect 3445 3420 3515 3440
rect 3230 3405 3286 3411
rect 3230 3345 3234 3405
rect 3315 3395 3515 3420
rect 3570 3411 3600 3599
rect 3544 3405 3600 3411
rect 3286 3345 3544 3365
rect 3596 3345 3600 3405
rect 3230 3335 3600 3345
rect 3630 3665 4000 3675
rect 3630 3605 3634 3665
rect 3686 3645 3944 3665
rect 3630 3599 3686 3605
rect 3630 3411 3660 3599
rect 3715 3590 3915 3615
rect 3996 3605 4000 3665
rect 3944 3599 4000 3605
rect 3715 3570 3785 3590
rect 3690 3530 3785 3570
rect 3845 3570 3915 3590
rect 3845 3530 3940 3570
rect 3690 3480 3940 3530
rect 3690 3440 3785 3480
rect 3715 3420 3785 3440
rect 3845 3440 3940 3480
rect 3845 3420 3915 3440
rect 3630 3405 3686 3411
rect 3630 3345 3634 3405
rect 3715 3395 3915 3420
rect 3970 3411 4000 3599
rect 3944 3405 4000 3411
rect 3686 3345 3944 3365
rect 3996 3345 4000 3405
rect 3630 3335 4000 3345
rect 4030 3665 4400 3675
rect 4030 3605 4034 3665
rect 4086 3645 4344 3665
rect 4030 3599 4086 3605
rect 4030 3411 4060 3599
rect 4115 3590 4315 3615
rect 4396 3605 4400 3665
rect 4344 3599 4400 3605
rect 4115 3570 4185 3590
rect 4090 3530 4185 3570
rect 4245 3570 4315 3590
rect 4245 3530 4340 3570
rect 4090 3480 4340 3530
rect 4090 3440 4185 3480
rect 4115 3420 4185 3440
rect 4245 3440 4340 3480
rect 4245 3420 4315 3440
rect 4030 3405 4086 3411
rect 4030 3345 4034 3405
rect 4115 3395 4315 3420
rect 4370 3411 4400 3599
rect 4344 3405 4400 3411
rect 4086 3345 4344 3365
rect 4396 3345 4400 3405
rect 4030 3335 4400 3345
rect 4430 3665 4800 3675
rect 4430 3605 4434 3665
rect 4486 3645 4744 3665
rect 4430 3599 4486 3605
rect 4430 3411 4460 3599
rect 4515 3590 4715 3615
rect 4796 3605 4800 3665
rect 4744 3599 4800 3605
rect 4515 3570 4585 3590
rect 4490 3530 4585 3570
rect 4645 3570 4715 3590
rect 4645 3530 4740 3570
rect 4490 3480 4740 3530
rect 4490 3440 4585 3480
rect 4515 3420 4585 3440
rect 4645 3440 4740 3480
rect 4645 3420 4715 3440
rect 4430 3405 4486 3411
rect 4430 3345 4434 3405
rect 4515 3395 4715 3420
rect 4770 3411 4800 3599
rect 4744 3405 4800 3411
rect 4486 3345 4744 3365
rect 4796 3345 4800 3405
rect 4430 3335 4800 3345
rect 4830 3665 5200 3675
rect 4830 3605 4834 3665
rect 4886 3645 5144 3665
rect 4830 3599 4886 3605
rect 4830 3411 4860 3599
rect 4915 3590 5115 3615
rect 5196 3605 5200 3665
rect 5144 3599 5200 3605
rect 4915 3570 4985 3590
rect 4890 3530 4985 3570
rect 5045 3570 5115 3590
rect 5045 3530 5140 3570
rect 4890 3480 5140 3530
rect 4890 3440 4985 3480
rect 4915 3420 4985 3440
rect 5045 3440 5140 3480
rect 5045 3420 5115 3440
rect 4830 3405 4886 3411
rect 4830 3345 4834 3405
rect 4915 3395 5115 3420
rect 5170 3411 5200 3599
rect 5144 3405 5200 3411
rect 4886 3345 5144 3365
rect 5196 3345 5200 3405
rect 4830 3335 5200 3345
rect 5230 3665 5600 3675
rect 5230 3605 5234 3665
rect 5286 3645 5544 3665
rect 5230 3599 5286 3605
rect 5230 3411 5260 3599
rect 5315 3590 5515 3615
rect 5596 3605 5600 3665
rect 5544 3599 5600 3605
rect 5315 3570 5385 3590
rect 5290 3530 5385 3570
rect 5445 3570 5515 3590
rect 5445 3530 5540 3570
rect 5290 3480 5540 3530
rect 5290 3440 5385 3480
rect 5315 3420 5385 3440
rect 5445 3440 5540 3480
rect 5445 3420 5515 3440
rect 5230 3405 5286 3411
rect 5230 3345 5234 3405
rect 5315 3395 5515 3420
rect 5570 3411 5600 3599
rect 5544 3405 5600 3411
rect 5286 3345 5544 3365
rect 5596 3345 5600 3405
rect 5230 3335 5600 3345
rect 5630 3665 6000 3675
rect 5630 3605 5634 3665
rect 5686 3645 5944 3665
rect 5630 3599 5686 3605
rect 5630 3411 5660 3599
rect 5715 3590 5915 3615
rect 5996 3605 6000 3665
rect 5944 3599 6000 3605
rect 5715 3570 5785 3590
rect 5690 3530 5785 3570
rect 5845 3570 5915 3590
rect 5845 3530 5940 3570
rect 5690 3480 5940 3530
rect 5690 3440 5785 3480
rect 5715 3420 5785 3440
rect 5845 3440 5940 3480
rect 5845 3420 5915 3440
rect 5630 3405 5686 3411
rect 5630 3345 5634 3405
rect 5715 3395 5915 3420
rect 5970 3411 6000 3599
rect 5944 3405 6000 3411
rect 5686 3345 5944 3365
rect 5996 3345 6000 3405
rect 5630 3335 6000 3345
rect 6030 3665 6400 3675
rect 6030 3605 6034 3665
rect 6086 3645 6344 3665
rect 6030 3599 6086 3605
rect 6030 3411 6060 3599
rect 6115 3590 6315 3615
rect 6396 3605 6400 3665
rect 6344 3599 6400 3605
rect 6115 3570 6185 3590
rect 6090 3530 6185 3570
rect 6245 3570 6315 3590
rect 6245 3530 6340 3570
rect 6090 3480 6340 3530
rect 6090 3440 6185 3480
rect 6115 3420 6185 3440
rect 6245 3440 6340 3480
rect 6245 3420 6315 3440
rect 6030 3405 6086 3411
rect 6030 3345 6034 3405
rect 6115 3395 6315 3420
rect 6370 3411 6400 3599
rect 6344 3405 6400 3411
rect 6086 3345 6344 3365
rect 6396 3345 6400 3405
rect 6030 3335 6400 3345
rect 6430 3665 6800 3675
rect 6430 3605 6434 3665
rect 6486 3645 6744 3665
rect 6430 3599 6486 3605
rect 6430 3411 6460 3599
rect 6515 3590 6715 3615
rect 6796 3605 6800 3665
rect 6744 3599 6800 3605
rect 6515 3570 6585 3590
rect 6490 3530 6585 3570
rect 6645 3570 6715 3590
rect 6645 3530 6740 3570
rect 6490 3480 6740 3530
rect 6490 3440 6585 3480
rect 6515 3420 6585 3440
rect 6645 3440 6740 3480
rect 6645 3420 6715 3440
rect 6430 3405 6486 3411
rect 6430 3345 6434 3405
rect 6515 3395 6715 3420
rect 6770 3411 6800 3599
rect 6744 3405 6800 3411
rect 6486 3345 6744 3365
rect 6796 3345 6800 3405
rect 6430 3335 6800 3345
rect 6830 3665 7200 3675
rect 6830 3605 6834 3665
rect 6886 3645 7144 3665
rect 6830 3599 6886 3605
rect 6830 3411 6860 3599
rect 6915 3590 7115 3615
rect 7196 3605 7200 3665
rect 7144 3599 7200 3605
rect 6915 3570 6985 3590
rect 6890 3530 6985 3570
rect 7045 3570 7115 3590
rect 7045 3530 7140 3570
rect 6890 3480 7140 3530
rect 6890 3440 6985 3480
rect 6915 3420 6985 3440
rect 7045 3440 7140 3480
rect 7045 3420 7115 3440
rect 6830 3405 6886 3411
rect 6830 3345 6834 3405
rect 6915 3395 7115 3420
rect 7170 3411 7200 3599
rect 7144 3405 7200 3411
rect 6886 3345 7144 3365
rect 7196 3345 7200 3405
rect 6830 3335 7200 3345
rect 7230 3665 7600 3675
rect 7230 3605 7234 3665
rect 7286 3645 7544 3665
rect 7230 3599 7286 3605
rect 7230 3411 7260 3599
rect 7315 3590 7515 3615
rect 7596 3605 7600 3665
rect 7544 3599 7600 3605
rect 7315 3570 7385 3590
rect 7290 3530 7385 3570
rect 7445 3570 7515 3590
rect 7445 3530 7540 3570
rect 7290 3480 7540 3530
rect 7290 3440 7385 3480
rect 7315 3420 7385 3440
rect 7445 3440 7540 3480
rect 7445 3420 7515 3440
rect 7230 3405 7286 3411
rect 7230 3345 7234 3405
rect 7315 3395 7515 3420
rect 7570 3411 7600 3599
rect 7544 3405 7600 3411
rect 7286 3345 7544 3365
rect 7596 3345 7600 3405
rect 7230 3335 7600 3345
rect 7630 3665 8000 3675
rect 7630 3605 7634 3665
rect 7686 3645 7944 3665
rect 7630 3599 7686 3605
rect 7630 3411 7660 3599
rect 7715 3590 7915 3615
rect 7996 3605 8000 3665
rect 7944 3599 8000 3605
rect 7715 3570 7785 3590
rect 7690 3530 7785 3570
rect 7845 3570 7915 3590
rect 7845 3530 7940 3570
rect 7690 3480 7940 3530
rect 7690 3440 7785 3480
rect 7715 3420 7785 3440
rect 7845 3440 7940 3480
rect 7845 3420 7915 3440
rect 7630 3405 7686 3411
rect 7630 3345 7634 3405
rect 7715 3395 7915 3420
rect 7970 3411 8000 3599
rect 7944 3405 8000 3411
rect 7686 3345 7944 3365
rect 7996 3345 8000 3405
rect 7630 3335 8000 3345
rect 8030 3665 8400 3675
rect 8030 3605 8034 3665
rect 8086 3645 8344 3665
rect 8030 3599 8086 3605
rect 8030 3411 8060 3599
rect 8115 3590 8315 3615
rect 8396 3605 8400 3665
rect 8344 3599 8400 3605
rect 8115 3570 8185 3590
rect 8090 3530 8185 3570
rect 8245 3570 8315 3590
rect 8245 3530 8340 3570
rect 8090 3480 8340 3530
rect 8090 3440 8185 3480
rect 8115 3420 8185 3440
rect 8245 3440 8340 3480
rect 8245 3420 8315 3440
rect 8030 3405 8086 3411
rect 8030 3345 8034 3405
rect 8115 3395 8315 3420
rect 8370 3411 8400 3599
rect 8344 3405 8400 3411
rect 8086 3345 8344 3365
rect 8396 3345 8400 3405
rect 8030 3335 8400 3345
rect 8430 3665 8800 3675
rect 8430 3605 8434 3665
rect 8486 3645 8744 3665
rect 8430 3599 8486 3605
rect 8430 3411 8460 3599
rect 8515 3590 8715 3615
rect 8796 3605 8800 3665
rect 8744 3599 8800 3605
rect 8515 3570 8585 3590
rect 8490 3530 8585 3570
rect 8645 3570 8715 3590
rect 8645 3530 8740 3570
rect 8490 3480 8740 3530
rect 8490 3440 8585 3480
rect 8515 3420 8585 3440
rect 8645 3440 8740 3480
rect 8645 3420 8715 3440
rect 8430 3405 8486 3411
rect 8430 3345 8434 3405
rect 8515 3395 8715 3420
rect 8770 3411 8800 3599
rect 8744 3405 8800 3411
rect 8486 3345 8744 3365
rect 8796 3345 8800 3405
rect 8430 3335 8800 3345
rect 8830 3665 9200 3675
rect 8830 3605 8834 3665
rect 8886 3645 9144 3665
rect 8830 3599 8886 3605
rect 8830 3411 8860 3599
rect 8915 3590 9115 3615
rect 9196 3605 9200 3665
rect 9144 3599 9200 3605
rect 8915 3570 8985 3590
rect 8890 3530 8985 3570
rect 9045 3570 9115 3590
rect 9045 3530 9140 3570
rect 8890 3480 9140 3530
rect 8890 3440 8985 3480
rect 8915 3420 8985 3440
rect 9045 3440 9140 3480
rect 9045 3420 9115 3440
rect 8830 3405 8886 3411
rect 8830 3345 8834 3405
rect 8915 3395 9115 3420
rect 9170 3411 9200 3599
rect 9144 3405 9200 3411
rect 8886 3345 9144 3365
rect 9196 3345 9200 3405
rect 8830 3335 9200 3345
rect 9230 3665 9600 3675
rect 9230 3605 9234 3665
rect 9286 3645 9544 3665
rect 9230 3599 9286 3605
rect 9230 3411 9260 3599
rect 9315 3590 9515 3615
rect 9596 3605 9600 3665
rect 9544 3599 9600 3605
rect 9315 3570 9385 3590
rect 9290 3530 9385 3570
rect 9445 3570 9515 3590
rect 9445 3530 9540 3570
rect 9290 3480 9540 3530
rect 9290 3440 9385 3480
rect 9315 3420 9385 3440
rect 9445 3440 9540 3480
rect 9445 3420 9515 3440
rect 9230 3405 9286 3411
rect 9230 3345 9234 3405
rect 9315 3395 9515 3420
rect 9570 3411 9600 3599
rect 9544 3405 9600 3411
rect 9286 3345 9544 3365
rect 9596 3345 9600 3405
rect 9230 3335 9600 3345
rect 9630 3665 10000 3675
rect 9630 3605 9634 3665
rect 9686 3645 9944 3665
rect 9630 3599 9686 3605
rect 9630 3411 9660 3599
rect 9715 3590 9915 3615
rect 9996 3605 10000 3665
rect 9944 3599 10000 3605
rect 9715 3570 9785 3590
rect 9690 3530 9785 3570
rect 9845 3570 9915 3590
rect 9845 3530 9940 3570
rect 9690 3480 9940 3530
rect 9690 3440 9785 3480
rect 9715 3420 9785 3440
rect 9845 3440 9940 3480
rect 9845 3420 9915 3440
rect 9630 3405 9686 3411
rect 9630 3345 9634 3405
rect 9715 3395 9915 3420
rect 9970 3411 10000 3599
rect 9944 3405 10000 3411
rect 9686 3345 9944 3365
rect 9996 3345 10000 3405
rect 9630 3335 10000 3345
rect 10030 3665 10400 3675
rect 10030 3605 10034 3665
rect 10086 3645 10344 3665
rect 10030 3599 10086 3605
rect 10030 3411 10060 3599
rect 10115 3590 10315 3615
rect 10396 3605 10400 3665
rect 10344 3599 10400 3605
rect 10115 3570 10185 3590
rect 10090 3530 10185 3570
rect 10245 3570 10315 3590
rect 10245 3530 10340 3570
rect 10090 3480 10340 3530
rect 10090 3440 10185 3480
rect 10115 3420 10185 3440
rect 10245 3440 10340 3480
rect 10245 3420 10315 3440
rect 10030 3405 10086 3411
rect 10030 3345 10034 3405
rect 10115 3395 10315 3420
rect 10370 3411 10400 3599
rect 10344 3405 10400 3411
rect 10086 3345 10344 3365
rect 10396 3345 10400 3405
rect 10030 3335 10400 3345
rect 10430 3665 10800 3675
rect 10430 3605 10434 3665
rect 10486 3645 10744 3665
rect 10430 3599 10486 3605
rect 10430 3411 10460 3599
rect 10515 3590 10715 3615
rect 10796 3605 10800 3665
rect 10744 3599 10800 3605
rect 10515 3570 10585 3590
rect 10490 3530 10585 3570
rect 10645 3570 10715 3590
rect 10645 3530 10740 3570
rect 10490 3480 10740 3530
rect 10490 3440 10585 3480
rect 10515 3420 10585 3440
rect 10645 3440 10740 3480
rect 10645 3420 10715 3440
rect 10430 3405 10486 3411
rect 10430 3345 10434 3405
rect 10515 3395 10715 3420
rect 10770 3411 10800 3599
rect 10744 3405 10800 3411
rect 10486 3345 10744 3365
rect 10796 3345 10800 3405
rect 10430 3335 10800 3345
rect 10830 3665 11200 3675
rect 10830 3605 10834 3665
rect 10886 3645 11144 3665
rect 10830 3599 10886 3605
rect 10830 3411 10860 3599
rect 10915 3590 11115 3615
rect 11196 3605 11200 3665
rect 11144 3599 11200 3605
rect 10915 3570 10985 3590
rect 10890 3530 10985 3570
rect 11045 3570 11115 3590
rect 11045 3530 11140 3570
rect 10890 3480 11140 3530
rect 10890 3440 10985 3480
rect 10915 3420 10985 3440
rect 11045 3440 11140 3480
rect 11045 3420 11115 3440
rect 10830 3405 10886 3411
rect 10830 3345 10834 3405
rect 10915 3395 11115 3420
rect 11170 3411 11200 3599
rect 11144 3405 11200 3411
rect 10886 3345 11144 3365
rect 11196 3345 11200 3405
rect 10830 3335 11200 3345
rect 11230 3665 11600 3675
rect 11230 3605 11234 3665
rect 11286 3645 11544 3665
rect 11230 3599 11286 3605
rect 11230 3411 11260 3599
rect 11315 3590 11515 3615
rect 11596 3605 11600 3665
rect 11544 3599 11600 3605
rect 11315 3570 11385 3590
rect 11290 3530 11385 3570
rect 11445 3570 11515 3590
rect 11445 3530 11540 3570
rect 11290 3480 11540 3530
rect 11290 3440 11385 3480
rect 11315 3420 11385 3440
rect 11445 3440 11540 3480
rect 11445 3420 11515 3440
rect 11230 3405 11286 3411
rect 11230 3345 11234 3405
rect 11315 3395 11515 3420
rect 11570 3411 11600 3599
rect 11544 3405 11600 3411
rect 11286 3345 11544 3365
rect 11596 3345 11600 3405
rect 11230 3335 11600 3345
rect 11630 3665 12000 3675
rect 11630 3605 11634 3665
rect 11686 3645 11944 3665
rect 11630 3599 11686 3605
rect 11630 3411 11660 3599
rect 11715 3590 11915 3615
rect 11996 3605 12000 3665
rect 11944 3599 12000 3605
rect 11715 3570 11785 3590
rect 11690 3530 11785 3570
rect 11845 3570 11915 3590
rect 11845 3530 11940 3570
rect 11690 3480 11940 3530
rect 11690 3440 11785 3480
rect 11715 3420 11785 3440
rect 11845 3440 11940 3480
rect 11845 3420 11915 3440
rect 11630 3405 11686 3411
rect 11630 3345 11634 3405
rect 11715 3395 11915 3420
rect 11970 3411 12000 3599
rect 11944 3405 12000 3411
rect 11686 3345 11944 3365
rect 11996 3345 12000 3405
rect 11630 3335 12000 3345
rect 12030 3665 12400 3675
rect 12030 3605 12034 3665
rect 12086 3645 12344 3665
rect 12030 3599 12086 3605
rect 12030 3411 12060 3599
rect 12115 3590 12315 3615
rect 12396 3605 12400 3665
rect 12344 3599 12400 3605
rect 12115 3570 12185 3590
rect 12090 3530 12185 3570
rect 12245 3570 12315 3590
rect 12245 3530 12340 3570
rect 12090 3480 12340 3530
rect 12090 3440 12185 3480
rect 12115 3420 12185 3440
rect 12245 3440 12340 3480
rect 12245 3420 12315 3440
rect 12030 3405 12086 3411
rect 12030 3345 12034 3405
rect 12115 3395 12315 3420
rect 12370 3411 12400 3599
rect 12344 3405 12400 3411
rect 12086 3345 12344 3365
rect 12396 3345 12400 3405
rect 12030 3335 12400 3345
rect 12430 3665 12800 3675
rect 12430 3605 12434 3665
rect 12486 3645 12744 3665
rect 12430 3599 12486 3605
rect 12430 3411 12460 3599
rect 12515 3590 12715 3615
rect 12796 3605 12800 3665
rect 12744 3599 12800 3605
rect 12515 3570 12585 3590
rect 12490 3530 12585 3570
rect 12645 3570 12715 3590
rect 12645 3530 12740 3570
rect 12490 3480 12740 3530
rect 12490 3440 12585 3480
rect 12515 3420 12585 3440
rect 12645 3440 12740 3480
rect 12645 3420 12715 3440
rect 12430 3405 12486 3411
rect 12430 3345 12434 3405
rect 12515 3395 12715 3420
rect 12770 3411 12800 3599
rect 12744 3405 12800 3411
rect 12486 3345 12744 3365
rect 12796 3345 12800 3405
rect 12430 3335 12800 3345
rect 12830 3665 13200 3675
rect 12830 3605 12834 3665
rect 12886 3645 13144 3665
rect 12830 3599 12886 3605
rect 12830 3411 12860 3599
rect 12915 3590 13115 3615
rect 13196 3605 13200 3665
rect 13144 3599 13200 3605
rect 12915 3570 12985 3590
rect 12890 3530 12985 3570
rect 13045 3570 13115 3590
rect 13045 3530 13140 3570
rect 12890 3480 13140 3530
rect 12890 3440 12985 3480
rect 12915 3420 12985 3440
rect 13045 3440 13140 3480
rect 13045 3420 13115 3440
rect 12830 3405 12886 3411
rect 12830 3345 12834 3405
rect 12915 3395 13115 3420
rect 13170 3411 13200 3599
rect 13144 3405 13200 3411
rect 12886 3345 13144 3365
rect 13196 3345 13200 3405
rect 12830 3335 13200 3345
rect -370 3295 0 3305
rect -370 3235 -366 3295
rect -314 3275 -56 3295
rect -370 3229 -314 3235
rect -370 3041 -340 3229
rect -285 3220 -85 3245
rect -4 3235 0 3295
rect -56 3229 0 3235
rect -285 3200 -215 3220
rect -310 3160 -215 3200
rect -155 3200 -85 3220
rect -155 3160 -60 3200
rect -310 3110 -60 3160
rect -310 3070 -215 3110
rect -285 3050 -215 3070
rect -155 3070 -60 3110
rect -155 3050 -85 3070
rect -370 3035 -314 3041
rect -370 2975 -366 3035
rect -285 3025 -85 3050
rect -30 3041 0 3229
rect -56 3035 0 3041
rect -314 2975 -56 2995
rect -4 2975 0 3035
rect -370 2965 0 2975
rect 30 3295 400 3305
rect 30 3235 34 3295
rect 86 3275 344 3295
rect 30 3229 86 3235
rect 30 3041 60 3229
rect 115 3220 315 3245
rect 396 3235 400 3295
rect 344 3229 400 3235
rect 115 3200 185 3220
rect 90 3160 185 3200
rect 245 3200 315 3220
rect 245 3160 340 3200
rect 90 3110 340 3160
rect 90 3070 185 3110
rect 115 3050 185 3070
rect 245 3070 340 3110
rect 245 3050 315 3070
rect 30 3035 86 3041
rect 30 2975 34 3035
rect 115 3025 315 3050
rect 370 3041 400 3229
rect 344 3035 400 3041
rect 86 2975 344 2995
rect 396 2975 400 3035
rect 30 2965 400 2975
rect 430 3295 800 3305
rect 430 3235 434 3295
rect 486 3275 744 3295
rect 430 3229 486 3235
rect 430 3041 460 3229
rect 515 3220 715 3245
rect 796 3235 800 3295
rect 744 3229 800 3235
rect 515 3200 585 3220
rect 490 3160 585 3200
rect 645 3200 715 3220
rect 645 3160 740 3200
rect 490 3110 740 3160
rect 490 3070 585 3110
rect 515 3050 585 3070
rect 645 3070 740 3110
rect 645 3050 715 3070
rect 430 3035 486 3041
rect 430 2975 434 3035
rect 515 3025 715 3050
rect 770 3041 800 3229
rect 744 3035 800 3041
rect 486 2975 744 2995
rect 796 2975 800 3035
rect 430 2965 800 2975
rect 830 3295 1200 3305
rect 830 3235 834 3295
rect 886 3275 1144 3295
rect 830 3229 886 3235
rect 830 3041 860 3229
rect 915 3220 1115 3245
rect 1196 3235 1200 3295
rect 1144 3229 1200 3235
rect 915 3200 985 3220
rect 890 3160 985 3200
rect 1045 3200 1115 3220
rect 1045 3160 1140 3200
rect 890 3110 1140 3160
rect 890 3070 985 3110
rect 915 3050 985 3070
rect 1045 3070 1140 3110
rect 1045 3050 1115 3070
rect 830 3035 886 3041
rect 830 2975 834 3035
rect 915 3025 1115 3050
rect 1170 3041 1200 3229
rect 1144 3035 1200 3041
rect 886 2975 1144 2995
rect 1196 2975 1200 3035
rect 830 2965 1200 2975
rect 1230 3295 1600 3305
rect 1230 3235 1234 3295
rect 1286 3275 1544 3295
rect 1230 3229 1286 3235
rect 1230 3041 1260 3229
rect 1315 3220 1515 3245
rect 1596 3235 1600 3295
rect 1544 3229 1600 3235
rect 1315 3200 1385 3220
rect 1290 3160 1385 3200
rect 1445 3200 1515 3220
rect 1445 3160 1540 3200
rect 1290 3110 1540 3160
rect 1290 3070 1385 3110
rect 1315 3050 1385 3070
rect 1445 3070 1540 3110
rect 1445 3050 1515 3070
rect 1230 3035 1286 3041
rect 1230 2975 1234 3035
rect 1315 3025 1515 3050
rect 1570 3041 1600 3229
rect 1544 3035 1600 3041
rect 1286 2975 1544 2995
rect 1596 2975 1600 3035
rect 1230 2965 1600 2975
rect 1630 3295 2000 3305
rect 1630 3235 1634 3295
rect 1686 3275 1944 3295
rect 1630 3229 1686 3235
rect 1630 3041 1660 3229
rect 1715 3220 1915 3245
rect 1996 3235 2000 3295
rect 1944 3229 2000 3235
rect 1715 3200 1785 3220
rect 1690 3160 1785 3200
rect 1845 3200 1915 3220
rect 1845 3160 1940 3200
rect 1690 3110 1940 3160
rect 1690 3070 1785 3110
rect 1715 3050 1785 3070
rect 1845 3070 1940 3110
rect 1845 3050 1915 3070
rect 1630 3035 1686 3041
rect 1630 2975 1634 3035
rect 1715 3025 1915 3050
rect 1970 3041 2000 3229
rect 1944 3035 2000 3041
rect 1686 2975 1944 2995
rect 1996 2975 2000 3035
rect 1630 2965 2000 2975
rect 2030 3295 2400 3305
rect 2030 3235 2034 3295
rect 2086 3275 2344 3295
rect 2030 3229 2086 3235
rect 2030 3041 2060 3229
rect 2115 3220 2315 3245
rect 2396 3235 2400 3295
rect 2344 3229 2400 3235
rect 2115 3200 2185 3220
rect 2090 3160 2185 3200
rect 2245 3200 2315 3220
rect 2245 3160 2340 3200
rect 2090 3110 2340 3160
rect 2090 3070 2185 3110
rect 2115 3050 2185 3070
rect 2245 3070 2340 3110
rect 2245 3050 2315 3070
rect 2030 3035 2086 3041
rect 2030 2975 2034 3035
rect 2115 3025 2315 3050
rect 2370 3041 2400 3229
rect 2344 3035 2400 3041
rect 2086 2975 2344 2995
rect 2396 2975 2400 3035
rect 2030 2965 2400 2975
rect 2430 3295 2800 3305
rect 2430 3235 2434 3295
rect 2486 3275 2744 3295
rect 2430 3229 2486 3235
rect 2430 3041 2460 3229
rect 2515 3220 2715 3245
rect 2796 3235 2800 3295
rect 2744 3229 2800 3235
rect 2515 3200 2585 3220
rect 2490 3160 2585 3200
rect 2645 3200 2715 3220
rect 2645 3160 2740 3200
rect 2490 3110 2740 3160
rect 2490 3070 2585 3110
rect 2515 3050 2585 3070
rect 2645 3070 2740 3110
rect 2645 3050 2715 3070
rect 2430 3035 2486 3041
rect 2430 2975 2434 3035
rect 2515 3025 2715 3050
rect 2770 3041 2800 3229
rect 2744 3035 2800 3041
rect 2486 2975 2744 2995
rect 2796 2975 2800 3035
rect 2430 2965 2800 2975
rect 2830 3295 3200 3305
rect 2830 3235 2834 3295
rect 2886 3275 3144 3295
rect 2830 3229 2886 3235
rect 2830 3041 2860 3229
rect 2915 3220 3115 3245
rect 3196 3235 3200 3295
rect 3144 3229 3200 3235
rect 2915 3200 2985 3220
rect 2890 3160 2985 3200
rect 3045 3200 3115 3220
rect 3045 3160 3140 3200
rect 2890 3110 3140 3160
rect 2890 3070 2985 3110
rect 2915 3050 2985 3070
rect 3045 3070 3140 3110
rect 3045 3050 3115 3070
rect 2830 3035 2886 3041
rect 2830 2975 2834 3035
rect 2915 3025 3115 3050
rect 3170 3041 3200 3229
rect 3144 3035 3200 3041
rect 2886 2975 3144 2995
rect 3196 2975 3200 3035
rect 2830 2965 3200 2975
rect 3230 3295 3600 3305
rect 3230 3235 3234 3295
rect 3286 3275 3544 3295
rect 3230 3229 3286 3235
rect 3230 3041 3260 3229
rect 3315 3220 3515 3245
rect 3596 3235 3600 3295
rect 3544 3229 3600 3235
rect 3315 3200 3385 3220
rect 3290 3160 3385 3200
rect 3445 3200 3515 3220
rect 3445 3160 3540 3200
rect 3290 3110 3540 3160
rect 3290 3070 3385 3110
rect 3315 3050 3385 3070
rect 3445 3070 3540 3110
rect 3445 3050 3515 3070
rect 3230 3035 3286 3041
rect 3230 2975 3234 3035
rect 3315 3025 3515 3050
rect 3570 3041 3600 3229
rect 3544 3035 3600 3041
rect 3286 2975 3544 2995
rect 3596 2975 3600 3035
rect 3230 2965 3600 2975
rect 3630 3295 4000 3305
rect 3630 3235 3634 3295
rect 3686 3275 3944 3295
rect 3630 3229 3686 3235
rect 3630 3041 3660 3229
rect 3715 3220 3915 3245
rect 3996 3235 4000 3295
rect 3944 3229 4000 3235
rect 3715 3200 3785 3220
rect 3690 3160 3785 3200
rect 3845 3200 3915 3220
rect 3845 3160 3940 3200
rect 3690 3110 3940 3160
rect 3690 3070 3785 3110
rect 3715 3050 3785 3070
rect 3845 3070 3940 3110
rect 3845 3050 3915 3070
rect 3630 3035 3686 3041
rect 3630 2975 3634 3035
rect 3715 3025 3915 3050
rect 3970 3041 4000 3229
rect 3944 3035 4000 3041
rect 3686 2975 3944 2995
rect 3996 2975 4000 3035
rect 3630 2965 4000 2975
rect 4030 3295 4400 3305
rect 4030 3235 4034 3295
rect 4086 3275 4344 3295
rect 4030 3229 4086 3235
rect 4030 3041 4060 3229
rect 4115 3220 4315 3245
rect 4396 3235 4400 3295
rect 4344 3229 4400 3235
rect 4115 3200 4185 3220
rect 4090 3160 4185 3200
rect 4245 3200 4315 3220
rect 4245 3160 4340 3200
rect 4090 3110 4340 3160
rect 4090 3070 4185 3110
rect 4115 3050 4185 3070
rect 4245 3070 4340 3110
rect 4245 3050 4315 3070
rect 4030 3035 4086 3041
rect 4030 2975 4034 3035
rect 4115 3025 4315 3050
rect 4370 3041 4400 3229
rect 4344 3035 4400 3041
rect 4086 2975 4344 2995
rect 4396 2975 4400 3035
rect 4030 2965 4400 2975
rect 4430 3295 4800 3305
rect 4430 3235 4434 3295
rect 4486 3275 4744 3295
rect 4430 3229 4486 3235
rect 4430 3041 4460 3229
rect 4515 3220 4715 3245
rect 4796 3235 4800 3295
rect 4744 3229 4800 3235
rect 4515 3200 4585 3220
rect 4490 3160 4585 3200
rect 4645 3200 4715 3220
rect 4645 3160 4740 3200
rect 4490 3110 4740 3160
rect 4490 3070 4585 3110
rect 4515 3050 4585 3070
rect 4645 3070 4740 3110
rect 4645 3050 4715 3070
rect 4430 3035 4486 3041
rect 4430 2975 4434 3035
rect 4515 3025 4715 3050
rect 4770 3041 4800 3229
rect 4744 3035 4800 3041
rect 4486 2975 4744 2995
rect 4796 2975 4800 3035
rect 4430 2965 4800 2975
rect 4830 3295 5200 3305
rect 4830 3235 4834 3295
rect 4886 3275 5144 3295
rect 4830 3229 4886 3235
rect 4830 3041 4860 3229
rect 4915 3220 5115 3245
rect 5196 3235 5200 3295
rect 5144 3229 5200 3235
rect 4915 3200 4985 3220
rect 4890 3160 4985 3200
rect 5045 3200 5115 3220
rect 5045 3160 5140 3200
rect 4890 3110 5140 3160
rect 4890 3070 4985 3110
rect 4915 3050 4985 3070
rect 5045 3070 5140 3110
rect 5045 3050 5115 3070
rect 4830 3035 4886 3041
rect 4830 2975 4834 3035
rect 4915 3025 5115 3050
rect 5170 3041 5200 3229
rect 5144 3035 5200 3041
rect 4886 2975 5144 2995
rect 5196 2975 5200 3035
rect 4830 2965 5200 2975
rect 5230 3295 5600 3305
rect 5230 3235 5234 3295
rect 5286 3275 5544 3295
rect 5230 3229 5286 3235
rect 5230 3041 5260 3229
rect 5315 3220 5515 3245
rect 5596 3235 5600 3295
rect 5544 3229 5600 3235
rect 5315 3200 5385 3220
rect 5290 3160 5385 3200
rect 5445 3200 5515 3220
rect 5445 3160 5540 3200
rect 5290 3110 5540 3160
rect 5290 3070 5385 3110
rect 5315 3050 5385 3070
rect 5445 3070 5540 3110
rect 5445 3050 5515 3070
rect 5230 3035 5286 3041
rect 5230 2975 5234 3035
rect 5315 3025 5515 3050
rect 5570 3041 5600 3229
rect 5544 3035 5600 3041
rect 5286 2975 5544 2995
rect 5596 2975 5600 3035
rect 5230 2965 5600 2975
rect 5630 3295 6000 3305
rect 5630 3235 5634 3295
rect 5686 3275 5944 3295
rect 5630 3229 5686 3235
rect 5630 3041 5660 3229
rect 5715 3220 5915 3245
rect 5996 3235 6000 3295
rect 5944 3229 6000 3235
rect 5715 3200 5785 3220
rect 5690 3160 5785 3200
rect 5845 3200 5915 3220
rect 5845 3160 5940 3200
rect 5690 3110 5940 3160
rect 5690 3070 5785 3110
rect 5715 3050 5785 3070
rect 5845 3070 5940 3110
rect 5845 3050 5915 3070
rect 5630 3035 5686 3041
rect 5630 2975 5634 3035
rect 5715 3025 5915 3050
rect 5970 3041 6000 3229
rect 5944 3035 6000 3041
rect 5686 2975 5944 2995
rect 5996 2975 6000 3035
rect 5630 2965 6000 2975
rect 6030 3295 6400 3305
rect 6030 3235 6034 3295
rect 6086 3275 6344 3295
rect 6030 3229 6086 3235
rect 6030 3041 6060 3229
rect 6115 3220 6315 3245
rect 6396 3235 6400 3295
rect 6344 3229 6400 3235
rect 6115 3200 6185 3220
rect 6090 3160 6185 3200
rect 6245 3200 6315 3220
rect 6245 3160 6340 3200
rect 6090 3110 6340 3160
rect 6090 3070 6185 3110
rect 6115 3050 6185 3070
rect 6245 3070 6340 3110
rect 6245 3050 6315 3070
rect 6030 3035 6086 3041
rect 6030 2975 6034 3035
rect 6115 3025 6315 3050
rect 6370 3041 6400 3229
rect 6344 3035 6400 3041
rect 6086 2975 6344 2995
rect 6396 2975 6400 3035
rect 6030 2965 6400 2975
rect 6430 3295 6800 3305
rect 6430 3235 6434 3295
rect 6486 3275 6744 3295
rect 6430 3229 6486 3235
rect 6430 3041 6460 3229
rect 6515 3220 6715 3245
rect 6796 3235 6800 3295
rect 6744 3229 6800 3235
rect 6515 3200 6585 3220
rect 6490 3160 6585 3200
rect 6645 3200 6715 3220
rect 6645 3160 6740 3200
rect 6490 3110 6740 3160
rect 6490 3070 6585 3110
rect 6515 3050 6585 3070
rect 6645 3070 6740 3110
rect 6645 3050 6715 3070
rect 6430 3035 6486 3041
rect 6430 2975 6434 3035
rect 6515 3025 6715 3050
rect 6770 3041 6800 3229
rect 6744 3035 6800 3041
rect 6486 2975 6744 2995
rect 6796 2975 6800 3035
rect 6430 2965 6800 2975
rect 6830 3295 7200 3305
rect 6830 3235 6834 3295
rect 6886 3275 7144 3295
rect 6830 3229 6886 3235
rect 6830 3041 6860 3229
rect 6915 3220 7115 3245
rect 7196 3235 7200 3295
rect 7144 3229 7200 3235
rect 6915 3200 6985 3220
rect 6890 3160 6985 3200
rect 7045 3200 7115 3220
rect 7045 3160 7140 3200
rect 6890 3110 7140 3160
rect 6890 3070 6985 3110
rect 6915 3050 6985 3070
rect 7045 3070 7140 3110
rect 7045 3050 7115 3070
rect 6830 3035 6886 3041
rect 6830 2975 6834 3035
rect 6915 3025 7115 3050
rect 7170 3041 7200 3229
rect 7144 3035 7200 3041
rect 6886 2975 7144 2995
rect 7196 2975 7200 3035
rect 6830 2965 7200 2975
rect 7230 3295 7600 3305
rect 7230 3235 7234 3295
rect 7286 3275 7544 3295
rect 7230 3229 7286 3235
rect 7230 3041 7260 3229
rect 7315 3220 7515 3245
rect 7596 3235 7600 3295
rect 7544 3229 7600 3235
rect 7315 3200 7385 3220
rect 7290 3160 7385 3200
rect 7445 3200 7515 3220
rect 7445 3160 7540 3200
rect 7290 3110 7540 3160
rect 7290 3070 7385 3110
rect 7315 3050 7385 3070
rect 7445 3070 7540 3110
rect 7445 3050 7515 3070
rect 7230 3035 7286 3041
rect 7230 2975 7234 3035
rect 7315 3025 7515 3050
rect 7570 3041 7600 3229
rect 7544 3035 7600 3041
rect 7286 2975 7544 2995
rect 7596 2975 7600 3035
rect 7230 2965 7600 2975
rect 7630 3295 8000 3305
rect 7630 3235 7634 3295
rect 7686 3275 7944 3295
rect 7630 3229 7686 3235
rect 7630 3041 7660 3229
rect 7715 3220 7915 3245
rect 7996 3235 8000 3295
rect 7944 3229 8000 3235
rect 7715 3200 7785 3220
rect 7690 3160 7785 3200
rect 7845 3200 7915 3220
rect 7845 3160 7940 3200
rect 7690 3110 7940 3160
rect 7690 3070 7785 3110
rect 7715 3050 7785 3070
rect 7845 3070 7940 3110
rect 7845 3050 7915 3070
rect 7630 3035 7686 3041
rect 7630 2975 7634 3035
rect 7715 3025 7915 3050
rect 7970 3041 8000 3229
rect 7944 3035 8000 3041
rect 7686 2975 7944 2995
rect 7996 2975 8000 3035
rect 7630 2965 8000 2975
rect 8030 3295 8400 3305
rect 8030 3235 8034 3295
rect 8086 3275 8344 3295
rect 8030 3229 8086 3235
rect 8030 3041 8060 3229
rect 8115 3220 8315 3245
rect 8396 3235 8400 3295
rect 8344 3229 8400 3235
rect 8115 3200 8185 3220
rect 8090 3160 8185 3200
rect 8245 3200 8315 3220
rect 8245 3160 8340 3200
rect 8090 3110 8340 3160
rect 8090 3070 8185 3110
rect 8115 3050 8185 3070
rect 8245 3070 8340 3110
rect 8245 3050 8315 3070
rect 8030 3035 8086 3041
rect 8030 2975 8034 3035
rect 8115 3025 8315 3050
rect 8370 3041 8400 3229
rect 8344 3035 8400 3041
rect 8086 2975 8344 2995
rect 8396 2975 8400 3035
rect 8030 2965 8400 2975
rect 8430 3295 8800 3305
rect 8430 3235 8434 3295
rect 8486 3275 8744 3295
rect 8430 3229 8486 3235
rect 8430 3041 8460 3229
rect 8515 3220 8715 3245
rect 8796 3235 8800 3295
rect 8744 3229 8800 3235
rect 8515 3200 8585 3220
rect 8490 3160 8585 3200
rect 8645 3200 8715 3220
rect 8645 3160 8740 3200
rect 8490 3110 8740 3160
rect 8490 3070 8585 3110
rect 8515 3050 8585 3070
rect 8645 3070 8740 3110
rect 8645 3050 8715 3070
rect 8430 3035 8486 3041
rect 8430 2975 8434 3035
rect 8515 3025 8715 3050
rect 8770 3041 8800 3229
rect 8744 3035 8800 3041
rect 8486 2975 8744 2995
rect 8796 2975 8800 3035
rect 8430 2965 8800 2975
rect 8830 3295 9200 3305
rect 8830 3235 8834 3295
rect 8886 3275 9144 3295
rect 8830 3229 8886 3235
rect 8830 3041 8860 3229
rect 8915 3220 9115 3245
rect 9196 3235 9200 3295
rect 9144 3229 9200 3235
rect 8915 3200 8985 3220
rect 8890 3160 8985 3200
rect 9045 3200 9115 3220
rect 9045 3160 9140 3200
rect 8890 3110 9140 3160
rect 8890 3070 8985 3110
rect 8915 3050 8985 3070
rect 9045 3070 9140 3110
rect 9045 3050 9115 3070
rect 8830 3035 8886 3041
rect 8830 2975 8834 3035
rect 8915 3025 9115 3050
rect 9170 3041 9200 3229
rect 9144 3035 9200 3041
rect 8886 2975 9144 2995
rect 9196 2975 9200 3035
rect 8830 2965 9200 2975
rect 9230 3295 9600 3305
rect 9230 3235 9234 3295
rect 9286 3275 9544 3295
rect 9230 3229 9286 3235
rect 9230 3041 9260 3229
rect 9315 3220 9515 3245
rect 9596 3235 9600 3295
rect 9544 3229 9600 3235
rect 9315 3200 9385 3220
rect 9290 3160 9385 3200
rect 9445 3200 9515 3220
rect 9445 3160 9540 3200
rect 9290 3110 9540 3160
rect 9290 3070 9385 3110
rect 9315 3050 9385 3070
rect 9445 3070 9540 3110
rect 9445 3050 9515 3070
rect 9230 3035 9286 3041
rect 9230 2975 9234 3035
rect 9315 3025 9515 3050
rect 9570 3041 9600 3229
rect 9544 3035 9600 3041
rect 9286 2975 9544 2995
rect 9596 2975 9600 3035
rect 9230 2965 9600 2975
rect 9630 3295 10000 3305
rect 9630 3235 9634 3295
rect 9686 3275 9944 3295
rect 9630 3229 9686 3235
rect 9630 3041 9660 3229
rect 9715 3220 9915 3245
rect 9996 3235 10000 3295
rect 9944 3229 10000 3235
rect 9715 3200 9785 3220
rect 9690 3160 9785 3200
rect 9845 3200 9915 3220
rect 9845 3160 9940 3200
rect 9690 3110 9940 3160
rect 9690 3070 9785 3110
rect 9715 3050 9785 3070
rect 9845 3070 9940 3110
rect 9845 3050 9915 3070
rect 9630 3035 9686 3041
rect 9630 2975 9634 3035
rect 9715 3025 9915 3050
rect 9970 3041 10000 3229
rect 9944 3035 10000 3041
rect 9686 2975 9944 2995
rect 9996 2975 10000 3035
rect 9630 2965 10000 2975
rect 10030 3295 10400 3305
rect 10030 3235 10034 3295
rect 10086 3275 10344 3295
rect 10030 3229 10086 3235
rect 10030 3041 10060 3229
rect 10115 3220 10315 3245
rect 10396 3235 10400 3295
rect 10344 3229 10400 3235
rect 10115 3200 10185 3220
rect 10090 3160 10185 3200
rect 10245 3200 10315 3220
rect 10245 3160 10340 3200
rect 10090 3110 10340 3160
rect 10090 3070 10185 3110
rect 10115 3050 10185 3070
rect 10245 3070 10340 3110
rect 10245 3050 10315 3070
rect 10030 3035 10086 3041
rect 10030 2975 10034 3035
rect 10115 3025 10315 3050
rect 10370 3041 10400 3229
rect 10344 3035 10400 3041
rect 10086 2975 10344 2995
rect 10396 2975 10400 3035
rect 10030 2965 10400 2975
rect 10430 3295 10800 3305
rect 10430 3235 10434 3295
rect 10486 3275 10744 3295
rect 10430 3229 10486 3235
rect 10430 3041 10460 3229
rect 10515 3220 10715 3245
rect 10796 3235 10800 3295
rect 10744 3229 10800 3235
rect 10515 3200 10585 3220
rect 10490 3160 10585 3200
rect 10645 3200 10715 3220
rect 10645 3160 10740 3200
rect 10490 3110 10740 3160
rect 10490 3070 10585 3110
rect 10515 3050 10585 3070
rect 10645 3070 10740 3110
rect 10645 3050 10715 3070
rect 10430 3035 10486 3041
rect 10430 2975 10434 3035
rect 10515 3025 10715 3050
rect 10770 3041 10800 3229
rect 10744 3035 10800 3041
rect 10486 2975 10744 2995
rect 10796 2975 10800 3035
rect 10430 2965 10800 2975
rect 10830 3295 11200 3305
rect 10830 3235 10834 3295
rect 10886 3275 11144 3295
rect 10830 3229 10886 3235
rect 10830 3041 10860 3229
rect 10915 3220 11115 3245
rect 11196 3235 11200 3295
rect 11144 3229 11200 3235
rect 10915 3200 10985 3220
rect 10890 3160 10985 3200
rect 11045 3200 11115 3220
rect 11045 3160 11140 3200
rect 10890 3110 11140 3160
rect 10890 3070 10985 3110
rect 10915 3050 10985 3070
rect 11045 3070 11140 3110
rect 11045 3050 11115 3070
rect 10830 3035 10886 3041
rect 10830 2975 10834 3035
rect 10915 3025 11115 3050
rect 11170 3041 11200 3229
rect 11144 3035 11200 3041
rect 10886 2975 11144 2995
rect 11196 2975 11200 3035
rect 10830 2965 11200 2975
rect 11230 3295 11600 3305
rect 11230 3235 11234 3295
rect 11286 3275 11544 3295
rect 11230 3229 11286 3235
rect 11230 3041 11260 3229
rect 11315 3220 11515 3245
rect 11596 3235 11600 3295
rect 11544 3229 11600 3235
rect 11315 3200 11385 3220
rect 11290 3160 11385 3200
rect 11445 3200 11515 3220
rect 11445 3160 11540 3200
rect 11290 3110 11540 3160
rect 11290 3070 11385 3110
rect 11315 3050 11385 3070
rect 11445 3070 11540 3110
rect 11445 3050 11515 3070
rect 11230 3035 11286 3041
rect 11230 2975 11234 3035
rect 11315 3025 11515 3050
rect 11570 3041 11600 3229
rect 11544 3035 11600 3041
rect 11286 2975 11544 2995
rect 11596 2975 11600 3035
rect 11230 2965 11600 2975
rect 11630 3295 12000 3305
rect 11630 3235 11634 3295
rect 11686 3275 11944 3295
rect 11630 3229 11686 3235
rect 11630 3041 11660 3229
rect 11715 3220 11915 3245
rect 11996 3235 12000 3295
rect 11944 3229 12000 3235
rect 11715 3200 11785 3220
rect 11690 3160 11785 3200
rect 11845 3200 11915 3220
rect 11845 3160 11940 3200
rect 11690 3110 11940 3160
rect 11690 3070 11785 3110
rect 11715 3050 11785 3070
rect 11845 3070 11940 3110
rect 11845 3050 11915 3070
rect 11630 3035 11686 3041
rect 11630 2975 11634 3035
rect 11715 3025 11915 3050
rect 11970 3041 12000 3229
rect 11944 3035 12000 3041
rect 11686 2975 11944 2995
rect 11996 2975 12000 3035
rect 11630 2965 12000 2975
rect 12030 3295 12400 3305
rect 12030 3235 12034 3295
rect 12086 3275 12344 3295
rect 12030 3229 12086 3235
rect 12030 3041 12060 3229
rect 12115 3220 12315 3245
rect 12396 3235 12400 3295
rect 12344 3229 12400 3235
rect 12115 3200 12185 3220
rect 12090 3160 12185 3200
rect 12245 3200 12315 3220
rect 12245 3160 12340 3200
rect 12090 3110 12340 3160
rect 12090 3070 12185 3110
rect 12115 3050 12185 3070
rect 12245 3070 12340 3110
rect 12245 3050 12315 3070
rect 12030 3035 12086 3041
rect 12030 2975 12034 3035
rect 12115 3025 12315 3050
rect 12370 3041 12400 3229
rect 12344 3035 12400 3041
rect 12086 2975 12344 2995
rect 12396 2975 12400 3035
rect 12030 2965 12400 2975
rect 12430 3295 12800 3305
rect 12430 3235 12434 3295
rect 12486 3275 12744 3295
rect 12430 3229 12486 3235
rect 12430 3041 12460 3229
rect 12515 3220 12715 3245
rect 12796 3235 12800 3295
rect 12744 3229 12800 3235
rect 12515 3200 12585 3220
rect 12490 3160 12585 3200
rect 12645 3200 12715 3220
rect 12645 3160 12740 3200
rect 12490 3110 12740 3160
rect 12490 3070 12585 3110
rect 12515 3050 12585 3070
rect 12645 3070 12740 3110
rect 12645 3050 12715 3070
rect 12430 3035 12486 3041
rect 12430 2975 12434 3035
rect 12515 3025 12715 3050
rect 12770 3041 12800 3229
rect 12744 3035 12800 3041
rect 12486 2975 12744 2995
rect 12796 2975 12800 3035
rect 12430 2965 12800 2975
rect 12830 3295 13200 3305
rect 12830 3235 12834 3295
rect 12886 3275 13144 3295
rect 12830 3229 12886 3235
rect 12830 3041 12860 3229
rect 12915 3220 13115 3245
rect 13196 3235 13200 3295
rect 13144 3229 13200 3235
rect 12915 3200 12985 3220
rect 12890 3160 12985 3200
rect 13045 3200 13115 3220
rect 13045 3160 13140 3200
rect 12890 3110 13140 3160
rect 12890 3070 12985 3110
rect 12915 3050 12985 3070
rect 13045 3070 13140 3110
rect 13045 3050 13115 3070
rect 12830 3035 12886 3041
rect 12830 2975 12834 3035
rect 12915 3025 13115 3050
rect 13170 3041 13200 3229
rect 13144 3035 13200 3041
rect 12886 2975 13144 2995
rect 13196 2975 13200 3035
rect 12830 2965 13200 2975
rect -370 2925 0 2935
rect -370 2865 -366 2925
rect -314 2905 -56 2925
rect -370 2859 -314 2865
rect -370 2671 -340 2859
rect -285 2850 -85 2875
rect -4 2865 0 2925
rect -56 2859 0 2865
rect -285 2830 -215 2850
rect -310 2790 -215 2830
rect -155 2830 -85 2850
rect -155 2790 -60 2830
rect -310 2740 -60 2790
rect -310 2700 -215 2740
rect -285 2680 -215 2700
rect -155 2700 -60 2740
rect -155 2680 -85 2700
rect -370 2665 -314 2671
rect -370 2605 -366 2665
rect -285 2655 -85 2680
rect -30 2671 0 2859
rect -56 2665 0 2671
rect -314 2605 -56 2625
rect -4 2605 0 2665
rect -370 2595 0 2605
rect 30 2925 400 2935
rect 30 2865 34 2925
rect 86 2905 344 2925
rect 30 2859 86 2865
rect 30 2671 60 2859
rect 115 2850 315 2875
rect 396 2865 400 2925
rect 344 2859 400 2865
rect 115 2830 185 2850
rect 90 2790 185 2830
rect 245 2830 315 2850
rect 245 2790 340 2830
rect 90 2740 340 2790
rect 90 2700 185 2740
rect 115 2680 185 2700
rect 245 2700 340 2740
rect 245 2680 315 2700
rect 30 2665 86 2671
rect 30 2605 34 2665
rect 115 2655 315 2680
rect 370 2671 400 2859
rect 344 2665 400 2671
rect 86 2605 344 2625
rect 396 2605 400 2665
rect 30 2595 400 2605
rect 430 2925 800 2935
rect 430 2865 434 2925
rect 486 2905 744 2925
rect 430 2859 486 2865
rect 430 2671 460 2859
rect 515 2850 715 2875
rect 796 2865 800 2925
rect 744 2859 800 2865
rect 515 2830 585 2850
rect 490 2790 585 2830
rect 645 2830 715 2850
rect 645 2790 740 2830
rect 490 2740 740 2790
rect 490 2700 585 2740
rect 515 2680 585 2700
rect 645 2700 740 2740
rect 645 2680 715 2700
rect 430 2665 486 2671
rect 430 2605 434 2665
rect 515 2655 715 2680
rect 770 2671 800 2859
rect 744 2665 800 2671
rect 486 2605 744 2625
rect 796 2605 800 2665
rect 430 2595 800 2605
rect 830 2925 1200 2935
rect 830 2865 834 2925
rect 886 2905 1144 2925
rect 830 2859 886 2865
rect 830 2671 860 2859
rect 915 2850 1115 2875
rect 1196 2865 1200 2925
rect 1144 2859 1200 2865
rect 915 2830 985 2850
rect 890 2790 985 2830
rect 1045 2830 1115 2850
rect 1045 2790 1140 2830
rect 890 2740 1140 2790
rect 890 2700 985 2740
rect 915 2680 985 2700
rect 1045 2700 1140 2740
rect 1045 2680 1115 2700
rect 830 2665 886 2671
rect 830 2605 834 2665
rect 915 2655 1115 2680
rect 1170 2671 1200 2859
rect 1144 2665 1200 2671
rect 886 2605 1144 2625
rect 1196 2605 1200 2665
rect 830 2595 1200 2605
rect 1230 2925 1600 2935
rect 1230 2865 1234 2925
rect 1286 2905 1544 2925
rect 1230 2859 1286 2865
rect 1230 2671 1260 2859
rect 1315 2850 1515 2875
rect 1596 2865 1600 2925
rect 1544 2859 1600 2865
rect 1315 2830 1385 2850
rect 1290 2790 1385 2830
rect 1445 2830 1515 2850
rect 1445 2790 1540 2830
rect 1290 2740 1540 2790
rect 1290 2700 1385 2740
rect 1315 2680 1385 2700
rect 1445 2700 1540 2740
rect 1445 2680 1515 2700
rect 1230 2665 1286 2671
rect 1230 2605 1234 2665
rect 1315 2655 1515 2680
rect 1570 2671 1600 2859
rect 1544 2665 1600 2671
rect 1286 2605 1544 2625
rect 1596 2605 1600 2665
rect 1230 2595 1600 2605
rect 1630 2925 2000 2935
rect 1630 2865 1634 2925
rect 1686 2905 1944 2925
rect 1630 2859 1686 2865
rect 1630 2671 1660 2859
rect 1715 2850 1915 2875
rect 1996 2865 2000 2925
rect 1944 2859 2000 2865
rect 1715 2830 1785 2850
rect 1690 2790 1785 2830
rect 1845 2830 1915 2850
rect 1845 2790 1940 2830
rect 1690 2740 1940 2790
rect 1690 2700 1785 2740
rect 1715 2680 1785 2700
rect 1845 2700 1940 2740
rect 1845 2680 1915 2700
rect 1630 2665 1686 2671
rect 1630 2605 1634 2665
rect 1715 2655 1915 2680
rect 1970 2671 2000 2859
rect 1944 2665 2000 2671
rect 1686 2605 1944 2625
rect 1996 2605 2000 2665
rect 1630 2595 2000 2605
rect 2030 2925 2400 2935
rect 2030 2865 2034 2925
rect 2086 2905 2344 2925
rect 2030 2859 2086 2865
rect 2030 2671 2060 2859
rect 2115 2850 2315 2875
rect 2396 2865 2400 2925
rect 2344 2859 2400 2865
rect 2115 2830 2185 2850
rect 2090 2790 2185 2830
rect 2245 2830 2315 2850
rect 2245 2790 2340 2830
rect 2090 2740 2340 2790
rect 2090 2700 2185 2740
rect 2115 2680 2185 2700
rect 2245 2700 2340 2740
rect 2245 2680 2315 2700
rect 2030 2665 2086 2671
rect 2030 2605 2034 2665
rect 2115 2655 2315 2680
rect 2370 2671 2400 2859
rect 2344 2665 2400 2671
rect 2086 2605 2344 2625
rect 2396 2605 2400 2665
rect 2030 2595 2400 2605
rect 2430 2925 2800 2935
rect 2430 2865 2434 2925
rect 2486 2905 2744 2925
rect 2430 2859 2486 2865
rect 2430 2671 2460 2859
rect 2515 2850 2715 2875
rect 2796 2865 2800 2925
rect 2744 2859 2800 2865
rect 2515 2830 2585 2850
rect 2490 2790 2585 2830
rect 2645 2830 2715 2850
rect 2645 2790 2740 2830
rect 2490 2740 2740 2790
rect 2490 2700 2585 2740
rect 2515 2680 2585 2700
rect 2645 2700 2740 2740
rect 2645 2680 2715 2700
rect 2430 2665 2486 2671
rect 2430 2605 2434 2665
rect 2515 2655 2715 2680
rect 2770 2671 2800 2859
rect 2744 2665 2800 2671
rect 2486 2605 2744 2625
rect 2796 2605 2800 2665
rect 2430 2595 2800 2605
rect 2830 2925 3200 2935
rect 2830 2865 2834 2925
rect 2886 2905 3144 2925
rect 2830 2859 2886 2865
rect 2830 2671 2860 2859
rect 2915 2850 3115 2875
rect 3196 2865 3200 2925
rect 3144 2859 3200 2865
rect 2915 2830 2985 2850
rect 2890 2790 2985 2830
rect 3045 2830 3115 2850
rect 3045 2790 3140 2830
rect 2890 2740 3140 2790
rect 2890 2700 2985 2740
rect 2915 2680 2985 2700
rect 3045 2700 3140 2740
rect 3045 2680 3115 2700
rect 2830 2665 2886 2671
rect 2830 2605 2834 2665
rect 2915 2655 3115 2680
rect 3170 2671 3200 2859
rect 3144 2665 3200 2671
rect 2886 2605 3144 2625
rect 3196 2605 3200 2665
rect 2830 2595 3200 2605
rect 3230 2925 3600 2935
rect 3230 2865 3234 2925
rect 3286 2905 3544 2925
rect 3230 2859 3286 2865
rect 3230 2671 3260 2859
rect 3315 2850 3515 2875
rect 3596 2865 3600 2925
rect 3544 2859 3600 2865
rect 3315 2830 3385 2850
rect 3290 2790 3385 2830
rect 3445 2830 3515 2850
rect 3445 2790 3540 2830
rect 3290 2740 3540 2790
rect 3290 2700 3385 2740
rect 3315 2680 3385 2700
rect 3445 2700 3540 2740
rect 3445 2680 3515 2700
rect 3230 2665 3286 2671
rect 3230 2605 3234 2665
rect 3315 2655 3515 2680
rect 3570 2671 3600 2859
rect 3544 2665 3600 2671
rect 3286 2605 3544 2625
rect 3596 2605 3600 2665
rect 3230 2595 3600 2605
rect 3630 2925 4000 2935
rect 3630 2865 3634 2925
rect 3686 2905 3944 2925
rect 3630 2859 3686 2865
rect 3630 2671 3660 2859
rect 3715 2850 3915 2875
rect 3996 2865 4000 2925
rect 3944 2859 4000 2865
rect 3715 2830 3785 2850
rect 3690 2790 3785 2830
rect 3845 2830 3915 2850
rect 3845 2790 3940 2830
rect 3690 2740 3940 2790
rect 3690 2700 3785 2740
rect 3715 2680 3785 2700
rect 3845 2700 3940 2740
rect 3845 2680 3915 2700
rect 3630 2665 3686 2671
rect 3630 2605 3634 2665
rect 3715 2655 3915 2680
rect 3970 2671 4000 2859
rect 3944 2665 4000 2671
rect 3686 2605 3944 2625
rect 3996 2605 4000 2665
rect 3630 2595 4000 2605
rect 4030 2925 4400 2935
rect 4030 2865 4034 2925
rect 4086 2905 4344 2925
rect 4030 2859 4086 2865
rect 4030 2671 4060 2859
rect 4115 2850 4315 2875
rect 4396 2865 4400 2925
rect 4344 2859 4400 2865
rect 4115 2830 4185 2850
rect 4090 2790 4185 2830
rect 4245 2830 4315 2850
rect 4245 2790 4340 2830
rect 4090 2740 4340 2790
rect 4090 2700 4185 2740
rect 4115 2680 4185 2700
rect 4245 2700 4340 2740
rect 4245 2680 4315 2700
rect 4030 2665 4086 2671
rect 4030 2605 4034 2665
rect 4115 2655 4315 2680
rect 4370 2671 4400 2859
rect 4344 2665 4400 2671
rect 4086 2605 4344 2625
rect 4396 2605 4400 2665
rect 4030 2595 4400 2605
rect 4430 2925 4800 2935
rect 4430 2865 4434 2925
rect 4486 2905 4744 2925
rect 4430 2859 4486 2865
rect 4430 2671 4460 2859
rect 4515 2850 4715 2875
rect 4796 2865 4800 2925
rect 4744 2859 4800 2865
rect 4515 2830 4585 2850
rect 4490 2790 4585 2830
rect 4645 2830 4715 2850
rect 4645 2790 4740 2830
rect 4490 2740 4740 2790
rect 4490 2700 4585 2740
rect 4515 2680 4585 2700
rect 4645 2700 4740 2740
rect 4645 2680 4715 2700
rect 4430 2665 4486 2671
rect 4430 2605 4434 2665
rect 4515 2655 4715 2680
rect 4770 2671 4800 2859
rect 4744 2665 4800 2671
rect 4486 2605 4744 2625
rect 4796 2605 4800 2665
rect 4430 2595 4800 2605
rect 4830 2925 5200 2935
rect 4830 2865 4834 2925
rect 4886 2905 5144 2925
rect 4830 2859 4886 2865
rect 4830 2671 4860 2859
rect 4915 2850 5115 2875
rect 5196 2865 5200 2925
rect 5144 2859 5200 2865
rect 4915 2830 4985 2850
rect 4890 2790 4985 2830
rect 5045 2830 5115 2850
rect 5045 2790 5140 2830
rect 4890 2740 5140 2790
rect 4890 2700 4985 2740
rect 4915 2680 4985 2700
rect 5045 2700 5140 2740
rect 5045 2680 5115 2700
rect 4830 2665 4886 2671
rect 4830 2605 4834 2665
rect 4915 2655 5115 2680
rect 5170 2671 5200 2859
rect 5144 2665 5200 2671
rect 4886 2605 5144 2625
rect 5196 2605 5200 2665
rect 4830 2595 5200 2605
rect 5230 2925 5600 2935
rect 5230 2865 5234 2925
rect 5286 2905 5544 2925
rect 5230 2859 5286 2865
rect 5230 2671 5260 2859
rect 5315 2850 5515 2875
rect 5596 2865 5600 2925
rect 5544 2859 5600 2865
rect 5315 2830 5385 2850
rect 5290 2790 5385 2830
rect 5445 2830 5515 2850
rect 5445 2790 5540 2830
rect 5290 2740 5540 2790
rect 5290 2700 5385 2740
rect 5315 2680 5385 2700
rect 5445 2700 5540 2740
rect 5445 2680 5515 2700
rect 5230 2665 5286 2671
rect 5230 2605 5234 2665
rect 5315 2655 5515 2680
rect 5570 2671 5600 2859
rect 5544 2665 5600 2671
rect 5286 2605 5544 2625
rect 5596 2605 5600 2665
rect 5230 2595 5600 2605
rect 5630 2925 6000 2935
rect 5630 2865 5634 2925
rect 5686 2905 5944 2925
rect 5630 2859 5686 2865
rect 5630 2671 5660 2859
rect 5715 2850 5915 2875
rect 5996 2865 6000 2925
rect 5944 2859 6000 2865
rect 5715 2830 5785 2850
rect 5690 2790 5785 2830
rect 5845 2830 5915 2850
rect 5845 2790 5940 2830
rect 5690 2740 5940 2790
rect 5690 2700 5785 2740
rect 5715 2680 5785 2700
rect 5845 2700 5940 2740
rect 5845 2680 5915 2700
rect 5630 2665 5686 2671
rect 5630 2605 5634 2665
rect 5715 2655 5915 2680
rect 5970 2671 6000 2859
rect 5944 2665 6000 2671
rect 5686 2605 5944 2625
rect 5996 2605 6000 2665
rect 5630 2595 6000 2605
rect 6030 2925 6400 2935
rect 6030 2865 6034 2925
rect 6086 2905 6344 2925
rect 6030 2859 6086 2865
rect 6030 2671 6060 2859
rect 6115 2850 6315 2875
rect 6396 2865 6400 2925
rect 6344 2859 6400 2865
rect 6115 2830 6185 2850
rect 6090 2790 6185 2830
rect 6245 2830 6315 2850
rect 6245 2790 6340 2830
rect 6090 2740 6340 2790
rect 6090 2700 6185 2740
rect 6115 2680 6185 2700
rect 6245 2700 6340 2740
rect 6245 2680 6315 2700
rect 6030 2665 6086 2671
rect 6030 2605 6034 2665
rect 6115 2655 6315 2680
rect 6370 2671 6400 2859
rect 6344 2665 6400 2671
rect 6086 2605 6344 2625
rect 6396 2605 6400 2665
rect 6030 2595 6400 2605
rect 6430 2925 6800 2935
rect 6430 2865 6434 2925
rect 6486 2905 6744 2925
rect 6430 2859 6486 2865
rect 6430 2671 6460 2859
rect 6515 2850 6715 2875
rect 6796 2865 6800 2925
rect 6744 2859 6800 2865
rect 6515 2830 6585 2850
rect 6490 2790 6585 2830
rect 6645 2830 6715 2850
rect 6645 2790 6740 2830
rect 6490 2740 6740 2790
rect 6490 2700 6585 2740
rect 6515 2680 6585 2700
rect 6645 2700 6740 2740
rect 6645 2680 6715 2700
rect 6430 2665 6486 2671
rect 6430 2605 6434 2665
rect 6515 2655 6715 2680
rect 6770 2671 6800 2859
rect 6744 2665 6800 2671
rect 6486 2605 6744 2625
rect 6796 2605 6800 2665
rect 6430 2595 6800 2605
rect 6830 2925 7200 2935
rect 6830 2865 6834 2925
rect 6886 2905 7144 2925
rect 6830 2859 6886 2865
rect 6830 2671 6860 2859
rect 6915 2850 7115 2875
rect 7196 2865 7200 2925
rect 7144 2859 7200 2865
rect 6915 2830 6985 2850
rect 6890 2790 6985 2830
rect 7045 2830 7115 2850
rect 7045 2790 7140 2830
rect 6890 2740 7140 2790
rect 6890 2700 6985 2740
rect 6915 2680 6985 2700
rect 7045 2700 7140 2740
rect 7045 2680 7115 2700
rect 6830 2665 6886 2671
rect 6830 2605 6834 2665
rect 6915 2655 7115 2680
rect 7170 2671 7200 2859
rect 7144 2665 7200 2671
rect 6886 2605 7144 2625
rect 7196 2605 7200 2665
rect 6830 2595 7200 2605
rect 7230 2925 7600 2935
rect 7230 2865 7234 2925
rect 7286 2905 7544 2925
rect 7230 2859 7286 2865
rect 7230 2671 7260 2859
rect 7315 2850 7515 2875
rect 7596 2865 7600 2925
rect 7544 2859 7600 2865
rect 7315 2830 7385 2850
rect 7290 2790 7385 2830
rect 7445 2830 7515 2850
rect 7445 2790 7540 2830
rect 7290 2740 7540 2790
rect 7290 2700 7385 2740
rect 7315 2680 7385 2700
rect 7445 2700 7540 2740
rect 7445 2680 7515 2700
rect 7230 2665 7286 2671
rect 7230 2605 7234 2665
rect 7315 2655 7515 2680
rect 7570 2671 7600 2859
rect 7544 2665 7600 2671
rect 7286 2605 7544 2625
rect 7596 2605 7600 2665
rect 7230 2595 7600 2605
rect 7630 2925 8000 2935
rect 7630 2865 7634 2925
rect 7686 2905 7944 2925
rect 7630 2859 7686 2865
rect 7630 2671 7660 2859
rect 7715 2850 7915 2875
rect 7996 2865 8000 2925
rect 7944 2859 8000 2865
rect 7715 2830 7785 2850
rect 7690 2790 7785 2830
rect 7845 2830 7915 2850
rect 7845 2790 7940 2830
rect 7690 2740 7940 2790
rect 7690 2700 7785 2740
rect 7715 2680 7785 2700
rect 7845 2700 7940 2740
rect 7845 2680 7915 2700
rect 7630 2665 7686 2671
rect 7630 2605 7634 2665
rect 7715 2655 7915 2680
rect 7970 2671 8000 2859
rect 7944 2665 8000 2671
rect 7686 2605 7944 2625
rect 7996 2605 8000 2665
rect 7630 2595 8000 2605
rect 8030 2925 8400 2935
rect 8030 2865 8034 2925
rect 8086 2905 8344 2925
rect 8030 2859 8086 2865
rect 8030 2671 8060 2859
rect 8115 2850 8315 2875
rect 8396 2865 8400 2925
rect 8344 2859 8400 2865
rect 8115 2830 8185 2850
rect 8090 2790 8185 2830
rect 8245 2830 8315 2850
rect 8245 2790 8340 2830
rect 8090 2740 8340 2790
rect 8090 2700 8185 2740
rect 8115 2680 8185 2700
rect 8245 2700 8340 2740
rect 8245 2680 8315 2700
rect 8030 2665 8086 2671
rect 8030 2605 8034 2665
rect 8115 2655 8315 2680
rect 8370 2671 8400 2859
rect 8344 2665 8400 2671
rect 8086 2605 8344 2625
rect 8396 2605 8400 2665
rect 8030 2595 8400 2605
rect 8430 2925 8800 2935
rect 8430 2865 8434 2925
rect 8486 2905 8744 2925
rect 8430 2859 8486 2865
rect 8430 2671 8460 2859
rect 8515 2850 8715 2875
rect 8796 2865 8800 2925
rect 8744 2859 8800 2865
rect 8515 2830 8585 2850
rect 8490 2790 8585 2830
rect 8645 2830 8715 2850
rect 8645 2790 8740 2830
rect 8490 2740 8740 2790
rect 8490 2700 8585 2740
rect 8515 2680 8585 2700
rect 8645 2700 8740 2740
rect 8645 2680 8715 2700
rect 8430 2665 8486 2671
rect 8430 2605 8434 2665
rect 8515 2655 8715 2680
rect 8770 2671 8800 2859
rect 8744 2665 8800 2671
rect 8486 2605 8744 2625
rect 8796 2605 8800 2665
rect 8430 2595 8800 2605
rect 8830 2925 9200 2935
rect 8830 2865 8834 2925
rect 8886 2905 9144 2925
rect 8830 2859 8886 2865
rect 8830 2671 8860 2859
rect 8915 2850 9115 2875
rect 9196 2865 9200 2925
rect 9144 2859 9200 2865
rect 8915 2830 8985 2850
rect 8890 2790 8985 2830
rect 9045 2830 9115 2850
rect 9045 2790 9140 2830
rect 8890 2740 9140 2790
rect 8890 2700 8985 2740
rect 8915 2680 8985 2700
rect 9045 2700 9140 2740
rect 9045 2680 9115 2700
rect 8830 2665 8886 2671
rect 8830 2605 8834 2665
rect 8915 2655 9115 2680
rect 9170 2671 9200 2859
rect 9144 2665 9200 2671
rect 8886 2605 9144 2625
rect 9196 2605 9200 2665
rect 8830 2595 9200 2605
rect 9230 2925 9600 2935
rect 9230 2865 9234 2925
rect 9286 2905 9544 2925
rect 9230 2859 9286 2865
rect 9230 2671 9260 2859
rect 9315 2850 9515 2875
rect 9596 2865 9600 2925
rect 9544 2859 9600 2865
rect 9315 2830 9385 2850
rect 9290 2790 9385 2830
rect 9445 2830 9515 2850
rect 9445 2790 9540 2830
rect 9290 2740 9540 2790
rect 9290 2700 9385 2740
rect 9315 2680 9385 2700
rect 9445 2700 9540 2740
rect 9445 2680 9515 2700
rect 9230 2665 9286 2671
rect 9230 2605 9234 2665
rect 9315 2655 9515 2680
rect 9570 2671 9600 2859
rect 9544 2665 9600 2671
rect 9286 2605 9544 2625
rect 9596 2605 9600 2665
rect 9230 2595 9600 2605
rect 9630 2925 10000 2935
rect 9630 2865 9634 2925
rect 9686 2905 9944 2925
rect 9630 2859 9686 2865
rect 9630 2671 9660 2859
rect 9715 2850 9915 2875
rect 9996 2865 10000 2925
rect 9944 2859 10000 2865
rect 9715 2830 9785 2850
rect 9690 2790 9785 2830
rect 9845 2830 9915 2850
rect 9845 2790 9940 2830
rect 9690 2740 9940 2790
rect 9690 2700 9785 2740
rect 9715 2680 9785 2700
rect 9845 2700 9940 2740
rect 9845 2680 9915 2700
rect 9630 2665 9686 2671
rect 9630 2605 9634 2665
rect 9715 2655 9915 2680
rect 9970 2671 10000 2859
rect 9944 2665 10000 2671
rect 9686 2605 9944 2625
rect 9996 2605 10000 2665
rect 9630 2595 10000 2605
rect 10030 2925 10400 2935
rect 10030 2865 10034 2925
rect 10086 2905 10344 2925
rect 10030 2859 10086 2865
rect 10030 2671 10060 2859
rect 10115 2850 10315 2875
rect 10396 2865 10400 2925
rect 10344 2859 10400 2865
rect 10115 2830 10185 2850
rect 10090 2790 10185 2830
rect 10245 2830 10315 2850
rect 10245 2790 10340 2830
rect 10090 2740 10340 2790
rect 10090 2700 10185 2740
rect 10115 2680 10185 2700
rect 10245 2700 10340 2740
rect 10245 2680 10315 2700
rect 10030 2665 10086 2671
rect 10030 2605 10034 2665
rect 10115 2655 10315 2680
rect 10370 2671 10400 2859
rect 10344 2665 10400 2671
rect 10086 2605 10344 2625
rect 10396 2605 10400 2665
rect 10030 2595 10400 2605
rect 10430 2925 10800 2935
rect 10430 2865 10434 2925
rect 10486 2905 10744 2925
rect 10430 2859 10486 2865
rect 10430 2671 10460 2859
rect 10515 2850 10715 2875
rect 10796 2865 10800 2925
rect 10744 2859 10800 2865
rect 10515 2830 10585 2850
rect 10490 2790 10585 2830
rect 10645 2830 10715 2850
rect 10645 2790 10740 2830
rect 10490 2740 10740 2790
rect 10490 2700 10585 2740
rect 10515 2680 10585 2700
rect 10645 2700 10740 2740
rect 10645 2680 10715 2700
rect 10430 2665 10486 2671
rect 10430 2605 10434 2665
rect 10515 2655 10715 2680
rect 10770 2671 10800 2859
rect 10744 2665 10800 2671
rect 10486 2605 10744 2625
rect 10796 2605 10800 2665
rect 10430 2595 10800 2605
rect 10830 2925 11200 2935
rect 10830 2865 10834 2925
rect 10886 2905 11144 2925
rect 10830 2859 10886 2865
rect 10830 2671 10860 2859
rect 10915 2850 11115 2875
rect 11196 2865 11200 2925
rect 11144 2859 11200 2865
rect 10915 2830 10985 2850
rect 10890 2790 10985 2830
rect 11045 2830 11115 2850
rect 11045 2790 11140 2830
rect 10890 2740 11140 2790
rect 10890 2700 10985 2740
rect 10915 2680 10985 2700
rect 11045 2700 11140 2740
rect 11045 2680 11115 2700
rect 10830 2665 10886 2671
rect 10830 2605 10834 2665
rect 10915 2655 11115 2680
rect 11170 2671 11200 2859
rect 11144 2665 11200 2671
rect 10886 2605 11144 2625
rect 11196 2605 11200 2665
rect 10830 2595 11200 2605
rect 11230 2925 11600 2935
rect 11230 2865 11234 2925
rect 11286 2905 11544 2925
rect 11230 2859 11286 2865
rect 11230 2671 11260 2859
rect 11315 2850 11515 2875
rect 11596 2865 11600 2925
rect 11544 2859 11600 2865
rect 11315 2830 11385 2850
rect 11290 2790 11385 2830
rect 11445 2830 11515 2850
rect 11445 2790 11540 2830
rect 11290 2740 11540 2790
rect 11290 2700 11385 2740
rect 11315 2680 11385 2700
rect 11445 2700 11540 2740
rect 11445 2680 11515 2700
rect 11230 2665 11286 2671
rect 11230 2605 11234 2665
rect 11315 2655 11515 2680
rect 11570 2671 11600 2859
rect 11544 2665 11600 2671
rect 11286 2605 11544 2625
rect 11596 2605 11600 2665
rect 11230 2595 11600 2605
rect 11630 2925 12000 2935
rect 11630 2865 11634 2925
rect 11686 2905 11944 2925
rect 11630 2859 11686 2865
rect 11630 2671 11660 2859
rect 11715 2850 11915 2875
rect 11996 2865 12000 2925
rect 11944 2859 12000 2865
rect 11715 2830 11785 2850
rect 11690 2790 11785 2830
rect 11845 2830 11915 2850
rect 11845 2790 11940 2830
rect 11690 2740 11940 2790
rect 11690 2700 11785 2740
rect 11715 2680 11785 2700
rect 11845 2700 11940 2740
rect 11845 2680 11915 2700
rect 11630 2665 11686 2671
rect 11630 2605 11634 2665
rect 11715 2655 11915 2680
rect 11970 2671 12000 2859
rect 11944 2665 12000 2671
rect 11686 2605 11944 2625
rect 11996 2605 12000 2665
rect 11630 2595 12000 2605
rect 12030 2925 12400 2935
rect 12030 2865 12034 2925
rect 12086 2905 12344 2925
rect 12030 2859 12086 2865
rect 12030 2671 12060 2859
rect 12115 2850 12315 2875
rect 12396 2865 12400 2925
rect 12344 2859 12400 2865
rect 12115 2830 12185 2850
rect 12090 2790 12185 2830
rect 12245 2830 12315 2850
rect 12245 2790 12340 2830
rect 12090 2740 12340 2790
rect 12090 2700 12185 2740
rect 12115 2680 12185 2700
rect 12245 2700 12340 2740
rect 12245 2680 12315 2700
rect 12030 2665 12086 2671
rect 12030 2605 12034 2665
rect 12115 2655 12315 2680
rect 12370 2671 12400 2859
rect 12344 2665 12400 2671
rect 12086 2605 12344 2625
rect 12396 2605 12400 2665
rect 12030 2595 12400 2605
rect 12430 2925 12800 2935
rect 12430 2865 12434 2925
rect 12486 2905 12744 2925
rect 12430 2859 12486 2865
rect 12430 2671 12460 2859
rect 12515 2850 12715 2875
rect 12796 2865 12800 2925
rect 12744 2859 12800 2865
rect 12515 2830 12585 2850
rect 12490 2790 12585 2830
rect 12645 2830 12715 2850
rect 12645 2790 12740 2830
rect 12490 2740 12740 2790
rect 12490 2700 12585 2740
rect 12515 2680 12585 2700
rect 12645 2700 12740 2740
rect 12645 2680 12715 2700
rect 12430 2665 12486 2671
rect 12430 2605 12434 2665
rect 12515 2655 12715 2680
rect 12770 2671 12800 2859
rect 12744 2665 12800 2671
rect 12486 2605 12744 2625
rect 12796 2605 12800 2665
rect 12430 2595 12800 2605
rect 12830 2925 13200 2935
rect 12830 2865 12834 2925
rect 12886 2905 13144 2925
rect 12830 2859 12886 2865
rect 12830 2671 12860 2859
rect 12915 2850 13115 2875
rect 13196 2865 13200 2925
rect 13144 2859 13200 2865
rect 12915 2830 12985 2850
rect 12890 2790 12985 2830
rect 13045 2830 13115 2850
rect 13045 2790 13140 2830
rect 12890 2740 13140 2790
rect 12890 2700 12985 2740
rect 12915 2680 12985 2700
rect 13045 2700 13140 2740
rect 13045 2680 13115 2700
rect 12830 2665 12886 2671
rect 12830 2605 12834 2665
rect 12915 2655 13115 2680
rect 13170 2671 13200 2859
rect 13144 2665 13200 2671
rect 12886 2605 13144 2625
rect 13196 2605 13200 2665
rect 12830 2595 13200 2605
rect -370 2555 0 2565
rect -370 2495 -366 2555
rect -314 2535 -56 2555
rect -370 2489 -314 2495
rect -370 2301 -340 2489
rect -285 2480 -85 2505
rect -4 2495 0 2555
rect -56 2489 0 2495
rect -285 2460 -215 2480
rect -310 2420 -215 2460
rect -155 2460 -85 2480
rect -155 2420 -60 2460
rect -310 2370 -60 2420
rect -310 2330 -215 2370
rect -285 2310 -215 2330
rect -155 2330 -60 2370
rect -155 2310 -85 2330
rect -370 2295 -314 2301
rect -370 2235 -366 2295
rect -285 2285 -85 2310
rect -30 2301 0 2489
rect -56 2295 0 2301
rect -314 2235 -56 2255
rect -4 2235 0 2295
rect -370 2225 0 2235
rect 30 2555 400 2565
rect 30 2495 34 2555
rect 86 2535 344 2555
rect 30 2489 86 2495
rect 30 2301 60 2489
rect 115 2480 315 2505
rect 396 2495 400 2555
rect 344 2489 400 2495
rect 115 2460 185 2480
rect 90 2420 185 2460
rect 245 2460 315 2480
rect 245 2420 340 2460
rect 90 2370 340 2420
rect 90 2330 185 2370
rect 115 2310 185 2330
rect 245 2330 340 2370
rect 245 2310 315 2330
rect 30 2295 86 2301
rect 30 2235 34 2295
rect 115 2285 315 2310
rect 370 2301 400 2489
rect 344 2295 400 2301
rect 86 2235 344 2255
rect 396 2235 400 2295
rect 30 2225 400 2235
rect 430 2555 800 2565
rect 430 2495 434 2555
rect 486 2535 744 2555
rect 430 2489 486 2495
rect 430 2301 460 2489
rect 515 2480 715 2505
rect 796 2495 800 2555
rect 744 2489 800 2495
rect 515 2460 585 2480
rect 490 2420 585 2460
rect 645 2460 715 2480
rect 645 2420 740 2460
rect 490 2370 740 2420
rect 490 2330 585 2370
rect 515 2310 585 2330
rect 645 2330 740 2370
rect 645 2310 715 2330
rect 430 2295 486 2301
rect 430 2235 434 2295
rect 515 2285 715 2310
rect 770 2301 800 2489
rect 744 2295 800 2301
rect 486 2235 744 2255
rect 796 2235 800 2295
rect 430 2225 800 2235
rect 830 2555 1200 2565
rect 830 2495 834 2555
rect 886 2535 1144 2555
rect 830 2489 886 2495
rect 830 2301 860 2489
rect 915 2480 1115 2505
rect 1196 2495 1200 2555
rect 1144 2489 1200 2495
rect 915 2460 985 2480
rect 890 2420 985 2460
rect 1045 2460 1115 2480
rect 1045 2420 1140 2460
rect 890 2370 1140 2420
rect 890 2330 985 2370
rect 915 2310 985 2330
rect 1045 2330 1140 2370
rect 1045 2310 1115 2330
rect 830 2295 886 2301
rect 830 2235 834 2295
rect 915 2285 1115 2310
rect 1170 2301 1200 2489
rect 1144 2295 1200 2301
rect 886 2235 1144 2255
rect 1196 2235 1200 2295
rect 830 2225 1200 2235
rect 1230 2555 1600 2565
rect 1230 2495 1234 2555
rect 1286 2535 1544 2555
rect 1230 2489 1286 2495
rect 1230 2301 1260 2489
rect 1315 2480 1515 2505
rect 1596 2495 1600 2555
rect 1544 2489 1600 2495
rect 1315 2460 1385 2480
rect 1290 2420 1385 2460
rect 1445 2460 1515 2480
rect 1445 2420 1540 2460
rect 1290 2370 1540 2420
rect 1290 2330 1385 2370
rect 1315 2310 1385 2330
rect 1445 2330 1540 2370
rect 1445 2310 1515 2330
rect 1230 2295 1286 2301
rect 1230 2235 1234 2295
rect 1315 2285 1515 2310
rect 1570 2301 1600 2489
rect 1544 2295 1600 2301
rect 1286 2235 1544 2255
rect 1596 2235 1600 2295
rect 1230 2225 1600 2235
rect 1630 2555 2000 2565
rect 1630 2495 1634 2555
rect 1686 2535 1944 2555
rect 1630 2489 1686 2495
rect 1630 2301 1660 2489
rect 1715 2480 1915 2505
rect 1996 2495 2000 2555
rect 1944 2489 2000 2495
rect 1715 2460 1785 2480
rect 1690 2420 1785 2460
rect 1845 2460 1915 2480
rect 1845 2420 1940 2460
rect 1690 2370 1940 2420
rect 1690 2330 1785 2370
rect 1715 2310 1785 2330
rect 1845 2330 1940 2370
rect 1845 2310 1915 2330
rect 1630 2295 1686 2301
rect 1630 2235 1634 2295
rect 1715 2285 1915 2310
rect 1970 2301 2000 2489
rect 1944 2295 2000 2301
rect 1686 2235 1944 2255
rect 1996 2235 2000 2295
rect 1630 2225 2000 2235
rect 2030 2555 2400 2565
rect 2030 2495 2034 2555
rect 2086 2535 2344 2555
rect 2030 2489 2086 2495
rect 2030 2301 2060 2489
rect 2115 2480 2315 2505
rect 2396 2495 2400 2555
rect 2344 2489 2400 2495
rect 2115 2460 2185 2480
rect 2090 2420 2185 2460
rect 2245 2460 2315 2480
rect 2245 2420 2340 2460
rect 2090 2370 2340 2420
rect 2090 2330 2185 2370
rect 2115 2310 2185 2330
rect 2245 2330 2340 2370
rect 2245 2310 2315 2330
rect 2030 2295 2086 2301
rect 2030 2235 2034 2295
rect 2115 2285 2315 2310
rect 2370 2301 2400 2489
rect 2344 2295 2400 2301
rect 2086 2235 2344 2255
rect 2396 2235 2400 2295
rect 2030 2225 2400 2235
rect 2430 2555 2800 2565
rect 2430 2495 2434 2555
rect 2486 2535 2744 2555
rect 2430 2489 2486 2495
rect 2430 2301 2460 2489
rect 2515 2480 2715 2505
rect 2796 2495 2800 2555
rect 2744 2489 2800 2495
rect 2515 2460 2585 2480
rect 2490 2420 2585 2460
rect 2645 2460 2715 2480
rect 2645 2420 2740 2460
rect 2490 2370 2740 2420
rect 2490 2330 2585 2370
rect 2515 2310 2585 2330
rect 2645 2330 2740 2370
rect 2645 2310 2715 2330
rect 2430 2295 2486 2301
rect 2430 2235 2434 2295
rect 2515 2285 2715 2310
rect 2770 2301 2800 2489
rect 2744 2295 2800 2301
rect 2486 2235 2744 2255
rect 2796 2235 2800 2295
rect 2430 2225 2800 2235
rect 2830 2555 3200 2565
rect 2830 2495 2834 2555
rect 2886 2535 3144 2555
rect 2830 2489 2886 2495
rect 2830 2301 2860 2489
rect 2915 2480 3115 2505
rect 3196 2495 3200 2555
rect 3144 2489 3200 2495
rect 2915 2460 2985 2480
rect 2890 2420 2985 2460
rect 3045 2460 3115 2480
rect 3045 2420 3140 2460
rect 2890 2370 3140 2420
rect 2890 2330 2985 2370
rect 2915 2310 2985 2330
rect 3045 2330 3140 2370
rect 3045 2310 3115 2330
rect 2830 2295 2886 2301
rect 2830 2235 2834 2295
rect 2915 2285 3115 2310
rect 3170 2301 3200 2489
rect 3144 2295 3200 2301
rect 2886 2235 3144 2255
rect 3196 2235 3200 2295
rect 2830 2225 3200 2235
rect 3230 2555 3600 2565
rect 3230 2495 3234 2555
rect 3286 2535 3544 2555
rect 3230 2489 3286 2495
rect 3230 2301 3260 2489
rect 3315 2480 3515 2505
rect 3596 2495 3600 2555
rect 3544 2489 3600 2495
rect 3315 2460 3385 2480
rect 3290 2420 3385 2460
rect 3445 2460 3515 2480
rect 3445 2420 3540 2460
rect 3290 2370 3540 2420
rect 3290 2330 3385 2370
rect 3315 2310 3385 2330
rect 3445 2330 3540 2370
rect 3445 2310 3515 2330
rect 3230 2295 3286 2301
rect 3230 2235 3234 2295
rect 3315 2285 3515 2310
rect 3570 2301 3600 2489
rect 3544 2295 3600 2301
rect 3286 2235 3544 2255
rect 3596 2235 3600 2295
rect 3230 2225 3600 2235
rect 3630 2555 4000 2565
rect 3630 2495 3634 2555
rect 3686 2535 3944 2555
rect 3630 2489 3686 2495
rect 3630 2301 3660 2489
rect 3715 2480 3915 2505
rect 3996 2495 4000 2555
rect 3944 2489 4000 2495
rect 3715 2460 3785 2480
rect 3690 2420 3785 2460
rect 3845 2460 3915 2480
rect 3845 2420 3940 2460
rect 3690 2370 3940 2420
rect 3690 2330 3785 2370
rect 3715 2310 3785 2330
rect 3845 2330 3940 2370
rect 3845 2310 3915 2330
rect 3630 2295 3686 2301
rect 3630 2235 3634 2295
rect 3715 2285 3915 2310
rect 3970 2301 4000 2489
rect 3944 2295 4000 2301
rect 3686 2235 3944 2255
rect 3996 2235 4000 2295
rect 3630 2225 4000 2235
rect 4030 2555 4400 2565
rect 4030 2495 4034 2555
rect 4086 2535 4344 2555
rect 4030 2489 4086 2495
rect 4030 2301 4060 2489
rect 4115 2480 4315 2505
rect 4396 2495 4400 2555
rect 4344 2489 4400 2495
rect 4115 2460 4185 2480
rect 4090 2420 4185 2460
rect 4245 2460 4315 2480
rect 4245 2420 4340 2460
rect 4090 2370 4340 2420
rect 4090 2330 4185 2370
rect 4115 2310 4185 2330
rect 4245 2330 4340 2370
rect 4245 2310 4315 2330
rect 4030 2295 4086 2301
rect 4030 2235 4034 2295
rect 4115 2285 4315 2310
rect 4370 2301 4400 2489
rect 4344 2295 4400 2301
rect 4086 2235 4344 2255
rect 4396 2235 4400 2295
rect 4030 2225 4400 2235
rect 4430 2555 4800 2565
rect 4430 2495 4434 2555
rect 4486 2535 4744 2555
rect 4430 2489 4486 2495
rect 4430 2301 4460 2489
rect 4515 2480 4715 2505
rect 4796 2495 4800 2555
rect 4744 2489 4800 2495
rect 4515 2460 4585 2480
rect 4490 2420 4585 2460
rect 4645 2460 4715 2480
rect 4645 2420 4740 2460
rect 4490 2370 4740 2420
rect 4490 2330 4585 2370
rect 4515 2310 4585 2330
rect 4645 2330 4740 2370
rect 4645 2310 4715 2330
rect 4430 2295 4486 2301
rect 4430 2235 4434 2295
rect 4515 2285 4715 2310
rect 4770 2301 4800 2489
rect 4744 2295 4800 2301
rect 4486 2235 4744 2255
rect 4796 2235 4800 2295
rect 4430 2225 4800 2235
rect 4830 2555 5200 2565
rect 4830 2495 4834 2555
rect 4886 2535 5144 2555
rect 4830 2489 4886 2495
rect 4830 2301 4860 2489
rect 4915 2480 5115 2505
rect 5196 2495 5200 2555
rect 5144 2489 5200 2495
rect 4915 2460 4985 2480
rect 4890 2420 4985 2460
rect 5045 2460 5115 2480
rect 5045 2420 5140 2460
rect 4890 2370 5140 2420
rect 4890 2330 4985 2370
rect 4915 2310 4985 2330
rect 5045 2330 5140 2370
rect 5045 2310 5115 2330
rect 4830 2295 4886 2301
rect 4830 2235 4834 2295
rect 4915 2285 5115 2310
rect 5170 2301 5200 2489
rect 5144 2295 5200 2301
rect 4886 2235 5144 2255
rect 5196 2235 5200 2295
rect 4830 2225 5200 2235
rect 5230 2555 5600 2565
rect 5230 2495 5234 2555
rect 5286 2535 5544 2555
rect 5230 2489 5286 2495
rect 5230 2301 5260 2489
rect 5315 2480 5515 2505
rect 5596 2495 5600 2555
rect 5544 2489 5600 2495
rect 5315 2460 5385 2480
rect 5290 2420 5385 2460
rect 5445 2460 5515 2480
rect 5445 2420 5540 2460
rect 5290 2370 5540 2420
rect 5290 2330 5385 2370
rect 5315 2310 5385 2330
rect 5445 2330 5540 2370
rect 5445 2310 5515 2330
rect 5230 2295 5286 2301
rect 5230 2235 5234 2295
rect 5315 2285 5515 2310
rect 5570 2301 5600 2489
rect 5544 2295 5600 2301
rect 5286 2235 5544 2255
rect 5596 2235 5600 2295
rect 5230 2225 5600 2235
rect 5630 2555 6000 2565
rect 5630 2495 5634 2555
rect 5686 2535 5944 2555
rect 5630 2489 5686 2495
rect 5630 2301 5660 2489
rect 5715 2480 5915 2505
rect 5996 2495 6000 2555
rect 5944 2489 6000 2495
rect 5715 2460 5785 2480
rect 5690 2420 5785 2460
rect 5845 2460 5915 2480
rect 5845 2420 5940 2460
rect 5690 2370 5940 2420
rect 5690 2330 5785 2370
rect 5715 2310 5785 2330
rect 5845 2330 5940 2370
rect 5845 2310 5915 2330
rect 5630 2295 5686 2301
rect 5630 2235 5634 2295
rect 5715 2285 5915 2310
rect 5970 2301 6000 2489
rect 5944 2295 6000 2301
rect 5686 2235 5944 2255
rect 5996 2235 6000 2295
rect 5630 2225 6000 2235
rect 6030 2555 6400 2565
rect 6030 2495 6034 2555
rect 6086 2535 6344 2555
rect 6030 2489 6086 2495
rect 6030 2301 6060 2489
rect 6115 2480 6315 2505
rect 6396 2495 6400 2555
rect 6344 2489 6400 2495
rect 6115 2460 6185 2480
rect 6090 2420 6185 2460
rect 6245 2460 6315 2480
rect 6245 2420 6340 2460
rect 6090 2370 6340 2420
rect 6090 2330 6185 2370
rect 6115 2310 6185 2330
rect 6245 2330 6340 2370
rect 6245 2310 6315 2330
rect 6030 2295 6086 2301
rect 6030 2235 6034 2295
rect 6115 2285 6315 2310
rect 6370 2301 6400 2489
rect 6344 2295 6400 2301
rect 6086 2235 6344 2255
rect 6396 2235 6400 2295
rect 6030 2225 6400 2235
rect 6430 2555 6800 2565
rect 6430 2495 6434 2555
rect 6486 2535 6744 2555
rect 6430 2489 6486 2495
rect 6430 2301 6460 2489
rect 6515 2480 6715 2505
rect 6796 2495 6800 2555
rect 6744 2489 6800 2495
rect 6515 2460 6585 2480
rect 6490 2420 6585 2460
rect 6645 2460 6715 2480
rect 6645 2420 6740 2460
rect 6490 2370 6740 2420
rect 6490 2330 6585 2370
rect 6515 2310 6585 2330
rect 6645 2330 6740 2370
rect 6645 2310 6715 2330
rect 6430 2295 6486 2301
rect 6430 2235 6434 2295
rect 6515 2285 6715 2310
rect 6770 2301 6800 2489
rect 6744 2295 6800 2301
rect 6486 2235 6744 2255
rect 6796 2235 6800 2295
rect 6430 2225 6800 2235
rect 6830 2555 7200 2565
rect 6830 2495 6834 2555
rect 6886 2535 7144 2555
rect 6830 2489 6886 2495
rect 6830 2301 6860 2489
rect 6915 2480 7115 2505
rect 7196 2495 7200 2555
rect 7144 2489 7200 2495
rect 6915 2460 6985 2480
rect 6890 2420 6985 2460
rect 7045 2460 7115 2480
rect 7045 2420 7140 2460
rect 6890 2370 7140 2420
rect 6890 2330 6985 2370
rect 6915 2310 6985 2330
rect 7045 2330 7140 2370
rect 7045 2310 7115 2330
rect 6830 2295 6886 2301
rect 6830 2235 6834 2295
rect 6915 2285 7115 2310
rect 7170 2301 7200 2489
rect 7144 2295 7200 2301
rect 6886 2235 7144 2255
rect 7196 2235 7200 2295
rect 6830 2225 7200 2235
rect 7230 2555 7600 2565
rect 7230 2495 7234 2555
rect 7286 2535 7544 2555
rect 7230 2489 7286 2495
rect 7230 2301 7260 2489
rect 7315 2480 7515 2505
rect 7596 2495 7600 2555
rect 7544 2489 7600 2495
rect 7315 2460 7385 2480
rect 7290 2420 7385 2460
rect 7445 2460 7515 2480
rect 7445 2420 7540 2460
rect 7290 2370 7540 2420
rect 7290 2330 7385 2370
rect 7315 2310 7385 2330
rect 7445 2330 7540 2370
rect 7445 2310 7515 2330
rect 7230 2295 7286 2301
rect 7230 2235 7234 2295
rect 7315 2285 7515 2310
rect 7570 2301 7600 2489
rect 7544 2295 7600 2301
rect 7286 2235 7544 2255
rect 7596 2235 7600 2295
rect 7230 2225 7600 2235
rect 7630 2555 8000 2565
rect 7630 2495 7634 2555
rect 7686 2535 7944 2555
rect 7630 2489 7686 2495
rect 7630 2301 7660 2489
rect 7715 2480 7915 2505
rect 7996 2495 8000 2555
rect 7944 2489 8000 2495
rect 7715 2460 7785 2480
rect 7690 2420 7785 2460
rect 7845 2460 7915 2480
rect 7845 2420 7940 2460
rect 7690 2370 7940 2420
rect 7690 2330 7785 2370
rect 7715 2310 7785 2330
rect 7845 2330 7940 2370
rect 7845 2310 7915 2330
rect 7630 2295 7686 2301
rect 7630 2235 7634 2295
rect 7715 2285 7915 2310
rect 7970 2301 8000 2489
rect 7944 2295 8000 2301
rect 7686 2235 7944 2255
rect 7996 2235 8000 2295
rect 7630 2225 8000 2235
rect 8030 2555 8400 2565
rect 8030 2495 8034 2555
rect 8086 2535 8344 2555
rect 8030 2489 8086 2495
rect 8030 2301 8060 2489
rect 8115 2480 8315 2505
rect 8396 2495 8400 2555
rect 8344 2489 8400 2495
rect 8115 2460 8185 2480
rect 8090 2420 8185 2460
rect 8245 2460 8315 2480
rect 8245 2420 8340 2460
rect 8090 2370 8340 2420
rect 8090 2330 8185 2370
rect 8115 2310 8185 2330
rect 8245 2330 8340 2370
rect 8245 2310 8315 2330
rect 8030 2295 8086 2301
rect 8030 2235 8034 2295
rect 8115 2285 8315 2310
rect 8370 2301 8400 2489
rect 8344 2295 8400 2301
rect 8086 2235 8344 2255
rect 8396 2235 8400 2295
rect 8030 2225 8400 2235
rect 8430 2555 8800 2565
rect 8430 2495 8434 2555
rect 8486 2535 8744 2555
rect 8430 2489 8486 2495
rect 8430 2301 8460 2489
rect 8515 2480 8715 2505
rect 8796 2495 8800 2555
rect 8744 2489 8800 2495
rect 8515 2460 8585 2480
rect 8490 2420 8585 2460
rect 8645 2460 8715 2480
rect 8645 2420 8740 2460
rect 8490 2370 8740 2420
rect 8490 2330 8585 2370
rect 8515 2310 8585 2330
rect 8645 2330 8740 2370
rect 8645 2310 8715 2330
rect 8430 2295 8486 2301
rect 8430 2235 8434 2295
rect 8515 2285 8715 2310
rect 8770 2301 8800 2489
rect 8744 2295 8800 2301
rect 8486 2235 8744 2255
rect 8796 2235 8800 2295
rect 8430 2225 8800 2235
rect 8830 2555 9200 2565
rect 8830 2495 8834 2555
rect 8886 2535 9144 2555
rect 8830 2489 8886 2495
rect 8830 2301 8860 2489
rect 8915 2480 9115 2505
rect 9196 2495 9200 2555
rect 9144 2489 9200 2495
rect 8915 2460 8985 2480
rect 8890 2420 8985 2460
rect 9045 2460 9115 2480
rect 9045 2420 9140 2460
rect 8890 2370 9140 2420
rect 8890 2330 8985 2370
rect 8915 2310 8985 2330
rect 9045 2330 9140 2370
rect 9045 2310 9115 2330
rect 8830 2295 8886 2301
rect 8830 2235 8834 2295
rect 8915 2285 9115 2310
rect 9170 2301 9200 2489
rect 9144 2295 9200 2301
rect 8886 2235 9144 2255
rect 9196 2235 9200 2295
rect 8830 2225 9200 2235
rect 9230 2555 9600 2565
rect 9230 2495 9234 2555
rect 9286 2535 9544 2555
rect 9230 2489 9286 2495
rect 9230 2301 9260 2489
rect 9315 2480 9515 2505
rect 9596 2495 9600 2555
rect 9544 2489 9600 2495
rect 9315 2460 9385 2480
rect 9290 2420 9385 2460
rect 9445 2460 9515 2480
rect 9445 2420 9540 2460
rect 9290 2370 9540 2420
rect 9290 2330 9385 2370
rect 9315 2310 9385 2330
rect 9445 2330 9540 2370
rect 9445 2310 9515 2330
rect 9230 2295 9286 2301
rect 9230 2235 9234 2295
rect 9315 2285 9515 2310
rect 9570 2301 9600 2489
rect 9544 2295 9600 2301
rect 9286 2235 9544 2255
rect 9596 2235 9600 2295
rect 9230 2225 9600 2235
rect 9630 2555 10000 2565
rect 9630 2495 9634 2555
rect 9686 2535 9944 2555
rect 9630 2489 9686 2495
rect 9630 2301 9660 2489
rect 9715 2480 9915 2505
rect 9996 2495 10000 2555
rect 9944 2489 10000 2495
rect 9715 2460 9785 2480
rect 9690 2420 9785 2460
rect 9845 2460 9915 2480
rect 9845 2420 9940 2460
rect 9690 2370 9940 2420
rect 9690 2330 9785 2370
rect 9715 2310 9785 2330
rect 9845 2330 9940 2370
rect 9845 2310 9915 2330
rect 9630 2295 9686 2301
rect 9630 2235 9634 2295
rect 9715 2285 9915 2310
rect 9970 2301 10000 2489
rect 9944 2295 10000 2301
rect 9686 2235 9944 2255
rect 9996 2235 10000 2295
rect 9630 2225 10000 2235
rect 10030 2555 10400 2565
rect 10030 2495 10034 2555
rect 10086 2535 10344 2555
rect 10030 2489 10086 2495
rect 10030 2301 10060 2489
rect 10115 2480 10315 2505
rect 10396 2495 10400 2555
rect 10344 2489 10400 2495
rect 10115 2460 10185 2480
rect 10090 2420 10185 2460
rect 10245 2460 10315 2480
rect 10245 2420 10340 2460
rect 10090 2370 10340 2420
rect 10090 2330 10185 2370
rect 10115 2310 10185 2330
rect 10245 2330 10340 2370
rect 10245 2310 10315 2330
rect 10030 2295 10086 2301
rect 10030 2235 10034 2295
rect 10115 2285 10315 2310
rect 10370 2301 10400 2489
rect 10344 2295 10400 2301
rect 10086 2235 10344 2255
rect 10396 2235 10400 2295
rect 10030 2225 10400 2235
rect 10430 2555 10800 2565
rect 10430 2495 10434 2555
rect 10486 2535 10744 2555
rect 10430 2489 10486 2495
rect 10430 2301 10460 2489
rect 10515 2480 10715 2505
rect 10796 2495 10800 2555
rect 10744 2489 10800 2495
rect 10515 2460 10585 2480
rect 10490 2420 10585 2460
rect 10645 2460 10715 2480
rect 10645 2420 10740 2460
rect 10490 2370 10740 2420
rect 10490 2330 10585 2370
rect 10515 2310 10585 2330
rect 10645 2330 10740 2370
rect 10645 2310 10715 2330
rect 10430 2295 10486 2301
rect 10430 2235 10434 2295
rect 10515 2285 10715 2310
rect 10770 2301 10800 2489
rect 10744 2295 10800 2301
rect 10486 2235 10744 2255
rect 10796 2235 10800 2295
rect 10430 2225 10800 2235
rect 10830 2555 11200 2565
rect 10830 2495 10834 2555
rect 10886 2535 11144 2555
rect 10830 2489 10886 2495
rect 10830 2301 10860 2489
rect 10915 2480 11115 2505
rect 11196 2495 11200 2555
rect 11144 2489 11200 2495
rect 10915 2460 10985 2480
rect 10890 2420 10985 2460
rect 11045 2460 11115 2480
rect 11045 2420 11140 2460
rect 10890 2370 11140 2420
rect 10890 2330 10985 2370
rect 10915 2310 10985 2330
rect 11045 2330 11140 2370
rect 11045 2310 11115 2330
rect 10830 2295 10886 2301
rect 10830 2235 10834 2295
rect 10915 2285 11115 2310
rect 11170 2301 11200 2489
rect 11144 2295 11200 2301
rect 10886 2235 11144 2255
rect 11196 2235 11200 2295
rect 10830 2225 11200 2235
rect 11230 2555 11600 2565
rect 11230 2495 11234 2555
rect 11286 2535 11544 2555
rect 11230 2489 11286 2495
rect 11230 2301 11260 2489
rect 11315 2480 11515 2505
rect 11596 2495 11600 2555
rect 11544 2489 11600 2495
rect 11315 2460 11385 2480
rect 11290 2420 11385 2460
rect 11445 2460 11515 2480
rect 11445 2420 11540 2460
rect 11290 2370 11540 2420
rect 11290 2330 11385 2370
rect 11315 2310 11385 2330
rect 11445 2330 11540 2370
rect 11445 2310 11515 2330
rect 11230 2295 11286 2301
rect 11230 2235 11234 2295
rect 11315 2285 11515 2310
rect 11570 2301 11600 2489
rect 11544 2295 11600 2301
rect 11286 2235 11544 2255
rect 11596 2235 11600 2295
rect 11230 2225 11600 2235
rect 11630 2555 12000 2565
rect 11630 2495 11634 2555
rect 11686 2535 11944 2555
rect 11630 2489 11686 2495
rect 11630 2301 11660 2489
rect 11715 2480 11915 2505
rect 11996 2495 12000 2555
rect 11944 2489 12000 2495
rect 11715 2460 11785 2480
rect 11690 2420 11785 2460
rect 11845 2460 11915 2480
rect 11845 2420 11940 2460
rect 11690 2370 11940 2420
rect 11690 2330 11785 2370
rect 11715 2310 11785 2330
rect 11845 2330 11940 2370
rect 11845 2310 11915 2330
rect 11630 2295 11686 2301
rect 11630 2235 11634 2295
rect 11715 2285 11915 2310
rect 11970 2301 12000 2489
rect 11944 2295 12000 2301
rect 11686 2235 11944 2255
rect 11996 2235 12000 2295
rect 11630 2225 12000 2235
rect 12030 2555 12400 2565
rect 12030 2495 12034 2555
rect 12086 2535 12344 2555
rect 12030 2489 12086 2495
rect 12030 2301 12060 2489
rect 12115 2480 12315 2505
rect 12396 2495 12400 2555
rect 12344 2489 12400 2495
rect 12115 2460 12185 2480
rect 12090 2420 12185 2460
rect 12245 2460 12315 2480
rect 12245 2420 12340 2460
rect 12090 2370 12340 2420
rect 12090 2330 12185 2370
rect 12115 2310 12185 2330
rect 12245 2330 12340 2370
rect 12245 2310 12315 2330
rect 12030 2295 12086 2301
rect 12030 2235 12034 2295
rect 12115 2285 12315 2310
rect 12370 2301 12400 2489
rect 12344 2295 12400 2301
rect 12086 2235 12344 2255
rect 12396 2235 12400 2295
rect 12030 2225 12400 2235
rect 12430 2555 12800 2565
rect 12430 2495 12434 2555
rect 12486 2535 12744 2555
rect 12430 2489 12486 2495
rect 12430 2301 12460 2489
rect 12515 2480 12715 2505
rect 12796 2495 12800 2555
rect 12744 2489 12800 2495
rect 12515 2460 12585 2480
rect 12490 2420 12585 2460
rect 12645 2460 12715 2480
rect 12645 2420 12740 2460
rect 12490 2370 12740 2420
rect 12490 2330 12585 2370
rect 12515 2310 12585 2330
rect 12645 2330 12740 2370
rect 12645 2310 12715 2330
rect 12430 2295 12486 2301
rect 12430 2235 12434 2295
rect 12515 2285 12715 2310
rect 12770 2301 12800 2489
rect 12744 2295 12800 2301
rect 12486 2235 12744 2255
rect 12796 2235 12800 2295
rect 12430 2225 12800 2235
rect 12830 2555 13200 2565
rect 12830 2495 12834 2555
rect 12886 2535 13144 2555
rect 12830 2489 12886 2495
rect 12830 2301 12860 2489
rect 12915 2480 13115 2505
rect 13196 2495 13200 2555
rect 13144 2489 13200 2495
rect 12915 2460 12985 2480
rect 12890 2420 12985 2460
rect 13045 2460 13115 2480
rect 13045 2420 13140 2460
rect 12890 2370 13140 2420
rect 12890 2330 12985 2370
rect 12915 2310 12985 2330
rect 13045 2330 13140 2370
rect 13045 2310 13115 2330
rect 12830 2295 12886 2301
rect 12830 2235 12834 2295
rect 12915 2285 13115 2310
rect 13170 2301 13200 2489
rect 13144 2295 13200 2301
rect 12886 2235 13144 2255
rect 13196 2235 13200 2295
rect 12830 2225 13200 2235
rect -370 2185 0 2195
rect -370 2125 -366 2185
rect -314 2165 -56 2185
rect -370 2119 -314 2125
rect -370 1931 -340 2119
rect -285 2110 -85 2135
rect -4 2125 0 2185
rect -56 2119 0 2125
rect -285 2090 -215 2110
rect -310 2050 -215 2090
rect -155 2090 -85 2110
rect -155 2050 -60 2090
rect -310 2000 -60 2050
rect -310 1960 -215 2000
rect -285 1940 -215 1960
rect -155 1960 -60 2000
rect -155 1940 -85 1960
rect -370 1925 -314 1931
rect -370 1865 -366 1925
rect -285 1915 -85 1940
rect -30 1931 0 2119
rect -56 1925 0 1931
rect -314 1865 -56 1885
rect -4 1865 0 1925
rect -370 1855 0 1865
rect 30 2185 400 2195
rect 30 2125 34 2185
rect 86 2165 344 2185
rect 30 2119 86 2125
rect 30 1931 60 2119
rect 115 2110 315 2135
rect 396 2125 400 2185
rect 344 2119 400 2125
rect 115 2090 185 2110
rect 90 2050 185 2090
rect 245 2090 315 2110
rect 245 2050 340 2090
rect 90 2000 340 2050
rect 90 1960 185 2000
rect 115 1940 185 1960
rect 245 1960 340 2000
rect 245 1940 315 1960
rect 30 1925 86 1931
rect 30 1865 34 1925
rect 115 1915 315 1940
rect 370 1931 400 2119
rect 344 1925 400 1931
rect 86 1865 344 1885
rect 396 1865 400 1925
rect 30 1855 400 1865
rect 430 2185 800 2195
rect 430 2125 434 2185
rect 486 2165 744 2185
rect 430 2119 486 2125
rect 430 1931 460 2119
rect 515 2110 715 2135
rect 796 2125 800 2185
rect 744 2119 800 2125
rect 515 2090 585 2110
rect 490 2050 585 2090
rect 645 2090 715 2110
rect 645 2050 740 2090
rect 490 2000 740 2050
rect 490 1960 585 2000
rect 515 1940 585 1960
rect 645 1960 740 2000
rect 645 1940 715 1960
rect 430 1925 486 1931
rect 430 1865 434 1925
rect 515 1915 715 1940
rect 770 1931 800 2119
rect 744 1925 800 1931
rect 486 1865 744 1885
rect 796 1865 800 1925
rect 430 1855 800 1865
rect 830 2185 1200 2195
rect 830 2125 834 2185
rect 886 2165 1144 2185
rect 830 2119 886 2125
rect 830 1931 860 2119
rect 915 2110 1115 2135
rect 1196 2125 1200 2185
rect 1144 2119 1200 2125
rect 915 2090 985 2110
rect 890 2050 985 2090
rect 1045 2090 1115 2110
rect 1045 2050 1140 2090
rect 890 2000 1140 2050
rect 890 1960 985 2000
rect 915 1940 985 1960
rect 1045 1960 1140 2000
rect 1045 1940 1115 1960
rect 830 1925 886 1931
rect 830 1865 834 1925
rect 915 1915 1115 1940
rect 1170 1931 1200 2119
rect 1144 1925 1200 1931
rect 886 1865 1144 1885
rect 1196 1865 1200 1925
rect 830 1855 1200 1865
rect 1230 2185 1600 2195
rect 1230 2125 1234 2185
rect 1286 2165 1544 2185
rect 1230 2119 1286 2125
rect 1230 1931 1260 2119
rect 1315 2110 1515 2135
rect 1596 2125 1600 2185
rect 1544 2119 1600 2125
rect 1315 2090 1385 2110
rect 1290 2050 1385 2090
rect 1445 2090 1515 2110
rect 1445 2050 1540 2090
rect 1290 2000 1540 2050
rect 1290 1960 1385 2000
rect 1315 1940 1385 1960
rect 1445 1960 1540 2000
rect 1445 1940 1515 1960
rect 1230 1925 1286 1931
rect 1230 1865 1234 1925
rect 1315 1915 1515 1940
rect 1570 1931 1600 2119
rect 1544 1925 1600 1931
rect 1286 1865 1544 1885
rect 1596 1865 1600 1925
rect 1230 1855 1600 1865
rect 1630 2185 2000 2195
rect 1630 2125 1634 2185
rect 1686 2165 1944 2185
rect 1630 2119 1686 2125
rect 1630 1931 1660 2119
rect 1715 2110 1915 2135
rect 1996 2125 2000 2185
rect 1944 2119 2000 2125
rect 1715 2090 1785 2110
rect 1690 2050 1785 2090
rect 1845 2090 1915 2110
rect 1845 2050 1940 2090
rect 1690 2000 1940 2050
rect 1690 1960 1785 2000
rect 1715 1940 1785 1960
rect 1845 1960 1940 2000
rect 1845 1940 1915 1960
rect 1630 1925 1686 1931
rect 1630 1865 1634 1925
rect 1715 1915 1915 1940
rect 1970 1931 2000 2119
rect 1944 1925 2000 1931
rect 1686 1865 1944 1885
rect 1996 1865 2000 1925
rect 1630 1855 2000 1865
rect 2030 2185 2400 2195
rect 2030 2125 2034 2185
rect 2086 2165 2344 2185
rect 2030 2119 2086 2125
rect 2030 1931 2060 2119
rect 2115 2110 2315 2135
rect 2396 2125 2400 2185
rect 2344 2119 2400 2125
rect 2115 2090 2185 2110
rect 2090 2050 2185 2090
rect 2245 2090 2315 2110
rect 2245 2050 2340 2090
rect 2090 2000 2340 2050
rect 2090 1960 2185 2000
rect 2115 1940 2185 1960
rect 2245 1960 2340 2000
rect 2245 1940 2315 1960
rect 2030 1925 2086 1931
rect 2030 1865 2034 1925
rect 2115 1915 2315 1940
rect 2370 1931 2400 2119
rect 2344 1925 2400 1931
rect 2086 1865 2344 1885
rect 2396 1865 2400 1925
rect 2030 1855 2400 1865
rect 2430 2185 2800 2195
rect 2430 2125 2434 2185
rect 2486 2165 2744 2185
rect 2430 2119 2486 2125
rect 2430 1931 2460 2119
rect 2515 2110 2715 2135
rect 2796 2125 2800 2185
rect 2744 2119 2800 2125
rect 2515 2090 2585 2110
rect 2490 2050 2585 2090
rect 2645 2090 2715 2110
rect 2645 2050 2740 2090
rect 2490 2000 2740 2050
rect 2490 1960 2585 2000
rect 2515 1940 2585 1960
rect 2645 1960 2740 2000
rect 2645 1940 2715 1960
rect 2430 1925 2486 1931
rect 2430 1865 2434 1925
rect 2515 1915 2715 1940
rect 2770 1931 2800 2119
rect 2744 1925 2800 1931
rect 2486 1865 2744 1885
rect 2796 1865 2800 1925
rect 2430 1855 2800 1865
rect 2830 2185 3200 2195
rect 2830 2125 2834 2185
rect 2886 2165 3144 2185
rect 2830 2119 2886 2125
rect 2830 1931 2860 2119
rect 2915 2110 3115 2135
rect 3196 2125 3200 2185
rect 3144 2119 3200 2125
rect 2915 2090 2985 2110
rect 2890 2050 2985 2090
rect 3045 2090 3115 2110
rect 3045 2050 3140 2090
rect 2890 2000 3140 2050
rect 2890 1960 2985 2000
rect 2915 1940 2985 1960
rect 3045 1960 3140 2000
rect 3045 1940 3115 1960
rect 2830 1925 2886 1931
rect 2830 1865 2834 1925
rect 2915 1915 3115 1940
rect 3170 1931 3200 2119
rect 3144 1925 3200 1931
rect 2886 1865 3144 1885
rect 3196 1865 3200 1925
rect 2830 1855 3200 1865
rect 3230 2185 3600 2195
rect 3230 2125 3234 2185
rect 3286 2165 3544 2185
rect 3230 2119 3286 2125
rect 3230 1931 3260 2119
rect 3315 2110 3515 2135
rect 3596 2125 3600 2185
rect 3544 2119 3600 2125
rect 3315 2090 3385 2110
rect 3290 2050 3385 2090
rect 3445 2090 3515 2110
rect 3445 2050 3540 2090
rect 3290 2000 3540 2050
rect 3290 1960 3385 2000
rect 3315 1940 3385 1960
rect 3445 1960 3540 2000
rect 3445 1940 3515 1960
rect 3230 1925 3286 1931
rect 3230 1865 3234 1925
rect 3315 1915 3515 1940
rect 3570 1931 3600 2119
rect 3544 1925 3600 1931
rect 3286 1865 3544 1885
rect 3596 1865 3600 1925
rect 3230 1855 3600 1865
rect 3630 2185 4000 2195
rect 3630 2125 3634 2185
rect 3686 2165 3944 2185
rect 3630 2119 3686 2125
rect 3630 1931 3660 2119
rect 3715 2110 3915 2135
rect 3996 2125 4000 2185
rect 3944 2119 4000 2125
rect 3715 2090 3785 2110
rect 3690 2050 3785 2090
rect 3845 2090 3915 2110
rect 3845 2050 3940 2090
rect 3690 2000 3940 2050
rect 3690 1960 3785 2000
rect 3715 1940 3785 1960
rect 3845 1960 3940 2000
rect 3845 1940 3915 1960
rect 3630 1925 3686 1931
rect 3630 1865 3634 1925
rect 3715 1915 3915 1940
rect 3970 1931 4000 2119
rect 3944 1925 4000 1931
rect 3686 1865 3944 1885
rect 3996 1865 4000 1925
rect 3630 1855 4000 1865
rect 4030 2185 4400 2195
rect 4030 2125 4034 2185
rect 4086 2165 4344 2185
rect 4030 2119 4086 2125
rect 4030 1931 4060 2119
rect 4115 2110 4315 2135
rect 4396 2125 4400 2185
rect 4344 2119 4400 2125
rect 4115 2090 4185 2110
rect 4090 2050 4185 2090
rect 4245 2090 4315 2110
rect 4245 2050 4340 2090
rect 4090 2000 4340 2050
rect 4090 1960 4185 2000
rect 4115 1940 4185 1960
rect 4245 1960 4340 2000
rect 4245 1940 4315 1960
rect 4030 1925 4086 1931
rect 4030 1865 4034 1925
rect 4115 1915 4315 1940
rect 4370 1931 4400 2119
rect 4344 1925 4400 1931
rect 4086 1865 4344 1885
rect 4396 1865 4400 1925
rect 4030 1855 4400 1865
rect 4430 2185 4800 2195
rect 4430 2125 4434 2185
rect 4486 2165 4744 2185
rect 4430 2119 4486 2125
rect 4430 1931 4460 2119
rect 4515 2110 4715 2135
rect 4796 2125 4800 2185
rect 4744 2119 4800 2125
rect 4515 2090 4585 2110
rect 4490 2050 4585 2090
rect 4645 2090 4715 2110
rect 4645 2050 4740 2090
rect 4490 2000 4740 2050
rect 4490 1960 4585 2000
rect 4515 1940 4585 1960
rect 4645 1960 4740 2000
rect 4645 1940 4715 1960
rect 4430 1925 4486 1931
rect 4430 1865 4434 1925
rect 4515 1915 4715 1940
rect 4770 1931 4800 2119
rect 4744 1925 4800 1931
rect 4486 1865 4744 1885
rect 4796 1865 4800 1925
rect 4430 1855 4800 1865
rect 4830 2185 5200 2195
rect 4830 2125 4834 2185
rect 4886 2165 5144 2185
rect 4830 2119 4886 2125
rect 4830 1931 4860 2119
rect 4915 2110 5115 2135
rect 5196 2125 5200 2185
rect 5144 2119 5200 2125
rect 4915 2090 4985 2110
rect 4890 2050 4985 2090
rect 5045 2090 5115 2110
rect 5045 2050 5140 2090
rect 4890 2000 5140 2050
rect 4890 1960 4985 2000
rect 4915 1940 4985 1960
rect 5045 1960 5140 2000
rect 5045 1940 5115 1960
rect 4830 1925 4886 1931
rect 4830 1865 4834 1925
rect 4915 1915 5115 1940
rect 5170 1931 5200 2119
rect 5144 1925 5200 1931
rect 4886 1865 5144 1885
rect 5196 1865 5200 1925
rect 4830 1855 5200 1865
rect 5230 2185 5600 2195
rect 5230 2125 5234 2185
rect 5286 2165 5544 2185
rect 5230 2119 5286 2125
rect 5230 1931 5260 2119
rect 5315 2110 5515 2135
rect 5596 2125 5600 2185
rect 5544 2119 5600 2125
rect 5315 2090 5385 2110
rect 5290 2050 5385 2090
rect 5445 2090 5515 2110
rect 5445 2050 5540 2090
rect 5290 2000 5540 2050
rect 5290 1960 5385 2000
rect 5315 1940 5385 1960
rect 5445 1960 5540 2000
rect 5445 1940 5515 1960
rect 5230 1925 5286 1931
rect 5230 1865 5234 1925
rect 5315 1915 5515 1940
rect 5570 1931 5600 2119
rect 5544 1925 5600 1931
rect 5286 1865 5544 1885
rect 5596 1865 5600 1925
rect 5230 1855 5600 1865
rect 5630 2185 6000 2195
rect 5630 2125 5634 2185
rect 5686 2165 5944 2185
rect 5630 2119 5686 2125
rect 5630 1931 5660 2119
rect 5715 2110 5915 2135
rect 5996 2125 6000 2185
rect 5944 2119 6000 2125
rect 5715 2090 5785 2110
rect 5690 2050 5785 2090
rect 5845 2090 5915 2110
rect 5845 2050 5940 2090
rect 5690 2000 5940 2050
rect 5690 1960 5785 2000
rect 5715 1940 5785 1960
rect 5845 1960 5940 2000
rect 5845 1940 5915 1960
rect 5630 1925 5686 1931
rect 5630 1865 5634 1925
rect 5715 1915 5915 1940
rect 5970 1931 6000 2119
rect 5944 1925 6000 1931
rect 5686 1865 5944 1885
rect 5996 1865 6000 1925
rect 5630 1855 6000 1865
rect 6030 2185 6400 2195
rect 6030 2125 6034 2185
rect 6086 2165 6344 2185
rect 6030 2119 6086 2125
rect 6030 1931 6060 2119
rect 6115 2110 6315 2135
rect 6396 2125 6400 2185
rect 6344 2119 6400 2125
rect 6115 2090 6185 2110
rect 6090 2050 6185 2090
rect 6245 2090 6315 2110
rect 6245 2050 6340 2090
rect 6090 2000 6340 2050
rect 6090 1960 6185 2000
rect 6115 1940 6185 1960
rect 6245 1960 6340 2000
rect 6245 1940 6315 1960
rect 6030 1925 6086 1931
rect 6030 1865 6034 1925
rect 6115 1915 6315 1940
rect 6370 1931 6400 2119
rect 6344 1925 6400 1931
rect 6086 1865 6344 1885
rect 6396 1865 6400 1925
rect 6030 1855 6400 1865
rect 6430 2185 6800 2195
rect 6430 2125 6434 2185
rect 6486 2165 6744 2185
rect 6430 2119 6486 2125
rect 6430 1931 6460 2119
rect 6515 2110 6715 2135
rect 6796 2125 6800 2185
rect 6744 2119 6800 2125
rect 6515 2090 6585 2110
rect 6490 2050 6585 2090
rect 6645 2090 6715 2110
rect 6645 2050 6740 2090
rect 6490 2000 6740 2050
rect 6490 1960 6585 2000
rect 6515 1940 6585 1960
rect 6645 1960 6740 2000
rect 6645 1940 6715 1960
rect 6430 1925 6486 1931
rect 6430 1865 6434 1925
rect 6515 1915 6715 1940
rect 6770 1931 6800 2119
rect 6744 1925 6800 1931
rect 6486 1865 6744 1885
rect 6796 1865 6800 1925
rect 6430 1855 6800 1865
rect 6830 2185 7200 2195
rect 6830 2125 6834 2185
rect 6886 2165 7144 2185
rect 6830 2119 6886 2125
rect 6830 1931 6860 2119
rect 6915 2110 7115 2135
rect 7196 2125 7200 2185
rect 7144 2119 7200 2125
rect 6915 2090 6985 2110
rect 6890 2050 6985 2090
rect 7045 2090 7115 2110
rect 7045 2050 7140 2090
rect 6890 2000 7140 2050
rect 6890 1960 6985 2000
rect 6915 1940 6985 1960
rect 7045 1960 7140 2000
rect 7045 1940 7115 1960
rect 6830 1925 6886 1931
rect 6830 1865 6834 1925
rect 6915 1915 7115 1940
rect 7170 1931 7200 2119
rect 7144 1925 7200 1931
rect 6886 1865 7144 1885
rect 7196 1865 7200 1925
rect 6830 1855 7200 1865
rect 7230 2185 7600 2195
rect 7230 2125 7234 2185
rect 7286 2165 7544 2185
rect 7230 2119 7286 2125
rect 7230 1931 7260 2119
rect 7315 2110 7515 2135
rect 7596 2125 7600 2185
rect 7544 2119 7600 2125
rect 7315 2090 7385 2110
rect 7290 2050 7385 2090
rect 7445 2090 7515 2110
rect 7445 2050 7540 2090
rect 7290 2000 7540 2050
rect 7290 1960 7385 2000
rect 7315 1940 7385 1960
rect 7445 1960 7540 2000
rect 7445 1940 7515 1960
rect 7230 1925 7286 1931
rect 7230 1865 7234 1925
rect 7315 1915 7515 1940
rect 7570 1931 7600 2119
rect 7544 1925 7600 1931
rect 7286 1865 7544 1885
rect 7596 1865 7600 1925
rect 7230 1855 7600 1865
rect 7630 2185 8000 2195
rect 7630 2125 7634 2185
rect 7686 2165 7944 2185
rect 7630 2119 7686 2125
rect 7630 1931 7660 2119
rect 7715 2110 7915 2135
rect 7996 2125 8000 2185
rect 7944 2119 8000 2125
rect 7715 2090 7785 2110
rect 7690 2050 7785 2090
rect 7845 2090 7915 2110
rect 7845 2050 7940 2090
rect 7690 2000 7940 2050
rect 7690 1960 7785 2000
rect 7715 1940 7785 1960
rect 7845 1960 7940 2000
rect 7845 1940 7915 1960
rect 7630 1925 7686 1931
rect 7630 1865 7634 1925
rect 7715 1915 7915 1940
rect 7970 1931 8000 2119
rect 7944 1925 8000 1931
rect 7686 1865 7944 1885
rect 7996 1865 8000 1925
rect 7630 1855 8000 1865
rect 8030 2185 8400 2195
rect 8030 2125 8034 2185
rect 8086 2165 8344 2185
rect 8030 2119 8086 2125
rect 8030 1931 8060 2119
rect 8115 2110 8315 2135
rect 8396 2125 8400 2185
rect 8344 2119 8400 2125
rect 8115 2090 8185 2110
rect 8090 2050 8185 2090
rect 8245 2090 8315 2110
rect 8245 2050 8340 2090
rect 8090 2000 8340 2050
rect 8090 1960 8185 2000
rect 8115 1940 8185 1960
rect 8245 1960 8340 2000
rect 8245 1940 8315 1960
rect 8030 1925 8086 1931
rect 8030 1865 8034 1925
rect 8115 1915 8315 1940
rect 8370 1931 8400 2119
rect 8344 1925 8400 1931
rect 8086 1865 8344 1885
rect 8396 1865 8400 1925
rect 8030 1855 8400 1865
rect 8430 2185 8800 2195
rect 8430 2125 8434 2185
rect 8486 2165 8744 2185
rect 8430 2119 8486 2125
rect 8430 1931 8460 2119
rect 8515 2110 8715 2135
rect 8796 2125 8800 2185
rect 8744 2119 8800 2125
rect 8515 2090 8585 2110
rect 8490 2050 8585 2090
rect 8645 2090 8715 2110
rect 8645 2050 8740 2090
rect 8490 2000 8740 2050
rect 8490 1960 8585 2000
rect 8515 1940 8585 1960
rect 8645 1960 8740 2000
rect 8645 1940 8715 1960
rect 8430 1925 8486 1931
rect 8430 1865 8434 1925
rect 8515 1915 8715 1940
rect 8770 1931 8800 2119
rect 8744 1925 8800 1931
rect 8486 1865 8744 1885
rect 8796 1865 8800 1925
rect 8430 1855 8800 1865
rect 8830 2185 9200 2195
rect 8830 2125 8834 2185
rect 8886 2165 9144 2185
rect 8830 2119 8886 2125
rect 8830 1931 8860 2119
rect 8915 2110 9115 2135
rect 9196 2125 9200 2185
rect 9144 2119 9200 2125
rect 8915 2090 8985 2110
rect 8890 2050 8985 2090
rect 9045 2090 9115 2110
rect 9045 2050 9140 2090
rect 8890 2000 9140 2050
rect 8890 1960 8985 2000
rect 8915 1940 8985 1960
rect 9045 1960 9140 2000
rect 9045 1940 9115 1960
rect 8830 1925 8886 1931
rect 8830 1865 8834 1925
rect 8915 1915 9115 1940
rect 9170 1931 9200 2119
rect 9144 1925 9200 1931
rect 8886 1865 9144 1885
rect 9196 1865 9200 1925
rect 8830 1855 9200 1865
rect 9230 2185 9600 2195
rect 9230 2125 9234 2185
rect 9286 2165 9544 2185
rect 9230 2119 9286 2125
rect 9230 1931 9260 2119
rect 9315 2110 9515 2135
rect 9596 2125 9600 2185
rect 9544 2119 9600 2125
rect 9315 2090 9385 2110
rect 9290 2050 9385 2090
rect 9445 2090 9515 2110
rect 9445 2050 9540 2090
rect 9290 2000 9540 2050
rect 9290 1960 9385 2000
rect 9315 1940 9385 1960
rect 9445 1960 9540 2000
rect 9445 1940 9515 1960
rect 9230 1925 9286 1931
rect 9230 1865 9234 1925
rect 9315 1915 9515 1940
rect 9570 1931 9600 2119
rect 9544 1925 9600 1931
rect 9286 1865 9544 1885
rect 9596 1865 9600 1925
rect 9230 1855 9600 1865
rect 9630 2185 10000 2195
rect 9630 2125 9634 2185
rect 9686 2165 9944 2185
rect 9630 2119 9686 2125
rect 9630 1931 9660 2119
rect 9715 2110 9915 2135
rect 9996 2125 10000 2185
rect 9944 2119 10000 2125
rect 9715 2090 9785 2110
rect 9690 2050 9785 2090
rect 9845 2090 9915 2110
rect 9845 2050 9940 2090
rect 9690 2000 9940 2050
rect 9690 1960 9785 2000
rect 9715 1940 9785 1960
rect 9845 1960 9940 2000
rect 9845 1940 9915 1960
rect 9630 1925 9686 1931
rect 9630 1865 9634 1925
rect 9715 1915 9915 1940
rect 9970 1931 10000 2119
rect 9944 1925 10000 1931
rect 9686 1865 9944 1885
rect 9996 1865 10000 1925
rect 9630 1855 10000 1865
rect 10030 2185 10400 2195
rect 10030 2125 10034 2185
rect 10086 2165 10344 2185
rect 10030 2119 10086 2125
rect 10030 1931 10060 2119
rect 10115 2110 10315 2135
rect 10396 2125 10400 2185
rect 10344 2119 10400 2125
rect 10115 2090 10185 2110
rect 10090 2050 10185 2090
rect 10245 2090 10315 2110
rect 10245 2050 10340 2090
rect 10090 2000 10340 2050
rect 10090 1960 10185 2000
rect 10115 1940 10185 1960
rect 10245 1960 10340 2000
rect 10245 1940 10315 1960
rect 10030 1925 10086 1931
rect 10030 1865 10034 1925
rect 10115 1915 10315 1940
rect 10370 1931 10400 2119
rect 10344 1925 10400 1931
rect 10086 1865 10344 1885
rect 10396 1865 10400 1925
rect 10030 1855 10400 1865
rect 10430 2185 10800 2195
rect 10430 2125 10434 2185
rect 10486 2165 10744 2185
rect 10430 2119 10486 2125
rect 10430 1931 10460 2119
rect 10515 2110 10715 2135
rect 10796 2125 10800 2185
rect 10744 2119 10800 2125
rect 10515 2090 10585 2110
rect 10490 2050 10585 2090
rect 10645 2090 10715 2110
rect 10645 2050 10740 2090
rect 10490 2000 10740 2050
rect 10490 1960 10585 2000
rect 10515 1940 10585 1960
rect 10645 1960 10740 2000
rect 10645 1940 10715 1960
rect 10430 1925 10486 1931
rect 10430 1865 10434 1925
rect 10515 1915 10715 1940
rect 10770 1931 10800 2119
rect 10744 1925 10800 1931
rect 10486 1865 10744 1885
rect 10796 1865 10800 1925
rect 10430 1855 10800 1865
rect 10830 2185 11200 2195
rect 10830 2125 10834 2185
rect 10886 2165 11144 2185
rect 10830 2119 10886 2125
rect 10830 1931 10860 2119
rect 10915 2110 11115 2135
rect 11196 2125 11200 2185
rect 11144 2119 11200 2125
rect 10915 2090 10985 2110
rect 10890 2050 10985 2090
rect 11045 2090 11115 2110
rect 11045 2050 11140 2090
rect 10890 2000 11140 2050
rect 10890 1960 10985 2000
rect 10915 1940 10985 1960
rect 11045 1960 11140 2000
rect 11045 1940 11115 1960
rect 10830 1925 10886 1931
rect 10830 1865 10834 1925
rect 10915 1915 11115 1940
rect 11170 1931 11200 2119
rect 11144 1925 11200 1931
rect 10886 1865 11144 1885
rect 11196 1865 11200 1925
rect 10830 1855 11200 1865
rect 11230 2185 11600 2195
rect 11230 2125 11234 2185
rect 11286 2165 11544 2185
rect 11230 2119 11286 2125
rect 11230 1931 11260 2119
rect 11315 2110 11515 2135
rect 11596 2125 11600 2185
rect 11544 2119 11600 2125
rect 11315 2090 11385 2110
rect 11290 2050 11385 2090
rect 11445 2090 11515 2110
rect 11445 2050 11540 2090
rect 11290 2000 11540 2050
rect 11290 1960 11385 2000
rect 11315 1940 11385 1960
rect 11445 1960 11540 2000
rect 11445 1940 11515 1960
rect 11230 1925 11286 1931
rect 11230 1865 11234 1925
rect 11315 1915 11515 1940
rect 11570 1931 11600 2119
rect 11544 1925 11600 1931
rect 11286 1865 11544 1885
rect 11596 1865 11600 1925
rect 11230 1855 11600 1865
rect 11630 2185 12000 2195
rect 11630 2125 11634 2185
rect 11686 2165 11944 2185
rect 11630 2119 11686 2125
rect 11630 1931 11660 2119
rect 11715 2110 11915 2135
rect 11996 2125 12000 2185
rect 11944 2119 12000 2125
rect 11715 2090 11785 2110
rect 11690 2050 11785 2090
rect 11845 2090 11915 2110
rect 11845 2050 11940 2090
rect 11690 2000 11940 2050
rect 11690 1960 11785 2000
rect 11715 1940 11785 1960
rect 11845 1960 11940 2000
rect 11845 1940 11915 1960
rect 11630 1925 11686 1931
rect 11630 1865 11634 1925
rect 11715 1915 11915 1940
rect 11970 1931 12000 2119
rect 11944 1925 12000 1931
rect 11686 1865 11944 1885
rect 11996 1865 12000 1925
rect 11630 1855 12000 1865
rect 12030 2185 12400 2195
rect 12030 2125 12034 2185
rect 12086 2165 12344 2185
rect 12030 2119 12086 2125
rect 12030 1931 12060 2119
rect 12115 2110 12315 2135
rect 12396 2125 12400 2185
rect 12344 2119 12400 2125
rect 12115 2090 12185 2110
rect 12090 2050 12185 2090
rect 12245 2090 12315 2110
rect 12245 2050 12340 2090
rect 12090 2000 12340 2050
rect 12090 1960 12185 2000
rect 12115 1940 12185 1960
rect 12245 1960 12340 2000
rect 12245 1940 12315 1960
rect 12030 1925 12086 1931
rect 12030 1865 12034 1925
rect 12115 1915 12315 1940
rect 12370 1931 12400 2119
rect 12344 1925 12400 1931
rect 12086 1865 12344 1885
rect 12396 1865 12400 1925
rect 12030 1855 12400 1865
rect 12430 2185 12800 2195
rect 12430 2125 12434 2185
rect 12486 2165 12744 2185
rect 12430 2119 12486 2125
rect 12430 1931 12460 2119
rect 12515 2110 12715 2135
rect 12796 2125 12800 2185
rect 12744 2119 12800 2125
rect 12515 2090 12585 2110
rect 12490 2050 12585 2090
rect 12645 2090 12715 2110
rect 12645 2050 12740 2090
rect 12490 2000 12740 2050
rect 12490 1960 12585 2000
rect 12515 1940 12585 1960
rect 12645 1960 12740 2000
rect 12645 1940 12715 1960
rect 12430 1925 12486 1931
rect 12430 1865 12434 1925
rect 12515 1915 12715 1940
rect 12770 1931 12800 2119
rect 12744 1925 12800 1931
rect 12486 1865 12744 1885
rect 12796 1865 12800 1925
rect 12430 1855 12800 1865
rect 12830 2185 13200 2195
rect 12830 2125 12834 2185
rect 12886 2165 13144 2185
rect 12830 2119 12886 2125
rect 12830 1931 12860 2119
rect 12915 2110 13115 2135
rect 13196 2125 13200 2185
rect 13144 2119 13200 2125
rect 12915 2090 12985 2110
rect 12890 2050 12985 2090
rect 13045 2090 13115 2110
rect 13045 2050 13140 2090
rect 12890 2000 13140 2050
rect 12890 1960 12985 2000
rect 12915 1940 12985 1960
rect 13045 1960 13140 2000
rect 13045 1940 13115 1960
rect 12830 1925 12886 1931
rect 12830 1865 12834 1925
rect 12915 1915 13115 1940
rect 13170 1931 13200 2119
rect 13144 1925 13200 1931
rect 12886 1865 13144 1885
rect 13196 1865 13200 1925
rect 12830 1855 13200 1865
rect -370 1815 0 1825
rect -370 1755 -366 1815
rect -314 1795 -56 1815
rect -370 1749 -314 1755
rect -370 1561 -340 1749
rect -285 1740 -85 1765
rect -4 1755 0 1815
rect -56 1749 0 1755
rect -285 1720 -215 1740
rect -310 1680 -215 1720
rect -155 1720 -85 1740
rect -155 1680 -60 1720
rect -310 1630 -60 1680
rect -310 1590 -215 1630
rect -285 1570 -215 1590
rect -155 1590 -60 1630
rect -155 1570 -85 1590
rect -370 1555 -314 1561
rect -370 1495 -366 1555
rect -285 1545 -85 1570
rect -30 1561 0 1749
rect -56 1555 0 1561
rect -314 1495 -56 1515
rect -4 1495 0 1555
rect -370 1485 0 1495
rect 30 1815 400 1825
rect 30 1755 34 1815
rect 86 1795 344 1815
rect 30 1749 86 1755
rect 30 1561 60 1749
rect 115 1740 315 1765
rect 396 1755 400 1815
rect 344 1749 400 1755
rect 115 1720 185 1740
rect 90 1680 185 1720
rect 245 1720 315 1740
rect 245 1680 340 1720
rect 90 1630 340 1680
rect 90 1590 185 1630
rect 115 1570 185 1590
rect 245 1590 340 1630
rect 245 1570 315 1590
rect 30 1555 86 1561
rect 30 1495 34 1555
rect 115 1545 315 1570
rect 370 1561 400 1749
rect 344 1555 400 1561
rect 86 1495 344 1515
rect 396 1495 400 1555
rect 30 1485 400 1495
rect 430 1815 800 1825
rect 430 1755 434 1815
rect 486 1795 744 1815
rect 430 1749 486 1755
rect 430 1561 460 1749
rect 515 1740 715 1765
rect 796 1755 800 1815
rect 744 1749 800 1755
rect 515 1720 585 1740
rect 490 1680 585 1720
rect 645 1720 715 1740
rect 645 1680 740 1720
rect 490 1630 740 1680
rect 490 1590 585 1630
rect 515 1570 585 1590
rect 645 1590 740 1630
rect 645 1570 715 1590
rect 430 1555 486 1561
rect 430 1495 434 1555
rect 515 1545 715 1570
rect 770 1561 800 1749
rect 744 1555 800 1561
rect 486 1495 744 1515
rect 796 1495 800 1555
rect 430 1485 800 1495
rect 830 1815 1200 1825
rect 830 1755 834 1815
rect 886 1795 1144 1815
rect 830 1749 886 1755
rect 830 1561 860 1749
rect 915 1740 1115 1765
rect 1196 1755 1200 1815
rect 1144 1749 1200 1755
rect 915 1720 985 1740
rect 890 1680 985 1720
rect 1045 1720 1115 1740
rect 1045 1680 1140 1720
rect 890 1630 1140 1680
rect 890 1590 985 1630
rect 915 1570 985 1590
rect 1045 1590 1140 1630
rect 1045 1570 1115 1590
rect 830 1555 886 1561
rect 830 1495 834 1555
rect 915 1545 1115 1570
rect 1170 1561 1200 1749
rect 1144 1555 1200 1561
rect 886 1495 1144 1515
rect 1196 1495 1200 1555
rect 830 1485 1200 1495
rect 1230 1815 1600 1825
rect 1230 1755 1234 1815
rect 1286 1795 1544 1815
rect 1230 1749 1286 1755
rect 1230 1561 1260 1749
rect 1315 1740 1515 1765
rect 1596 1755 1600 1815
rect 1544 1749 1600 1755
rect 1315 1720 1385 1740
rect 1290 1680 1385 1720
rect 1445 1720 1515 1740
rect 1445 1680 1540 1720
rect 1290 1630 1540 1680
rect 1290 1590 1385 1630
rect 1315 1570 1385 1590
rect 1445 1590 1540 1630
rect 1445 1570 1515 1590
rect 1230 1555 1286 1561
rect 1230 1495 1234 1555
rect 1315 1545 1515 1570
rect 1570 1561 1600 1749
rect 1544 1555 1600 1561
rect 1286 1495 1544 1515
rect 1596 1495 1600 1555
rect 1230 1485 1600 1495
rect 1630 1815 2000 1825
rect 1630 1755 1634 1815
rect 1686 1795 1944 1815
rect 1630 1749 1686 1755
rect 1630 1561 1660 1749
rect 1715 1740 1915 1765
rect 1996 1755 2000 1815
rect 1944 1749 2000 1755
rect 1715 1720 1785 1740
rect 1690 1680 1785 1720
rect 1845 1720 1915 1740
rect 1845 1680 1940 1720
rect 1690 1630 1940 1680
rect 1690 1590 1785 1630
rect 1715 1570 1785 1590
rect 1845 1590 1940 1630
rect 1845 1570 1915 1590
rect 1630 1555 1686 1561
rect 1630 1495 1634 1555
rect 1715 1545 1915 1570
rect 1970 1561 2000 1749
rect 1944 1555 2000 1561
rect 1686 1495 1944 1515
rect 1996 1495 2000 1555
rect 1630 1485 2000 1495
rect 2030 1815 2400 1825
rect 2030 1755 2034 1815
rect 2086 1795 2344 1815
rect 2030 1749 2086 1755
rect 2030 1561 2060 1749
rect 2115 1740 2315 1765
rect 2396 1755 2400 1815
rect 2344 1749 2400 1755
rect 2115 1720 2185 1740
rect 2090 1680 2185 1720
rect 2245 1720 2315 1740
rect 2245 1680 2340 1720
rect 2090 1630 2340 1680
rect 2090 1590 2185 1630
rect 2115 1570 2185 1590
rect 2245 1590 2340 1630
rect 2245 1570 2315 1590
rect 2030 1555 2086 1561
rect 2030 1495 2034 1555
rect 2115 1545 2315 1570
rect 2370 1561 2400 1749
rect 2344 1555 2400 1561
rect 2086 1495 2344 1515
rect 2396 1495 2400 1555
rect 2030 1485 2400 1495
rect 2430 1815 2800 1825
rect 2430 1755 2434 1815
rect 2486 1795 2744 1815
rect 2430 1749 2486 1755
rect 2430 1561 2460 1749
rect 2515 1740 2715 1765
rect 2796 1755 2800 1815
rect 2744 1749 2800 1755
rect 2515 1720 2585 1740
rect 2490 1680 2585 1720
rect 2645 1720 2715 1740
rect 2645 1680 2740 1720
rect 2490 1630 2740 1680
rect 2490 1590 2585 1630
rect 2515 1570 2585 1590
rect 2645 1590 2740 1630
rect 2645 1570 2715 1590
rect 2430 1555 2486 1561
rect 2430 1495 2434 1555
rect 2515 1545 2715 1570
rect 2770 1561 2800 1749
rect 2744 1555 2800 1561
rect 2486 1495 2744 1515
rect 2796 1495 2800 1555
rect 2430 1485 2800 1495
rect 2830 1815 3200 1825
rect 2830 1755 2834 1815
rect 2886 1795 3144 1815
rect 2830 1749 2886 1755
rect 2830 1561 2860 1749
rect 2915 1740 3115 1765
rect 3196 1755 3200 1815
rect 3144 1749 3200 1755
rect 2915 1720 2985 1740
rect 2890 1680 2985 1720
rect 3045 1720 3115 1740
rect 3045 1680 3140 1720
rect 2890 1630 3140 1680
rect 2890 1590 2985 1630
rect 2915 1570 2985 1590
rect 3045 1590 3140 1630
rect 3045 1570 3115 1590
rect 2830 1555 2886 1561
rect 2830 1495 2834 1555
rect 2915 1545 3115 1570
rect 3170 1561 3200 1749
rect 3144 1555 3200 1561
rect 2886 1495 3144 1515
rect 3196 1495 3200 1555
rect 2830 1485 3200 1495
rect 3230 1815 3600 1825
rect 3230 1755 3234 1815
rect 3286 1795 3544 1815
rect 3230 1749 3286 1755
rect 3230 1561 3260 1749
rect 3315 1740 3515 1765
rect 3596 1755 3600 1815
rect 3544 1749 3600 1755
rect 3315 1720 3385 1740
rect 3290 1680 3385 1720
rect 3445 1720 3515 1740
rect 3445 1680 3540 1720
rect 3290 1630 3540 1680
rect 3290 1590 3385 1630
rect 3315 1570 3385 1590
rect 3445 1590 3540 1630
rect 3445 1570 3515 1590
rect 3230 1555 3286 1561
rect 3230 1495 3234 1555
rect 3315 1545 3515 1570
rect 3570 1561 3600 1749
rect 3544 1555 3600 1561
rect 3286 1495 3544 1515
rect 3596 1495 3600 1555
rect 3230 1485 3600 1495
rect 3630 1815 4000 1825
rect 3630 1755 3634 1815
rect 3686 1795 3944 1815
rect 3630 1749 3686 1755
rect 3630 1561 3660 1749
rect 3715 1740 3915 1765
rect 3996 1755 4000 1815
rect 3944 1749 4000 1755
rect 3715 1720 3785 1740
rect 3690 1680 3785 1720
rect 3845 1720 3915 1740
rect 3845 1680 3940 1720
rect 3690 1630 3940 1680
rect 3690 1590 3785 1630
rect 3715 1570 3785 1590
rect 3845 1590 3940 1630
rect 3845 1570 3915 1590
rect 3630 1555 3686 1561
rect 3630 1495 3634 1555
rect 3715 1545 3915 1570
rect 3970 1561 4000 1749
rect 3944 1555 4000 1561
rect 3686 1495 3944 1515
rect 3996 1495 4000 1555
rect 3630 1485 4000 1495
rect 4030 1815 4400 1825
rect 4030 1755 4034 1815
rect 4086 1795 4344 1815
rect 4030 1749 4086 1755
rect 4030 1561 4060 1749
rect 4115 1740 4315 1765
rect 4396 1755 4400 1815
rect 4344 1749 4400 1755
rect 4115 1720 4185 1740
rect 4090 1680 4185 1720
rect 4245 1720 4315 1740
rect 4245 1680 4340 1720
rect 4090 1630 4340 1680
rect 4090 1590 4185 1630
rect 4115 1570 4185 1590
rect 4245 1590 4340 1630
rect 4245 1570 4315 1590
rect 4030 1555 4086 1561
rect 4030 1495 4034 1555
rect 4115 1545 4315 1570
rect 4370 1561 4400 1749
rect 4344 1555 4400 1561
rect 4086 1495 4344 1515
rect 4396 1495 4400 1555
rect 4030 1485 4400 1495
rect 4430 1815 4800 1825
rect 4430 1755 4434 1815
rect 4486 1795 4744 1815
rect 4430 1749 4486 1755
rect 4430 1561 4460 1749
rect 4515 1740 4715 1765
rect 4796 1755 4800 1815
rect 4744 1749 4800 1755
rect 4515 1720 4585 1740
rect 4490 1680 4585 1720
rect 4645 1720 4715 1740
rect 4645 1680 4740 1720
rect 4490 1630 4740 1680
rect 4490 1590 4585 1630
rect 4515 1570 4585 1590
rect 4645 1590 4740 1630
rect 4645 1570 4715 1590
rect 4430 1555 4486 1561
rect 4430 1495 4434 1555
rect 4515 1545 4715 1570
rect 4770 1561 4800 1749
rect 4744 1555 4800 1561
rect 4486 1495 4744 1515
rect 4796 1495 4800 1555
rect 4430 1485 4800 1495
rect 4830 1815 5200 1825
rect 4830 1755 4834 1815
rect 4886 1795 5144 1815
rect 4830 1749 4886 1755
rect 4830 1561 4860 1749
rect 4915 1740 5115 1765
rect 5196 1755 5200 1815
rect 5144 1749 5200 1755
rect 4915 1720 4985 1740
rect 4890 1680 4985 1720
rect 5045 1720 5115 1740
rect 5045 1680 5140 1720
rect 4890 1630 5140 1680
rect 4890 1590 4985 1630
rect 4915 1570 4985 1590
rect 5045 1590 5140 1630
rect 5045 1570 5115 1590
rect 4830 1555 4886 1561
rect 4830 1495 4834 1555
rect 4915 1545 5115 1570
rect 5170 1561 5200 1749
rect 5144 1555 5200 1561
rect 4886 1495 5144 1515
rect 5196 1495 5200 1555
rect 4830 1485 5200 1495
rect 5230 1815 5600 1825
rect 5230 1755 5234 1815
rect 5286 1795 5544 1815
rect 5230 1749 5286 1755
rect 5230 1561 5260 1749
rect 5315 1740 5515 1765
rect 5596 1755 5600 1815
rect 5544 1749 5600 1755
rect 5315 1720 5385 1740
rect 5290 1680 5385 1720
rect 5445 1720 5515 1740
rect 5445 1680 5540 1720
rect 5290 1630 5540 1680
rect 5290 1590 5385 1630
rect 5315 1570 5385 1590
rect 5445 1590 5540 1630
rect 5445 1570 5515 1590
rect 5230 1555 5286 1561
rect 5230 1495 5234 1555
rect 5315 1545 5515 1570
rect 5570 1561 5600 1749
rect 5544 1555 5600 1561
rect 5286 1495 5544 1515
rect 5596 1495 5600 1555
rect 5230 1485 5600 1495
rect 5630 1815 6000 1825
rect 5630 1755 5634 1815
rect 5686 1795 5944 1815
rect 5630 1749 5686 1755
rect 5630 1561 5660 1749
rect 5715 1740 5915 1765
rect 5996 1755 6000 1815
rect 5944 1749 6000 1755
rect 5715 1720 5785 1740
rect 5690 1680 5785 1720
rect 5845 1720 5915 1740
rect 5845 1680 5940 1720
rect 5690 1630 5940 1680
rect 5690 1590 5785 1630
rect 5715 1570 5785 1590
rect 5845 1590 5940 1630
rect 5845 1570 5915 1590
rect 5630 1555 5686 1561
rect 5630 1495 5634 1555
rect 5715 1545 5915 1570
rect 5970 1561 6000 1749
rect 5944 1555 6000 1561
rect 5686 1495 5944 1515
rect 5996 1495 6000 1555
rect 5630 1485 6000 1495
rect 6030 1815 6400 1825
rect 6030 1755 6034 1815
rect 6086 1795 6344 1815
rect 6030 1749 6086 1755
rect 6030 1561 6060 1749
rect 6115 1740 6315 1765
rect 6396 1755 6400 1815
rect 6344 1749 6400 1755
rect 6115 1720 6185 1740
rect 6090 1680 6185 1720
rect 6245 1720 6315 1740
rect 6245 1680 6340 1720
rect 6090 1630 6340 1680
rect 6090 1590 6185 1630
rect 6115 1570 6185 1590
rect 6245 1590 6340 1630
rect 6245 1570 6315 1590
rect 6030 1555 6086 1561
rect 6030 1495 6034 1555
rect 6115 1545 6315 1570
rect 6370 1561 6400 1749
rect 6344 1555 6400 1561
rect 6086 1495 6344 1515
rect 6396 1495 6400 1555
rect 6030 1485 6400 1495
rect 6430 1815 6800 1825
rect 6430 1755 6434 1815
rect 6486 1795 6744 1815
rect 6430 1749 6486 1755
rect 6430 1561 6460 1749
rect 6515 1740 6715 1765
rect 6796 1755 6800 1815
rect 6744 1749 6800 1755
rect 6515 1720 6585 1740
rect 6490 1680 6585 1720
rect 6645 1720 6715 1740
rect 6645 1680 6740 1720
rect 6490 1630 6740 1680
rect 6490 1590 6585 1630
rect 6515 1570 6585 1590
rect 6645 1590 6740 1630
rect 6645 1570 6715 1590
rect 6430 1555 6486 1561
rect 6430 1495 6434 1555
rect 6515 1545 6715 1570
rect 6770 1561 6800 1749
rect 6744 1555 6800 1561
rect 6486 1495 6744 1515
rect 6796 1495 6800 1555
rect 6430 1485 6800 1495
rect 6830 1815 7200 1825
rect 6830 1755 6834 1815
rect 6886 1795 7144 1815
rect 6830 1749 6886 1755
rect 6830 1561 6860 1749
rect 6915 1740 7115 1765
rect 7196 1755 7200 1815
rect 7144 1749 7200 1755
rect 6915 1720 6985 1740
rect 6890 1680 6985 1720
rect 7045 1720 7115 1740
rect 7045 1680 7140 1720
rect 6890 1630 7140 1680
rect 6890 1590 6985 1630
rect 6915 1570 6985 1590
rect 7045 1590 7140 1630
rect 7045 1570 7115 1590
rect 6830 1555 6886 1561
rect 6830 1495 6834 1555
rect 6915 1545 7115 1570
rect 7170 1561 7200 1749
rect 7144 1555 7200 1561
rect 6886 1495 7144 1515
rect 7196 1495 7200 1555
rect 6830 1485 7200 1495
rect 7230 1815 7600 1825
rect 7230 1755 7234 1815
rect 7286 1795 7544 1815
rect 7230 1749 7286 1755
rect 7230 1561 7260 1749
rect 7315 1740 7515 1765
rect 7596 1755 7600 1815
rect 7544 1749 7600 1755
rect 7315 1720 7385 1740
rect 7290 1680 7385 1720
rect 7445 1720 7515 1740
rect 7445 1680 7540 1720
rect 7290 1630 7540 1680
rect 7290 1590 7385 1630
rect 7315 1570 7385 1590
rect 7445 1590 7540 1630
rect 7445 1570 7515 1590
rect 7230 1555 7286 1561
rect 7230 1495 7234 1555
rect 7315 1545 7515 1570
rect 7570 1561 7600 1749
rect 7544 1555 7600 1561
rect 7286 1495 7544 1515
rect 7596 1495 7600 1555
rect 7230 1485 7600 1495
rect 7630 1815 8000 1825
rect 7630 1755 7634 1815
rect 7686 1795 7944 1815
rect 7630 1749 7686 1755
rect 7630 1561 7660 1749
rect 7715 1740 7915 1765
rect 7996 1755 8000 1815
rect 7944 1749 8000 1755
rect 7715 1720 7785 1740
rect 7690 1680 7785 1720
rect 7845 1720 7915 1740
rect 7845 1680 7940 1720
rect 7690 1630 7940 1680
rect 7690 1590 7785 1630
rect 7715 1570 7785 1590
rect 7845 1590 7940 1630
rect 7845 1570 7915 1590
rect 7630 1555 7686 1561
rect 7630 1495 7634 1555
rect 7715 1545 7915 1570
rect 7970 1561 8000 1749
rect 7944 1555 8000 1561
rect 7686 1495 7944 1515
rect 7996 1495 8000 1555
rect 7630 1485 8000 1495
rect 8030 1815 8400 1825
rect 8030 1755 8034 1815
rect 8086 1795 8344 1815
rect 8030 1749 8086 1755
rect 8030 1561 8060 1749
rect 8115 1740 8315 1765
rect 8396 1755 8400 1815
rect 8344 1749 8400 1755
rect 8115 1720 8185 1740
rect 8090 1680 8185 1720
rect 8245 1720 8315 1740
rect 8245 1680 8340 1720
rect 8090 1630 8340 1680
rect 8090 1590 8185 1630
rect 8115 1570 8185 1590
rect 8245 1590 8340 1630
rect 8245 1570 8315 1590
rect 8030 1555 8086 1561
rect 8030 1495 8034 1555
rect 8115 1545 8315 1570
rect 8370 1561 8400 1749
rect 8344 1555 8400 1561
rect 8086 1495 8344 1515
rect 8396 1495 8400 1555
rect 8030 1485 8400 1495
rect 8430 1815 8800 1825
rect 8430 1755 8434 1815
rect 8486 1795 8744 1815
rect 8430 1749 8486 1755
rect 8430 1561 8460 1749
rect 8515 1740 8715 1765
rect 8796 1755 8800 1815
rect 8744 1749 8800 1755
rect 8515 1720 8585 1740
rect 8490 1680 8585 1720
rect 8645 1720 8715 1740
rect 8645 1680 8740 1720
rect 8490 1630 8740 1680
rect 8490 1590 8585 1630
rect 8515 1570 8585 1590
rect 8645 1590 8740 1630
rect 8645 1570 8715 1590
rect 8430 1555 8486 1561
rect 8430 1495 8434 1555
rect 8515 1545 8715 1570
rect 8770 1561 8800 1749
rect 8744 1555 8800 1561
rect 8486 1495 8744 1515
rect 8796 1495 8800 1555
rect 8430 1485 8800 1495
rect 8830 1815 9200 1825
rect 8830 1755 8834 1815
rect 8886 1795 9144 1815
rect 8830 1749 8886 1755
rect 8830 1561 8860 1749
rect 8915 1740 9115 1765
rect 9196 1755 9200 1815
rect 9144 1749 9200 1755
rect 8915 1720 8985 1740
rect 8890 1680 8985 1720
rect 9045 1720 9115 1740
rect 9045 1680 9140 1720
rect 8890 1630 9140 1680
rect 8890 1590 8985 1630
rect 8915 1570 8985 1590
rect 9045 1590 9140 1630
rect 9045 1570 9115 1590
rect 8830 1555 8886 1561
rect 8830 1495 8834 1555
rect 8915 1545 9115 1570
rect 9170 1561 9200 1749
rect 9144 1555 9200 1561
rect 8886 1495 9144 1515
rect 9196 1495 9200 1555
rect 8830 1485 9200 1495
rect 9230 1815 9600 1825
rect 9230 1755 9234 1815
rect 9286 1795 9544 1815
rect 9230 1749 9286 1755
rect 9230 1561 9260 1749
rect 9315 1740 9515 1765
rect 9596 1755 9600 1815
rect 9544 1749 9600 1755
rect 9315 1720 9385 1740
rect 9290 1680 9385 1720
rect 9445 1720 9515 1740
rect 9445 1680 9540 1720
rect 9290 1630 9540 1680
rect 9290 1590 9385 1630
rect 9315 1570 9385 1590
rect 9445 1590 9540 1630
rect 9445 1570 9515 1590
rect 9230 1555 9286 1561
rect 9230 1495 9234 1555
rect 9315 1545 9515 1570
rect 9570 1561 9600 1749
rect 9544 1555 9600 1561
rect 9286 1495 9544 1515
rect 9596 1495 9600 1555
rect 9230 1485 9600 1495
rect 9630 1815 10000 1825
rect 9630 1755 9634 1815
rect 9686 1795 9944 1815
rect 9630 1749 9686 1755
rect 9630 1561 9660 1749
rect 9715 1740 9915 1765
rect 9996 1755 10000 1815
rect 9944 1749 10000 1755
rect 9715 1720 9785 1740
rect 9690 1680 9785 1720
rect 9845 1720 9915 1740
rect 9845 1680 9940 1720
rect 9690 1630 9940 1680
rect 9690 1590 9785 1630
rect 9715 1570 9785 1590
rect 9845 1590 9940 1630
rect 9845 1570 9915 1590
rect 9630 1555 9686 1561
rect 9630 1495 9634 1555
rect 9715 1545 9915 1570
rect 9970 1561 10000 1749
rect 9944 1555 10000 1561
rect 9686 1495 9944 1515
rect 9996 1495 10000 1555
rect 9630 1485 10000 1495
rect 10030 1815 10400 1825
rect 10030 1755 10034 1815
rect 10086 1795 10344 1815
rect 10030 1749 10086 1755
rect 10030 1561 10060 1749
rect 10115 1740 10315 1765
rect 10396 1755 10400 1815
rect 10344 1749 10400 1755
rect 10115 1720 10185 1740
rect 10090 1680 10185 1720
rect 10245 1720 10315 1740
rect 10245 1680 10340 1720
rect 10090 1630 10340 1680
rect 10090 1590 10185 1630
rect 10115 1570 10185 1590
rect 10245 1590 10340 1630
rect 10245 1570 10315 1590
rect 10030 1555 10086 1561
rect 10030 1495 10034 1555
rect 10115 1545 10315 1570
rect 10370 1561 10400 1749
rect 10344 1555 10400 1561
rect 10086 1495 10344 1515
rect 10396 1495 10400 1555
rect 10030 1485 10400 1495
rect 10430 1815 10800 1825
rect 10430 1755 10434 1815
rect 10486 1795 10744 1815
rect 10430 1749 10486 1755
rect 10430 1561 10460 1749
rect 10515 1740 10715 1765
rect 10796 1755 10800 1815
rect 10744 1749 10800 1755
rect 10515 1720 10585 1740
rect 10490 1680 10585 1720
rect 10645 1720 10715 1740
rect 10645 1680 10740 1720
rect 10490 1630 10740 1680
rect 10490 1590 10585 1630
rect 10515 1570 10585 1590
rect 10645 1590 10740 1630
rect 10645 1570 10715 1590
rect 10430 1555 10486 1561
rect 10430 1495 10434 1555
rect 10515 1545 10715 1570
rect 10770 1561 10800 1749
rect 10744 1555 10800 1561
rect 10486 1495 10744 1515
rect 10796 1495 10800 1555
rect 10430 1485 10800 1495
rect 10830 1815 11200 1825
rect 10830 1755 10834 1815
rect 10886 1795 11144 1815
rect 10830 1749 10886 1755
rect 10830 1561 10860 1749
rect 10915 1740 11115 1765
rect 11196 1755 11200 1815
rect 11144 1749 11200 1755
rect 10915 1720 10985 1740
rect 10890 1680 10985 1720
rect 11045 1720 11115 1740
rect 11045 1680 11140 1720
rect 10890 1630 11140 1680
rect 10890 1590 10985 1630
rect 10915 1570 10985 1590
rect 11045 1590 11140 1630
rect 11045 1570 11115 1590
rect 10830 1555 10886 1561
rect 10830 1495 10834 1555
rect 10915 1545 11115 1570
rect 11170 1561 11200 1749
rect 11144 1555 11200 1561
rect 10886 1495 11144 1515
rect 11196 1495 11200 1555
rect 10830 1485 11200 1495
rect 11230 1815 11600 1825
rect 11230 1755 11234 1815
rect 11286 1795 11544 1815
rect 11230 1749 11286 1755
rect 11230 1561 11260 1749
rect 11315 1740 11515 1765
rect 11596 1755 11600 1815
rect 11544 1749 11600 1755
rect 11315 1720 11385 1740
rect 11290 1680 11385 1720
rect 11445 1720 11515 1740
rect 11445 1680 11540 1720
rect 11290 1630 11540 1680
rect 11290 1590 11385 1630
rect 11315 1570 11385 1590
rect 11445 1590 11540 1630
rect 11445 1570 11515 1590
rect 11230 1555 11286 1561
rect 11230 1495 11234 1555
rect 11315 1545 11515 1570
rect 11570 1561 11600 1749
rect 11544 1555 11600 1561
rect 11286 1495 11544 1515
rect 11596 1495 11600 1555
rect 11230 1485 11600 1495
rect 11630 1815 12000 1825
rect 11630 1755 11634 1815
rect 11686 1795 11944 1815
rect 11630 1749 11686 1755
rect 11630 1561 11660 1749
rect 11715 1740 11915 1765
rect 11996 1755 12000 1815
rect 11944 1749 12000 1755
rect 11715 1720 11785 1740
rect 11690 1680 11785 1720
rect 11845 1720 11915 1740
rect 11845 1680 11940 1720
rect 11690 1630 11940 1680
rect 11690 1590 11785 1630
rect 11715 1570 11785 1590
rect 11845 1590 11940 1630
rect 11845 1570 11915 1590
rect 11630 1555 11686 1561
rect 11630 1495 11634 1555
rect 11715 1545 11915 1570
rect 11970 1561 12000 1749
rect 11944 1555 12000 1561
rect 11686 1495 11944 1515
rect 11996 1495 12000 1555
rect 11630 1485 12000 1495
rect 12030 1815 12400 1825
rect 12030 1755 12034 1815
rect 12086 1795 12344 1815
rect 12030 1749 12086 1755
rect 12030 1561 12060 1749
rect 12115 1740 12315 1765
rect 12396 1755 12400 1815
rect 12344 1749 12400 1755
rect 12115 1720 12185 1740
rect 12090 1680 12185 1720
rect 12245 1720 12315 1740
rect 12245 1680 12340 1720
rect 12090 1630 12340 1680
rect 12090 1590 12185 1630
rect 12115 1570 12185 1590
rect 12245 1590 12340 1630
rect 12245 1570 12315 1590
rect 12030 1555 12086 1561
rect 12030 1495 12034 1555
rect 12115 1545 12315 1570
rect 12370 1561 12400 1749
rect 12344 1555 12400 1561
rect 12086 1495 12344 1515
rect 12396 1495 12400 1555
rect 12030 1485 12400 1495
rect 12430 1815 12800 1825
rect 12430 1755 12434 1815
rect 12486 1795 12744 1815
rect 12430 1749 12486 1755
rect 12430 1561 12460 1749
rect 12515 1740 12715 1765
rect 12796 1755 12800 1815
rect 12744 1749 12800 1755
rect 12515 1720 12585 1740
rect 12490 1680 12585 1720
rect 12645 1720 12715 1740
rect 12645 1680 12740 1720
rect 12490 1630 12740 1680
rect 12490 1590 12585 1630
rect 12515 1570 12585 1590
rect 12645 1590 12740 1630
rect 12645 1570 12715 1590
rect 12430 1555 12486 1561
rect 12430 1495 12434 1555
rect 12515 1545 12715 1570
rect 12770 1561 12800 1749
rect 12744 1555 12800 1561
rect 12486 1495 12744 1515
rect 12796 1495 12800 1555
rect 12430 1485 12800 1495
rect 12830 1815 13200 1825
rect 12830 1755 12834 1815
rect 12886 1795 13144 1815
rect 12830 1749 12886 1755
rect 12830 1561 12860 1749
rect 12915 1740 13115 1765
rect 13196 1755 13200 1815
rect 13144 1749 13200 1755
rect 12915 1720 12985 1740
rect 12890 1680 12985 1720
rect 13045 1720 13115 1740
rect 13045 1680 13140 1720
rect 12890 1630 13140 1680
rect 12890 1590 12985 1630
rect 12915 1570 12985 1590
rect 13045 1590 13140 1630
rect 13045 1570 13115 1590
rect 12830 1555 12886 1561
rect 12830 1495 12834 1555
rect 12915 1545 13115 1570
rect 13170 1561 13200 1749
rect 13144 1555 13200 1561
rect 12886 1495 13144 1515
rect 13196 1495 13200 1555
rect 12830 1485 13200 1495
rect -370 1445 0 1455
rect -370 1385 -366 1445
rect -314 1425 -56 1445
rect -370 1379 -314 1385
rect -370 1191 -340 1379
rect -285 1370 -85 1395
rect -4 1385 0 1445
rect -56 1379 0 1385
rect -285 1350 -215 1370
rect -310 1310 -215 1350
rect -155 1350 -85 1370
rect -155 1310 -60 1350
rect -310 1260 -60 1310
rect -310 1220 -215 1260
rect -285 1200 -215 1220
rect -155 1220 -60 1260
rect -155 1200 -85 1220
rect -370 1185 -314 1191
rect -370 1125 -366 1185
rect -285 1175 -85 1200
rect -30 1191 0 1379
rect -56 1185 0 1191
rect -314 1125 -56 1145
rect -4 1125 0 1185
rect -370 1115 0 1125
rect 30 1445 400 1455
rect 30 1385 34 1445
rect 86 1425 344 1445
rect 30 1379 86 1385
rect 30 1191 60 1379
rect 115 1370 315 1395
rect 396 1385 400 1445
rect 344 1379 400 1385
rect 115 1350 185 1370
rect 90 1310 185 1350
rect 245 1350 315 1370
rect 245 1310 340 1350
rect 90 1260 340 1310
rect 90 1220 185 1260
rect 115 1200 185 1220
rect 245 1220 340 1260
rect 245 1200 315 1220
rect 30 1185 86 1191
rect 30 1125 34 1185
rect 115 1175 315 1200
rect 370 1191 400 1379
rect 344 1185 400 1191
rect 86 1125 344 1145
rect 396 1125 400 1185
rect 30 1115 400 1125
rect 430 1445 800 1455
rect 430 1385 434 1445
rect 486 1425 744 1445
rect 430 1379 486 1385
rect 430 1191 460 1379
rect 515 1370 715 1395
rect 796 1385 800 1445
rect 744 1379 800 1385
rect 515 1350 585 1370
rect 490 1310 585 1350
rect 645 1350 715 1370
rect 645 1310 740 1350
rect 490 1260 740 1310
rect 490 1220 585 1260
rect 515 1200 585 1220
rect 645 1220 740 1260
rect 645 1200 715 1220
rect 430 1185 486 1191
rect 430 1125 434 1185
rect 515 1175 715 1200
rect 770 1191 800 1379
rect 744 1185 800 1191
rect 486 1125 744 1145
rect 796 1125 800 1185
rect 430 1115 800 1125
rect 830 1445 1200 1455
rect 830 1385 834 1445
rect 886 1425 1144 1445
rect 830 1379 886 1385
rect 830 1191 860 1379
rect 915 1370 1115 1395
rect 1196 1385 1200 1445
rect 1144 1379 1200 1385
rect 915 1350 985 1370
rect 890 1310 985 1350
rect 1045 1350 1115 1370
rect 1045 1310 1140 1350
rect 890 1260 1140 1310
rect 890 1220 985 1260
rect 915 1200 985 1220
rect 1045 1220 1140 1260
rect 1045 1200 1115 1220
rect 830 1185 886 1191
rect 830 1125 834 1185
rect 915 1175 1115 1200
rect 1170 1191 1200 1379
rect 1144 1185 1200 1191
rect 886 1125 1144 1145
rect 1196 1125 1200 1185
rect 830 1115 1200 1125
rect 1230 1445 1600 1455
rect 1230 1385 1234 1445
rect 1286 1425 1544 1445
rect 1230 1379 1286 1385
rect 1230 1191 1260 1379
rect 1315 1370 1515 1395
rect 1596 1385 1600 1445
rect 1544 1379 1600 1385
rect 1315 1350 1385 1370
rect 1290 1310 1385 1350
rect 1445 1350 1515 1370
rect 1445 1310 1540 1350
rect 1290 1260 1540 1310
rect 1290 1220 1385 1260
rect 1315 1200 1385 1220
rect 1445 1220 1540 1260
rect 1445 1200 1515 1220
rect 1230 1185 1286 1191
rect 1230 1125 1234 1185
rect 1315 1175 1515 1200
rect 1570 1191 1600 1379
rect 1544 1185 1600 1191
rect 1286 1125 1544 1145
rect 1596 1125 1600 1185
rect 1230 1115 1600 1125
rect 1630 1445 2000 1455
rect 1630 1385 1634 1445
rect 1686 1425 1944 1445
rect 1630 1379 1686 1385
rect 1630 1191 1660 1379
rect 1715 1370 1915 1395
rect 1996 1385 2000 1445
rect 1944 1379 2000 1385
rect 1715 1350 1785 1370
rect 1690 1310 1785 1350
rect 1845 1350 1915 1370
rect 1845 1310 1940 1350
rect 1690 1260 1940 1310
rect 1690 1220 1785 1260
rect 1715 1200 1785 1220
rect 1845 1220 1940 1260
rect 1845 1200 1915 1220
rect 1630 1185 1686 1191
rect 1630 1125 1634 1185
rect 1715 1175 1915 1200
rect 1970 1191 2000 1379
rect 1944 1185 2000 1191
rect 1686 1125 1944 1145
rect 1996 1125 2000 1185
rect 1630 1115 2000 1125
rect 2030 1445 2400 1455
rect 2030 1385 2034 1445
rect 2086 1425 2344 1445
rect 2030 1379 2086 1385
rect 2030 1191 2060 1379
rect 2115 1370 2315 1395
rect 2396 1385 2400 1445
rect 2344 1379 2400 1385
rect 2115 1350 2185 1370
rect 2090 1310 2185 1350
rect 2245 1350 2315 1370
rect 2245 1310 2340 1350
rect 2090 1260 2340 1310
rect 2090 1220 2185 1260
rect 2115 1200 2185 1220
rect 2245 1220 2340 1260
rect 2245 1200 2315 1220
rect 2030 1185 2086 1191
rect 2030 1125 2034 1185
rect 2115 1175 2315 1200
rect 2370 1191 2400 1379
rect 2344 1185 2400 1191
rect 2086 1125 2344 1145
rect 2396 1125 2400 1185
rect 2030 1115 2400 1125
rect 2430 1445 2800 1455
rect 2430 1385 2434 1445
rect 2486 1425 2744 1445
rect 2430 1379 2486 1385
rect 2430 1191 2460 1379
rect 2515 1370 2715 1395
rect 2796 1385 2800 1445
rect 2744 1379 2800 1385
rect 2515 1350 2585 1370
rect 2490 1310 2585 1350
rect 2645 1350 2715 1370
rect 2645 1310 2740 1350
rect 2490 1260 2740 1310
rect 2490 1220 2585 1260
rect 2515 1200 2585 1220
rect 2645 1220 2740 1260
rect 2645 1200 2715 1220
rect 2430 1185 2486 1191
rect 2430 1125 2434 1185
rect 2515 1175 2715 1200
rect 2770 1191 2800 1379
rect 2744 1185 2800 1191
rect 2486 1125 2744 1145
rect 2796 1125 2800 1185
rect 2430 1115 2800 1125
rect 2830 1445 3200 1455
rect 2830 1385 2834 1445
rect 2886 1425 3144 1445
rect 2830 1379 2886 1385
rect 2830 1191 2860 1379
rect 2915 1370 3115 1395
rect 3196 1385 3200 1445
rect 3144 1379 3200 1385
rect 2915 1350 2985 1370
rect 2890 1310 2985 1350
rect 3045 1350 3115 1370
rect 3045 1310 3140 1350
rect 2890 1260 3140 1310
rect 2890 1220 2985 1260
rect 2915 1200 2985 1220
rect 3045 1220 3140 1260
rect 3045 1200 3115 1220
rect 2830 1185 2886 1191
rect 2830 1125 2834 1185
rect 2915 1175 3115 1200
rect 3170 1191 3200 1379
rect 3144 1185 3200 1191
rect 2886 1125 3144 1145
rect 3196 1125 3200 1185
rect 2830 1115 3200 1125
rect 3230 1445 3600 1455
rect 3230 1385 3234 1445
rect 3286 1425 3544 1445
rect 3230 1379 3286 1385
rect 3230 1191 3260 1379
rect 3315 1370 3515 1395
rect 3596 1385 3600 1445
rect 3544 1379 3600 1385
rect 3315 1350 3385 1370
rect 3290 1310 3385 1350
rect 3445 1350 3515 1370
rect 3445 1310 3540 1350
rect 3290 1260 3540 1310
rect 3290 1220 3385 1260
rect 3315 1200 3385 1220
rect 3445 1220 3540 1260
rect 3445 1200 3515 1220
rect 3230 1185 3286 1191
rect 3230 1125 3234 1185
rect 3315 1175 3515 1200
rect 3570 1191 3600 1379
rect 3544 1185 3600 1191
rect 3286 1125 3544 1145
rect 3596 1125 3600 1185
rect 3230 1115 3600 1125
rect 3630 1445 4000 1455
rect 3630 1385 3634 1445
rect 3686 1425 3944 1445
rect 3630 1379 3686 1385
rect 3630 1191 3660 1379
rect 3715 1370 3915 1395
rect 3996 1385 4000 1445
rect 3944 1379 4000 1385
rect 3715 1350 3785 1370
rect 3690 1310 3785 1350
rect 3845 1350 3915 1370
rect 3845 1310 3940 1350
rect 3690 1260 3940 1310
rect 3690 1220 3785 1260
rect 3715 1200 3785 1220
rect 3845 1220 3940 1260
rect 3845 1200 3915 1220
rect 3630 1185 3686 1191
rect 3630 1125 3634 1185
rect 3715 1175 3915 1200
rect 3970 1191 4000 1379
rect 3944 1185 4000 1191
rect 3686 1125 3944 1145
rect 3996 1125 4000 1185
rect 3630 1115 4000 1125
rect 4030 1445 4400 1455
rect 4030 1385 4034 1445
rect 4086 1425 4344 1445
rect 4030 1379 4086 1385
rect 4030 1191 4060 1379
rect 4115 1370 4315 1395
rect 4396 1385 4400 1445
rect 4344 1379 4400 1385
rect 4115 1350 4185 1370
rect 4090 1310 4185 1350
rect 4245 1350 4315 1370
rect 4245 1310 4340 1350
rect 4090 1260 4340 1310
rect 4090 1220 4185 1260
rect 4115 1200 4185 1220
rect 4245 1220 4340 1260
rect 4245 1200 4315 1220
rect 4030 1185 4086 1191
rect 4030 1125 4034 1185
rect 4115 1175 4315 1200
rect 4370 1191 4400 1379
rect 4344 1185 4400 1191
rect 4086 1125 4344 1145
rect 4396 1125 4400 1185
rect 4030 1115 4400 1125
rect 4430 1445 4800 1455
rect 4430 1385 4434 1445
rect 4486 1425 4744 1445
rect 4430 1379 4486 1385
rect 4430 1191 4460 1379
rect 4515 1370 4715 1395
rect 4796 1385 4800 1445
rect 4744 1379 4800 1385
rect 4515 1350 4585 1370
rect 4490 1310 4585 1350
rect 4645 1350 4715 1370
rect 4645 1310 4740 1350
rect 4490 1260 4740 1310
rect 4490 1220 4585 1260
rect 4515 1200 4585 1220
rect 4645 1220 4740 1260
rect 4645 1200 4715 1220
rect 4430 1185 4486 1191
rect 4430 1125 4434 1185
rect 4515 1175 4715 1200
rect 4770 1191 4800 1379
rect 4744 1185 4800 1191
rect 4486 1125 4744 1145
rect 4796 1125 4800 1185
rect 4430 1115 4800 1125
rect 4830 1445 5200 1455
rect 4830 1385 4834 1445
rect 4886 1425 5144 1445
rect 4830 1379 4886 1385
rect 4830 1191 4860 1379
rect 4915 1370 5115 1395
rect 5196 1385 5200 1445
rect 5144 1379 5200 1385
rect 4915 1350 4985 1370
rect 4890 1310 4985 1350
rect 5045 1350 5115 1370
rect 5045 1310 5140 1350
rect 4890 1260 5140 1310
rect 4890 1220 4985 1260
rect 4915 1200 4985 1220
rect 5045 1220 5140 1260
rect 5045 1200 5115 1220
rect 4830 1185 4886 1191
rect 4830 1125 4834 1185
rect 4915 1175 5115 1200
rect 5170 1191 5200 1379
rect 5144 1185 5200 1191
rect 4886 1125 5144 1145
rect 5196 1125 5200 1185
rect 4830 1115 5200 1125
rect 5230 1445 5600 1455
rect 5230 1385 5234 1445
rect 5286 1425 5544 1445
rect 5230 1379 5286 1385
rect 5230 1191 5260 1379
rect 5315 1370 5515 1395
rect 5596 1385 5600 1445
rect 5544 1379 5600 1385
rect 5315 1350 5385 1370
rect 5290 1310 5385 1350
rect 5445 1350 5515 1370
rect 5445 1310 5540 1350
rect 5290 1260 5540 1310
rect 5290 1220 5385 1260
rect 5315 1200 5385 1220
rect 5445 1220 5540 1260
rect 5445 1200 5515 1220
rect 5230 1185 5286 1191
rect 5230 1125 5234 1185
rect 5315 1175 5515 1200
rect 5570 1191 5600 1379
rect 5544 1185 5600 1191
rect 5286 1125 5544 1145
rect 5596 1125 5600 1185
rect 5230 1115 5600 1125
rect 5630 1445 6000 1455
rect 5630 1385 5634 1445
rect 5686 1425 5944 1445
rect 5630 1379 5686 1385
rect 5630 1191 5660 1379
rect 5715 1370 5915 1395
rect 5996 1385 6000 1445
rect 5944 1379 6000 1385
rect 5715 1350 5785 1370
rect 5690 1310 5785 1350
rect 5845 1350 5915 1370
rect 5845 1310 5940 1350
rect 5690 1260 5940 1310
rect 5690 1220 5785 1260
rect 5715 1200 5785 1220
rect 5845 1220 5940 1260
rect 5845 1200 5915 1220
rect 5630 1185 5686 1191
rect 5630 1125 5634 1185
rect 5715 1175 5915 1200
rect 5970 1191 6000 1379
rect 5944 1185 6000 1191
rect 5686 1125 5944 1145
rect 5996 1125 6000 1185
rect 5630 1115 6000 1125
rect 6030 1445 6400 1455
rect 6030 1385 6034 1445
rect 6086 1425 6344 1445
rect 6030 1379 6086 1385
rect 6030 1191 6060 1379
rect 6115 1370 6315 1395
rect 6396 1385 6400 1445
rect 6344 1379 6400 1385
rect 6115 1350 6185 1370
rect 6090 1310 6185 1350
rect 6245 1350 6315 1370
rect 6245 1310 6340 1350
rect 6090 1260 6340 1310
rect 6090 1220 6185 1260
rect 6115 1200 6185 1220
rect 6245 1220 6340 1260
rect 6245 1200 6315 1220
rect 6030 1185 6086 1191
rect 6030 1125 6034 1185
rect 6115 1175 6315 1200
rect 6370 1191 6400 1379
rect 6344 1185 6400 1191
rect 6086 1125 6344 1145
rect 6396 1125 6400 1185
rect 6030 1115 6400 1125
rect 6430 1445 6800 1455
rect 6430 1385 6434 1445
rect 6486 1425 6744 1445
rect 6430 1379 6486 1385
rect 6430 1191 6460 1379
rect 6515 1370 6715 1395
rect 6796 1385 6800 1445
rect 6744 1379 6800 1385
rect 6515 1350 6585 1370
rect 6490 1310 6585 1350
rect 6645 1350 6715 1370
rect 6645 1310 6740 1350
rect 6490 1260 6740 1310
rect 6490 1220 6585 1260
rect 6515 1200 6585 1220
rect 6645 1220 6740 1260
rect 6645 1200 6715 1220
rect 6430 1185 6486 1191
rect 6430 1125 6434 1185
rect 6515 1175 6715 1200
rect 6770 1191 6800 1379
rect 6744 1185 6800 1191
rect 6486 1125 6744 1145
rect 6796 1125 6800 1185
rect 6430 1115 6800 1125
rect 6830 1445 7200 1455
rect 6830 1385 6834 1445
rect 6886 1425 7144 1445
rect 6830 1379 6886 1385
rect 6830 1191 6860 1379
rect 6915 1370 7115 1395
rect 7196 1385 7200 1445
rect 7144 1379 7200 1385
rect 6915 1350 6985 1370
rect 6890 1310 6985 1350
rect 7045 1350 7115 1370
rect 7045 1310 7140 1350
rect 6890 1260 7140 1310
rect 6890 1220 6985 1260
rect 6915 1200 6985 1220
rect 7045 1220 7140 1260
rect 7045 1200 7115 1220
rect 6830 1185 6886 1191
rect 6830 1125 6834 1185
rect 6915 1175 7115 1200
rect 7170 1191 7200 1379
rect 7144 1185 7200 1191
rect 6886 1125 7144 1145
rect 7196 1125 7200 1185
rect 6830 1115 7200 1125
rect 7230 1445 7600 1455
rect 7230 1385 7234 1445
rect 7286 1425 7544 1445
rect 7230 1379 7286 1385
rect 7230 1191 7260 1379
rect 7315 1370 7515 1395
rect 7596 1385 7600 1445
rect 7544 1379 7600 1385
rect 7315 1350 7385 1370
rect 7290 1310 7385 1350
rect 7445 1350 7515 1370
rect 7445 1310 7540 1350
rect 7290 1260 7540 1310
rect 7290 1220 7385 1260
rect 7315 1200 7385 1220
rect 7445 1220 7540 1260
rect 7445 1200 7515 1220
rect 7230 1185 7286 1191
rect 7230 1125 7234 1185
rect 7315 1175 7515 1200
rect 7570 1191 7600 1379
rect 7544 1185 7600 1191
rect 7286 1125 7544 1145
rect 7596 1125 7600 1185
rect 7230 1115 7600 1125
rect 7630 1445 8000 1455
rect 7630 1385 7634 1445
rect 7686 1425 7944 1445
rect 7630 1379 7686 1385
rect 7630 1191 7660 1379
rect 7715 1370 7915 1395
rect 7996 1385 8000 1445
rect 7944 1379 8000 1385
rect 7715 1350 7785 1370
rect 7690 1310 7785 1350
rect 7845 1350 7915 1370
rect 7845 1310 7940 1350
rect 7690 1260 7940 1310
rect 7690 1220 7785 1260
rect 7715 1200 7785 1220
rect 7845 1220 7940 1260
rect 7845 1200 7915 1220
rect 7630 1185 7686 1191
rect 7630 1125 7634 1185
rect 7715 1175 7915 1200
rect 7970 1191 8000 1379
rect 7944 1185 8000 1191
rect 7686 1125 7944 1145
rect 7996 1125 8000 1185
rect 7630 1115 8000 1125
rect 8030 1445 8400 1455
rect 8030 1385 8034 1445
rect 8086 1425 8344 1445
rect 8030 1379 8086 1385
rect 8030 1191 8060 1379
rect 8115 1370 8315 1395
rect 8396 1385 8400 1445
rect 8344 1379 8400 1385
rect 8115 1350 8185 1370
rect 8090 1310 8185 1350
rect 8245 1350 8315 1370
rect 8245 1310 8340 1350
rect 8090 1260 8340 1310
rect 8090 1220 8185 1260
rect 8115 1200 8185 1220
rect 8245 1220 8340 1260
rect 8245 1200 8315 1220
rect 8030 1185 8086 1191
rect 8030 1125 8034 1185
rect 8115 1175 8315 1200
rect 8370 1191 8400 1379
rect 8344 1185 8400 1191
rect 8086 1125 8344 1145
rect 8396 1125 8400 1185
rect 8030 1115 8400 1125
rect 8430 1445 8800 1455
rect 8430 1385 8434 1445
rect 8486 1425 8744 1445
rect 8430 1379 8486 1385
rect 8430 1191 8460 1379
rect 8515 1370 8715 1395
rect 8796 1385 8800 1445
rect 8744 1379 8800 1385
rect 8515 1350 8585 1370
rect 8490 1310 8585 1350
rect 8645 1350 8715 1370
rect 8645 1310 8740 1350
rect 8490 1260 8740 1310
rect 8490 1220 8585 1260
rect 8515 1200 8585 1220
rect 8645 1220 8740 1260
rect 8645 1200 8715 1220
rect 8430 1185 8486 1191
rect 8430 1125 8434 1185
rect 8515 1175 8715 1200
rect 8770 1191 8800 1379
rect 8744 1185 8800 1191
rect 8486 1125 8744 1145
rect 8796 1125 8800 1185
rect 8430 1115 8800 1125
rect 8830 1445 9200 1455
rect 8830 1385 8834 1445
rect 8886 1425 9144 1445
rect 8830 1379 8886 1385
rect 8830 1191 8860 1379
rect 8915 1370 9115 1395
rect 9196 1385 9200 1445
rect 9144 1379 9200 1385
rect 8915 1350 8985 1370
rect 8890 1310 8985 1350
rect 9045 1350 9115 1370
rect 9045 1310 9140 1350
rect 8890 1260 9140 1310
rect 8890 1220 8985 1260
rect 8915 1200 8985 1220
rect 9045 1220 9140 1260
rect 9045 1200 9115 1220
rect 8830 1185 8886 1191
rect 8830 1125 8834 1185
rect 8915 1175 9115 1200
rect 9170 1191 9200 1379
rect 9144 1185 9200 1191
rect 8886 1125 9144 1145
rect 9196 1125 9200 1185
rect 8830 1115 9200 1125
rect 9230 1445 9600 1455
rect 9230 1385 9234 1445
rect 9286 1425 9544 1445
rect 9230 1379 9286 1385
rect 9230 1191 9260 1379
rect 9315 1370 9515 1395
rect 9596 1385 9600 1445
rect 9544 1379 9600 1385
rect 9315 1350 9385 1370
rect 9290 1310 9385 1350
rect 9445 1350 9515 1370
rect 9445 1310 9540 1350
rect 9290 1260 9540 1310
rect 9290 1220 9385 1260
rect 9315 1200 9385 1220
rect 9445 1220 9540 1260
rect 9445 1200 9515 1220
rect 9230 1185 9286 1191
rect 9230 1125 9234 1185
rect 9315 1175 9515 1200
rect 9570 1191 9600 1379
rect 9544 1185 9600 1191
rect 9286 1125 9544 1145
rect 9596 1125 9600 1185
rect 9230 1115 9600 1125
rect 9630 1445 10000 1455
rect 9630 1385 9634 1445
rect 9686 1425 9944 1445
rect 9630 1379 9686 1385
rect 9630 1191 9660 1379
rect 9715 1370 9915 1395
rect 9996 1385 10000 1445
rect 9944 1379 10000 1385
rect 9715 1350 9785 1370
rect 9690 1310 9785 1350
rect 9845 1350 9915 1370
rect 9845 1310 9940 1350
rect 9690 1260 9940 1310
rect 9690 1220 9785 1260
rect 9715 1200 9785 1220
rect 9845 1220 9940 1260
rect 9845 1200 9915 1220
rect 9630 1185 9686 1191
rect 9630 1125 9634 1185
rect 9715 1175 9915 1200
rect 9970 1191 10000 1379
rect 9944 1185 10000 1191
rect 9686 1125 9944 1145
rect 9996 1125 10000 1185
rect 9630 1115 10000 1125
rect 10030 1445 10400 1455
rect 10030 1385 10034 1445
rect 10086 1425 10344 1445
rect 10030 1379 10086 1385
rect 10030 1191 10060 1379
rect 10115 1370 10315 1395
rect 10396 1385 10400 1445
rect 10344 1379 10400 1385
rect 10115 1350 10185 1370
rect 10090 1310 10185 1350
rect 10245 1350 10315 1370
rect 10245 1310 10340 1350
rect 10090 1260 10340 1310
rect 10090 1220 10185 1260
rect 10115 1200 10185 1220
rect 10245 1220 10340 1260
rect 10245 1200 10315 1220
rect 10030 1185 10086 1191
rect 10030 1125 10034 1185
rect 10115 1175 10315 1200
rect 10370 1191 10400 1379
rect 10344 1185 10400 1191
rect 10086 1125 10344 1145
rect 10396 1125 10400 1185
rect 10030 1115 10400 1125
rect 10430 1445 10800 1455
rect 10430 1385 10434 1445
rect 10486 1425 10744 1445
rect 10430 1379 10486 1385
rect 10430 1191 10460 1379
rect 10515 1370 10715 1395
rect 10796 1385 10800 1445
rect 10744 1379 10800 1385
rect 10515 1350 10585 1370
rect 10490 1310 10585 1350
rect 10645 1350 10715 1370
rect 10645 1310 10740 1350
rect 10490 1260 10740 1310
rect 10490 1220 10585 1260
rect 10515 1200 10585 1220
rect 10645 1220 10740 1260
rect 10645 1200 10715 1220
rect 10430 1185 10486 1191
rect 10430 1125 10434 1185
rect 10515 1175 10715 1200
rect 10770 1191 10800 1379
rect 10744 1185 10800 1191
rect 10486 1125 10744 1145
rect 10796 1125 10800 1185
rect 10430 1115 10800 1125
rect 10830 1445 11200 1455
rect 10830 1385 10834 1445
rect 10886 1425 11144 1445
rect 10830 1379 10886 1385
rect 10830 1191 10860 1379
rect 10915 1370 11115 1395
rect 11196 1385 11200 1445
rect 11144 1379 11200 1385
rect 10915 1350 10985 1370
rect 10890 1310 10985 1350
rect 11045 1350 11115 1370
rect 11045 1310 11140 1350
rect 10890 1260 11140 1310
rect 10890 1220 10985 1260
rect 10915 1200 10985 1220
rect 11045 1220 11140 1260
rect 11045 1200 11115 1220
rect 10830 1185 10886 1191
rect 10830 1125 10834 1185
rect 10915 1175 11115 1200
rect 11170 1191 11200 1379
rect 11144 1185 11200 1191
rect 10886 1125 11144 1145
rect 11196 1125 11200 1185
rect 10830 1115 11200 1125
rect 11230 1445 11600 1455
rect 11230 1385 11234 1445
rect 11286 1425 11544 1445
rect 11230 1379 11286 1385
rect 11230 1191 11260 1379
rect 11315 1370 11515 1395
rect 11596 1385 11600 1445
rect 11544 1379 11600 1385
rect 11315 1350 11385 1370
rect 11290 1310 11385 1350
rect 11445 1350 11515 1370
rect 11445 1310 11540 1350
rect 11290 1260 11540 1310
rect 11290 1220 11385 1260
rect 11315 1200 11385 1220
rect 11445 1220 11540 1260
rect 11445 1200 11515 1220
rect 11230 1185 11286 1191
rect 11230 1125 11234 1185
rect 11315 1175 11515 1200
rect 11570 1191 11600 1379
rect 11544 1185 11600 1191
rect 11286 1125 11544 1145
rect 11596 1125 11600 1185
rect 11230 1115 11600 1125
rect 11630 1445 12000 1455
rect 11630 1385 11634 1445
rect 11686 1425 11944 1445
rect 11630 1379 11686 1385
rect 11630 1191 11660 1379
rect 11715 1370 11915 1395
rect 11996 1385 12000 1445
rect 11944 1379 12000 1385
rect 11715 1350 11785 1370
rect 11690 1310 11785 1350
rect 11845 1350 11915 1370
rect 11845 1310 11940 1350
rect 11690 1260 11940 1310
rect 11690 1220 11785 1260
rect 11715 1200 11785 1220
rect 11845 1220 11940 1260
rect 11845 1200 11915 1220
rect 11630 1185 11686 1191
rect 11630 1125 11634 1185
rect 11715 1175 11915 1200
rect 11970 1191 12000 1379
rect 11944 1185 12000 1191
rect 11686 1125 11944 1145
rect 11996 1125 12000 1185
rect 11630 1115 12000 1125
rect 12030 1445 12400 1455
rect 12030 1385 12034 1445
rect 12086 1425 12344 1445
rect 12030 1379 12086 1385
rect 12030 1191 12060 1379
rect 12115 1370 12315 1395
rect 12396 1385 12400 1445
rect 12344 1379 12400 1385
rect 12115 1350 12185 1370
rect 12090 1310 12185 1350
rect 12245 1350 12315 1370
rect 12245 1310 12340 1350
rect 12090 1260 12340 1310
rect 12090 1220 12185 1260
rect 12115 1200 12185 1220
rect 12245 1220 12340 1260
rect 12245 1200 12315 1220
rect 12030 1185 12086 1191
rect 12030 1125 12034 1185
rect 12115 1175 12315 1200
rect 12370 1191 12400 1379
rect 12344 1185 12400 1191
rect 12086 1125 12344 1145
rect 12396 1125 12400 1185
rect 12030 1115 12400 1125
rect 12430 1445 12800 1455
rect 12430 1385 12434 1445
rect 12486 1425 12744 1445
rect 12430 1379 12486 1385
rect 12430 1191 12460 1379
rect 12515 1370 12715 1395
rect 12796 1385 12800 1445
rect 12744 1379 12800 1385
rect 12515 1350 12585 1370
rect 12490 1310 12585 1350
rect 12645 1350 12715 1370
rect 12645 1310 12740 1350
rect 12490 1260 12740 1310
rect 12490 1220 12585 1260
rect 12515 1200 12585 1220
rect 12645 1220 12740 1260
rect 12645 1200 12715 1220
rect 12430 1185 12486 1191
rect 12430 1125 12434 1185
rect 12515 1175 12715 1200
rect 12770 1191 12800 1379
rect 12744 1185 12800 1191
rect 12486 1125 12744 1145
rect 12796 1125 12800 1185
rect 12430 1115 12800 1125
rect 12830 1445 13200 1455
rect 12830 1385 12834 1445
rect 12886 1425 13144 1445
rect 12830 1379 12886 1385
rect 12830 1191 12860 1379
rect 12915 1370 13115 1395
rect 13196 1385 13200 1445
rect 13144 1379 13200 1385
rect 12915 1350 12985 1370
rect 12890 1310 12985 1350
rect 13045 1350 13115 1370
rect 13045 1310 13140 1350
rect 12890 1260 13140 1310
rect 12890 1220 12985 1260
rect 12915 1200 12985 1220
rect 13045 1220 13140 1260
rect 13045 1200 13115 1220
rect 12830 1185 12886 1191
rect 12830 1125 12834 1185
rect 12915 1175 13115 1200
rect 13170 1191 13200 1379
rect 13144 1185 13200 1191
rect 12886 1125 13144 1145
rect 13196 1125 13200 1185
rect 12830 1115 13200 1125
rect -370 1075 0 1085
rect -370 1015 -366 1075
rect -314 1055 -56 1075
rect -370 1009 -314 1015
rect -370 821 -340 1009
rect -285 1000 -85 1025
rect -4 1015 0 1075
rect -56 1009 0 1015
rect -285 980 -215 1000
rect -310 940 -215 980
rect -155 980 -85 1000
rect -155 940 -60 980
rect -310 890 -60 940
rect -310 850 -215 890
rect -285 830 -215 850
rect -155 850 -60 890
rect -155 830 -85 850
rect -370 815 -314 821
rect -370 755 -366 815
rect -285 805 -85 830
rect -30 821 0 1009
rect -56 815 0 821
rect -314 755 -56 775
rect -4 755 0 815
rect -370 745 0 755
rect 30 1075 400 1085
rect 30 1015 34 1075
rect 86 1055 344 1075
rect 30 1009 86 1015
rect 30 821 60 1009
rect 115 1000 315 1025
rect 396 1015 400 1075
rect 344 1009 400 1015
rect 115 980 185 1000
rect 90 940 185 980
rect 245 980 315 1000
rect 245 940 340 980
rect 90 890 340 940
rect 90 850 185 890
rect 115 830 185 850
rect 245 850 340 890
rect 245 830 315 850
rect 30 815 86 821
rect 30 755 34 815
rect 115 805 315 830
rect 370 821 400 1009
rect 344 815 400 821
rect 86 755 344 775
rect 396 755 400 815
rect 30 745 400 755
rect 430 1075 800 1085
rect 430 1015 434 1075
rect 486 1055 744 1075
rect 430 1009 486 1015
rect 430 821 460 1009
rect 515 1000 715 1025
rect 796 1015 800 1075
rect 744 1009 800 1015
rect 515 980 585 1000
rect 490 940 585 980
rect 645 980 715 1000
rect 645 940 740 980
rect 490 890 740 940
rect 490 850 585 890
rect 515 830 585 850
rect 645 850 740 890
rect 645 830 715 850
rect 430 815 486 821
rect 430 755 434 815
rect 515 805 715 830
rect 770 821 800 1009
rect 744 815 800 821
rect 486 755 744 775
rect 796 755 800 815
rect 430 745 800 755
rect 830 1075 1200 1085
rect 830 1015 834 1075
rect 886 1055 1144 1075
rect 830 1009 886 1015
rect 830 821 860 1009
rect 915 1000 1115 1025
rect 1196 1015 1200 1075
rect 1144 1009 1200 1015
rect 915 980 985 1000
rect 890 940 985 980
rect 1045 980 1115 1000
rect 1045 940 1140 980
rect 890 890 1140 940
rect 890 850 985 890
rect 915 830 985 850
rect 1045 850 1140 890
rect 1045 830 1115 850
rect 830 815 886 821
rect 830 755 834 815
rect 915 805 1115 830
rect 1170 821 1200 1009
rect 1144 815 1200 821
rect 886 755 1144 775
rect 1196 755 1200 815
rect 830 745 1200 755
rect 1230 1075 1600 1085
rect 1230 1015 1234 1075
rect 1286 1055 1544 1075
rect 1230 1009 1286 1015
rect 1230 821 1260 1009
rect 1315 1000 1515 1025
rect 1596 1015 1600 1075
rect 1544 1009 1600 1015
rect 1315 980 1385 1000
rect 1290 940 1385 980
rect 1445 980 1515 1000
rect 1445 940 1540 980
rect 1290 890 1540 940
rect 1290 850 1385 890
rect 1315 830 1385 850
rect 1445 850 1540 890
rect 1445 830 1515 850
rect 1230 815 1286 821
rect 1230 755 1234 815
rect 1315 805 1515 830
rect 1570 821 1600 1009
rect 1544 815 1600 821
rect 1286 755 1544 775
rect 1596 755 1600 815
rect 1230 745 1600 755
rect 1630 1075 2000 1085
rect 1630 1015 1634 1075
rect 1686 1055 1944 1075
rect 1630 1009 1686 1015
rect 1630 821 1660 1009
rect 1715 1000 1915 1025
rect 1996 1015 2000 1075
rect 1944 1009 2000 1015
rect 1715 980 1785 1000
rect 1690 940 1785 980
rect 1845 980 1915 1000
rect 1845 940 1940 980
rect 1690 890 1940 940
rect 1690 850 1785 890
rect 1715 830 1785 850
rect 1845 850 1940 890
rect 1845 830 1915 850
rect 1630 815 1686 821
rect 1630 755 1634 815
rect 1715 805 1915 830
rect 1970 821 2000 1009
rect 1944 815 2000 821
rect 1686 755 1944 775
rect 1996 755 2000 815
rect 1630 745 2000 755
rect 2030 1075 2400 1085
rect 2030 1015 2034 1075
rect 2086 1055 2344 1075
rect 2030 1009 2086 1015
rect 2030 821 2060 1009
rect 2115 1000 2315 1025
rect 2396 1015 2400 1075
rect 2344 1009 2400 1015
rect 2115 980 2185 1000
rect 2090 940 2185 980
rect 2245 980 2315 1000
rect 2245 940 2340 980
rect 2090 890 2340 940
rect 2090 850 2185 890
rect 2115 830 2185 850
rect 2245 850 2340 890
rect 2245 830 2315 850
rect 2030 815 2086 821
rect 2030 755 2034 815
rect 2115 805 2315 830
rect 2370 821 2400 1009
rect 2344 815 2400 821
rect 2086 755 2344 775
rect 2396 755 2400 815
rect 2030 745 2400 755
rect 2430 1075 2800 1085
rect 2430 1015 2434 1075
rect 2486 1055 2744 1075
rect 2430 1009 2486 1015
rect 2430 821 2460 1009
rect 2515 1000 2715 1025
rect 2796 1015 2800 1075
rect 2744 1009 2800 1015
rect 2515 980 2585 1000
rect 2490 940 2585 980
rect 2645 980 2715 1000
rect 2645 940 2740 980
rect 2490 890 2740 940
rect 2490 850 2585 890
rect 2515 830 2585 850
rect 2645 850 2740 890
rect 2645 830 2715 850
rect 2430 815 2486 821
rect 2430 755 2434 815
rect 2515 805 2715 830
rect 2770 821 2800 1009
rect 2744 815 2800 821
rect 2486 755 2744 775
rect 2796 755 2800 815
rect 2430 745 2800 755
rect 2830 1075 3200 1085
rect 2830 1015 2834 1075
rect 2886 1055 3144 1075
rect 2830 1009 2886 1015
rect 2830 821 2860 1009
rect 2915 1000 3115 1025
rect 3196 1015 3200 1075
rect 3144 1009 3200 1015
rect 2915 980 2985 1000
rect 2890 940 2985 980
rect 3045 980 3115 1000
rect 3045 940 3140 980
rect 2890 890 3140 940
rect 2890 850 2985 890
rect 2915 830 2985 850
rect 3045 850 3140 890
rect 3045 830 3115 850
rect 2830 815 2886 821
rect 2830 755 2834 815
rect 2915 805 3115 830
rect 3170 821 3200 1009
rect 3144 815 3200 821
rect 2886 755 3144 775
rect 3196 755 3200 815
rect 2830 745 3200 755
rect 3230 1075 3600 1085
rect 3230 1015 3234 1075
rect 3286 1055 3544 1075
rect 3230 1009 3286 1015
rect 3230 821 3260 1009
rect 3315 1000 3515 1025
rect 3596 1015 3600 1075
rect 3544 1009 3600 1015
rect 3315 980 3385 1000
rect 3290 940 3385 980
rect 3445 980 3515 1000
rect 3445 940 3540 980
rect 3290 890 3540 940
rect 3290 850 3385 890
rect 3315 830 3385 850
rect 3445 850 3540 890
rect 3445 830 3515 850
rect 3230 815 3286 821
rect 3230 755 3234 815
rect 3315 805 3515 830
rect 3570 821 3600 1009
rect 3544 815 3600 821
rect 3286 755 3544 775
rect 3596 755 3600 815
rect 3230 745 3600 755
rect 3630 1075 4000 1085
rect 3630 1015 3634 1075
rect 3686 1055 3944 1075
rect 3630 1009 3686 1015
rect 3630 821 3660 1009
rect 3715 1000 3915 1025
rect 3996 1015 4000 1075
rect 3944 1009 4000 1015
rect 3715 980 3785 1000
rect 3690 940 3785 980
rect 3845 980 3915 1000
rect 3845 940 3940 980
rect 3690 890 3940 940
rect 3690 850 3785 890
rect 3715 830 3785 850
rect 3845 850 3940 890
rect 3845 830 3915 850
rect 3630 815 3686 821
rect 3630 755 3634 815
rect 3715 805 3915 830
rect 3970 821 4000 1009
rect 3944 815 4000 821
rect 3686 755 3944 775
rect 3996 755 4000 815
rect 3630 745 4000 755
rect 4030 1075 4400 1085
rect 4030 1015 4034 1075
rect 4086 1055 4344 1075
rect 4030 1009 4086 1015
rect 4030 821 4060 1009
rect 4115 1000 4315 1025
rect 4396 1015 4400 1075
rect 4344 1009 4400 1015
rect 4115 980 4185 1000
rect 4090 940 4185 980
rect 4245 980 4315 1000
rect 4245 940 4340 980
rect 4090 890 4340 940
rect 4090 850 4185 890
rect 4115 830 4185 850
rect 4245 850 4340 890
rect 4245 830 4315 850
rect 4030 815 4086 821
rect 4030 755 4034 815
rect 4115 805 4315 830
rect 4370 821 4400 1009
rect 4344 815 4400 821
rect 4086 755 4344 775
rect 4396 755 4400 815
rect 4030 745 4400 755
rect 4430 1075 4800 1085
rect 4430 1015 4434 1075
rect 4486 1055 4744 1075
rect 4430 1009 4486 1015
rect 4430 821 4460 1009
rect 4515 1000 4715 1025
rect 4796 1015 4800 1075
rect 4744 1009 4800 1015
rect 4515 980 4585 1000
rect 4490 940 4585 980
rect 4645 980 4715 1000
rect 4645 940 4740 980
rect 4490 890 4740 940
rect 4490 850 4585 890
rect 4515 830 4585 850
rect 4645 850 4740 890
rect 4645 830 4715 850
rect 4430 815 4486 821
rect 4430 755 4434 815
rect 4515 805 4715 830
rect 4770 821 4800 1009
rect 4744 815 4800 821
rect 4486 755 4744 775
rect 4796 755 4800 815
rect 4430 745 4800 755
rect 4830 1075 5200 1085
rect 4830 1015 4834 1075
rect 4886 1055 5144 1075
rect 4830 1009 4886 1015
rect 4830 821 4860 1009
rect 4915 1000 5115 1025
rect 5196 1015 5200 1075
rect 5144 1009 5200 1015
rect 4915 980 4985 1000
rect 4890 940 4985 980
rect 5045 980 5115 1000
rect 5045 940 5140 980
rect 4890 890 5140 940
rect 4890 850 4985 890
rect 4915 830 4985 850
rect 5045 850 5140 890
rect 5045 830 5115 850
rect 4830 815 4886 821
rect 4830 755 4834 815
rect 4915 805 5115 830
rect 5170 821 5200 1009
rect 5144 815 5200 821
rect 4886 755 5144 775
rect 5196 755 5200 815
rect 4830 745 5200 755
rect 5230 1075 5600 1085
rect 5230 1015 5234 1075
rect 5286 1055 5544 1075
rect 5230 1009 5286 1015
rect 5230 821 5260 1009
rect 5315 1000 5515 1025
rect 5596 1015 5600 1075
rect 5544 1009 5600 1015
rect 5315 980 5385 1000
rect 5290 940 5385 980
rect 5445 980 5515 1000
rect 5445 940 5540 980
rect 5290 890 5540 940
rect 5290 850 5385 890
rect 5315 830 5385 850
rect 5445 850 5540 890
rect 5445 830 5515 850
rect 5230 815 5286 821
rect 5230 755 5234 815
rect 5315 805 5515 830
rect 5570 821 5600 1009
rect 5544 815 5600 821
rect 5286 755 5544 775
rect 5596 755 5600 815
rect 5230 745 5600 755
rect 5630 1075 6000 1085
rect 5630 1015 5634 1075
rect 5686 1055 5944 1075
rect 5630 1009 5686 1015
rect 5630 821 5660 1009
rect 5715 1000 5915 1025
rect 5996 1015 6000 1075
rect 5944 1009 6000 1015
rect 5715 980 5785 1000
rect 5690 940 5785 980
rect 5845 980 5915 1000
rect 5845 940 5940 980
rect 5690 890 5940 940
rect 5690 850 5785 890
rect 5715 830 5785 850
rect 5845 850 5940 890
rect 5845 830 5915 850
rect 5630 815 5686 821
rect 5630 755 5634 815
rect 5715 805 5915 830
rect 5970 821 6000 1009
rect 5944 815 6000 821
rect 5686 755 5944 775
rect 5996 755 6000 815
rect 5630 745 6000 755
rect 6030 1075 6400 1085
rect 6030 1015 6034 1075
rect 6086 1055 6344 1075
rect 6030 1009 6086 1015
rect 6030 821 6060 1009
rect 6115 1000 6315 1025
rect 6396 1015 6400 1075
rect 6344 1009 6400 1015
rect 6115 980 6185 1000
rect 6090 940 6185 980
rect 6245 980 6315 1000
rect 6245 940 6340 980
rect 6090 890 6340 940
rect 6090 850 6185 890
rect 6115 830 6185 850
rect 6245 850 6340 890
rect 6245 830 6315 850
rect 6030 815 6086 821
rect 6030 755 6034 815
rect 6115 805 6315 830
rect 6370 821 6400 1009
rect 6344 815 6400 821
rect 6086 755 6344 775
rect 6396 755 6400 815
rect 6030 745 6400 755
rect 6430 1075 6800 1085
rect 6430 1015 6434 1075
rect 6486 1055 6744 1075
rect 6430 1009 6486 1015
rect 6430 821 6460 1009
rect 6515 1000 6715 1025
rect 6796 1015 6800 1075
rect 6744 1009 6800 1015
rect 6515 980 6585 1000
rect 6490 940 6585 980
rect 6645 980 6715 1000
rect 6645 940 6740 980
rect 6490 890 6740 940
rect 6490 850 6585 890
rect 6515 830 6585 850
rect 6645 850 6740 890
rect 6645 830 6715 850
rect 6430 815 6486 821
rect 6430 755 6434 815
rect 6515 805 6715 830
rect 6770 821 6800 1009
rect 6744 815 6800 821
rect 6486 755 6744 775
rect 6796 755 6800 815
rect 6430 745 6800 755
rect 6830 1075 7200 1085
rect 6830 1015 6834 1075
rect 6886 1055 7144 1075
rect 6830 1009 6886 1015
rect 6830 821 6860 1009
rect 6915 1000 7115 1025
rect 7196 1015 7200 1075
rect 7144 1009 7200 1015
rect 6915 980 6985 1000
rect 6890 940 6985 980
rect 7045 980 7115 1000
rect 7045 940 7140 980
rect 6890 890 7140 940
rect 6890 850 6985 890
rect 6915 830 6985 850
rect 7045 850 7140 890
rect 7045 830 7115 850
rect 6830 815 6886 821
rect 6830 755 6834 815
rect 6915 805 7115 830
rect 7170 821 7200 1009
rect 7144 815 7200 821
rect 6886 755 7144 775
rect 7196 755 7200 815
rect 6830 745 7200 755
rect 7230 1075 7600 1085
rect 7230 1015 7234 1075
rect 7286 1055 7544 1075
rect 7230 1009 7286 1015
rect 7230 821 7260 1009
rect 7315 1000 7515 1025
rect 7596 1015 7600 1075
rect 7544 1009 7600 1015
rect 7315 980 7385 1000
rect 7290 940 7385 980
rect 7445 980 7515 1000
rect 7445 940 7540 980
rect 7290 890 7540 940
rect 7290 850 7385 890
rect 7315 830 7385 850
rect 7445 850 7540 890
rect 7445 830 7515 850
rect 7230 815 7286 821
rect 7230 755 7234 815
rect 7315 805 7515 830
rect 7570 821 7600 1009
rect 7544 815 7600 821
rect 7286 755 7544 775
rect 7596 755 7600 815
rect 7230 745 7600 755
rect 7630 1075 8000 1085
rect 7630 1015 7634 1075
rect 7686 1055 7944 1075
rect 7630 1009 7686 1015
rect 7630 821 7660 1009
rect 7715 1000 7915 1025
rect 7996 1015 8000 1075
rect 7944 1009 8000 1015
rect 7715 980 7785 1000
rect 7690 940 7785 980
rect 7845 980 7915 1000
rect 7845 940 7940 980
rect 7690 890 7940 940
rect 7690 850 7785 890
rect 7715 830 7785 850
rect 7845 850 7940 890
rect 7845 830 7915 850
rect 7630 815 7686 821
rect 7630 755 7634 815
rect 7715 805 7915 830
rect 7970 821 8000 1009
rect 7944 815 8000 821
rect 7686 755 7944 775
rect 7996 755 8000 815
rect 7630 745 8000 755
rect 8030 1075 8400 1085
rect 8030 1015 8034 1075
rect 8086 1055 8344 1075
rect 8030 1009 8086 1015
rect 8030 821 8060 1009
rect 8115 1000 8315 1025
rect 8396 1015 8400 1075
rect 8344 1009 8400 1015
rect 8115 980 8185 1000
rect 8090 940 8185 980
rect 8245 980 8315 1000
rect 8245 940 8340 980
rect 8090 890 8340 940
rect 8090 850 8185 890
rect 8115 830 8185 850
rect 8245 850 8340 890
rect 8245 830 8315 850
rect 8030 815 8086 821
rect 8030 755 8034 815
rect 8115 805 8315 830
rect 8370 821 8400 1009
rect 8344 815 8400 821
rect 8086 755 8344 775
rect 8396 755 8400 815
rect 8030 745 8400 755
rect 8430 1075 8800 1085
rect 8430 1015 8434 1075
rect 8486 1055 8744 1075
rect 8430 1009 8486 1015
rect 8430 821 8460 1009
rect 8515 1000 8715 1025
rect 8796 1015 8800 1075
rect 8744 1009 8800 1015
rect 8515 980 8585 1000
rect 8490 940 8585 980
rect 8645 980 8715 1000
rect 8645 940 8740 980
rect 8490 890 8740 940
rect 8490 850 8585 890
rect 8515 830 8585 850
rect 8645 850 8740 890
rect 8645 830 8715 850
rect 8430 815 8486 821
rect 8430 755 8434 815
rect 8515 805 8715 830
rect 8770 821 8800 1009
rect 8744 815 8800 821
rect 8486 755 8744 775
rect 8796 755 8800 815
rect 8430 745 8800 755
rect 8830 1075 9200 1085
rect 8830 1015 8834 1075
rect 8886 1055 9144 1075
rect 8830 1009 8886 1015
rect 8830 821 8860 1009
rect 8915 1000 9115 1025
rect 9196 1015 9200 1075
rect 9144 1009 9200 1015
rect 8915 980 8985 1000
rect 8890 940 8985 980
rect 9045 980 9115 1000
rect 9045 940 9140 980
rect 8890 890 9140 940
rect 8890 850 8985 890
rect 8915 830 8985 850
rect 9045 850 9140 890
rect 9045 830 9115 850
rect 8830 815 8886 821
rect 8830 755 8834 815
rect 8915 805 9115 830
rect 9170 821 9200 1009
rect 9144 815 9200 821
rect 8886 755 9144 775
rect 9196 755 9200 815
rect 8830 745 9200 755
rect 9230 1075 9600 1085
rect 9230 1015 9234 1075
rect 9286 1055 9544 1075
rect 9230 1009 9286 1015
rect 9230 821 9260 1009
rect 9315 1000 9515 1025
rect 9596 1015 9600 1075
rect 9544 1009 9600 1015
rect 9315 980 9385 1000
rect 9290 940 9385 980
rect 9445 980 9515 1000
rect 9445 940 9540 980
rect 9290 890 9540 940
rect 9290 850 9385 890
rect 9315 830 9385 850
rect 9445 850 9540 890
rect 9445 830 9515 850
rect 9230 815 9286 821
rect 9230 755 9234 815
rect 9315 805 9515 830
rect 9570 821 9600 1009
rect 9544 815 9600 821
rect 9286 755 9544 775
rect 9596 755 9600 815
rect 9230 745 9600 755
rect 9630 1075 10000 1085
rect 9630 1015 9634 1075
rect 9686 1055 9944 1075
rect 9630 1009 9686 1015
rect 9630 821 9660 1009
rect 9715 1000 9915 1025
rect 9996 1015 10000 1075
rect 9944 1009 10000 1015
rect 9715 980 9785 1000
rect 9690 940 9785 980
rect 9845 980 9915 1000
rect 9845 940 9940 980
rect 9690 890 9940 940
rect 9690 850 9785 890
rect 9715 830 9785 850
rect 9845 850 9940 890
rect 9845 830 9915 850
rect 9630 815 9686 821
rect 9630 755 9634 815
rect 9715 805 9915 830
rect 9970 821 10000 1009
rect 9944 815 10000 821
rect 9686 755 9944 775
rect 9996 755 10000 815
rect 9630 745 10000 755
rect 10030 1075 10400 1085
rect 10030 1015 10034 1075
rect 10086 1055 10344 1075
rect 10030 1009 10086 1015
rect 10030 821 10060 1009
rect 10115 1000 10315 1025
rect 10396 1015 10400 1075
rect 10344 1009 10400 1015
rect 10115 980 10185 1000
rect 10090 940 10185 980
rect 10245 980 10315 1000
rect 10245 940 10340 980
rect 10090 890 10340 940
rect 10090 850 10185 890
rect 10115 830 10185 850
rect 10245 850 10340 890
rect 10245 830 10315 850
rect 10030 815 10086 821
rect 10030 755 10034 815
rect 10115 805 10315 830
rect 10370 821 10400 1009
rect 10344 815 10400 821
rect 10086 755 10344 775
rect 10396 755 10400 815
rect 10030 745 10400 755
rect 10430 1075 10800 1085
rect 10430 1015 10434 1075
rect 10486 1055 10744 1075
rect 10430 1009 10486 1015
rect 10430 821 10460 1009
rect 10515 1000 10715 1025
rect 10796 1015 10800 1075
rect 10744 1009 10800 1015
rect 10515 980 10585 1000
rect 10490 940 10585 980
rect 10645 980 10715 1000
rect 10645 940 10740 980
rect 10490 890 10740 940
rect 10490 850 10585 890
rect 10515 830 10585 850
rect 10645 850 10740 890
rect 10645 830 10715 850
rect 10430 815 10486 821
rect 10430 755 10434 815
rect 10515 805 10715 830
rect 10770 821 10800 1009
rect 10744 815 10800 821
rect 10486 755 10744 775
rect 10796 755 10800 815
rect 10430 745 10800 755
rect 10830 1075 11200 1085
rect 10830 1015 10834 1075
rect 10886 1055 11144 1075
rect 10830 1009 10886 1015
rect 10830 821 10860 1009
rect 10915 1000 11115 1025
rect 11196 1015 11200 1075
rect 11144 1009 11200 1015
rect 10915 980 10985 1000
rect 10890 940 10985 980
rect 11045 980 11115 1000
rect 11045 940 11140 980
rect 10890 890 11140 940
rect 10890 850 10985 890
rect 10915 830 10985 850
rect 11045 850 11140 890
rect 11045 830 11115 850
rect 10830 815 10886 821
rect 10830 755 10834 815
rect 10915 805 11115 830
rect 11170 821 11200 1009
rect 11144 815 11200 821
rect 10886 755 11144 775
rect 11196 755 11200 815
rect 10830 745 11200 755
rect 11230 1075 11600 1085
rect 11230 1015 11234 1075
rect 11286 1055 11544 1075
rect 11230 1009 11286 1015
rect 11230 821 11260 1009
rect 11315 1000 11515 1025
rect 11596 1015 11600 1075
rect 11544 1009 11600 1015
rect 11315 980 11385 1000
rect 11290 940 11385 980
rect 11445 980 11515 1000
rect 11445 940 11540 980
rect 11290 890 11540 940
rect 11290 850 11385 890
rect 11315 830 11385 850
rect 11445 850 11540 890
rect 11445 830 11515 850
rect 11230 815 11286 821
rect 11230 755 11234 815
rect 11315 805 11515 830
rect 11570 821 11600 1009
rect 11544 815 11600 821
rect 11286 755 11544 775
rect 11596 755 11600 815
rect 11230 745 11600 755
rect 11630 1075 12000 1085
rect 11630 1015 11634 1075
rect 11686 1055 11944 1075
rect 11630 1009 11686 1015
rect 11630 821 11660 1009
rect 11715 1000 11915 1025
rect 11996 1015 12000 1075
rect 11944 1009 12000 1015
rect 11715 980 11785 1000
rect 11690 940 11785 980
rect 11845 980 11915 1000
rect 11845 940 11940 980
rect 11690 890 11940 940
rect 11690 850 11785 890
rect 11715 830 11785 850
rect 11845 850 11940 890
rect 11845 830 11915 850
rect 11630 815 11686 821
rect 11630 755 11634 815
rect 11715 805 11915 830
rect 11970 821 12000 1009
rect 11944 815 12000 821
rect 11686 755 11944 775
rect 11996 755 12000 815
rect 11630 745 12000 755
rect 12030 1075 12400 1085
rect 12030 1015 12034 1075
rect 12086 1055 12344 1075
rect 12030 1009 12086 1015
rect 12030 821 12060 1009
rect 12115 1000 12315 1025
rect 12396 1015 12400 1075
rect 12344 1009 12400 1015
rect 12115 980 12185 1000
rect 12090 940 12185 980
rect 12245 980 12315 1000
rect 12245 940 12340 980
rect 12090 890 12340 940
rect 12090 850 12185 890
rect 12115 830 12185 850
rect 12245 850 12340 890
rect 12245 830 12315 850
rect 12030 815 12086 821
rect 12030 755 12034 815
rect 12115 805 12315 830
rect 12370 821 12400 1009
rect 12344 815 12400 821
rect 12086 755 12344 775
rect 12396 755 12400 815
rect 12030 745 12400 755
rect 12430 1075 12800 1085
rect 12430 1015 12434 1075
rect 12486 1055 12744 1075
rect 12430 1009 12486 1015
rect 12430 821 12460 1009
rect 12515 1000 12715 1025
rect 12796 1015 12800 1075
rect 12744 1009 12800 1015
rect 12515 980 12585 1000
rect 12490 940 12585 980
rect 12645 980 12715 1000
rect 12645 940 12740 980
rect 12490 890 12740 940
rect 12490 850 12585 890
rect 12515 830 12585 850
rect 12645 850 12740 890
rect 12645 830 12715 850
rect 12430 815 12486 821
rect 12430 755 12434 815
rect 12515 805 12715 830
rect 12770 821 12800 1009
rect 12744 815 12800 821
rect 12486 755 12744 775
rect 12796 755 12800 815
rect 12430 745 12800 755
rect 12830 1075 13200 1085
rect 12830 1015 12834 1075
rect 12886 1055 13144 1075
rect 12830 1009 12886 1015
rect 12830 821 12860 1009
rect 12915 1000 13115 1025
rect 13196 1015 13200 1075
rect 13144 1009 13200 1015
rect 12915 980 12985 1000
rect 12890 940 12985 980
rect 13045 980 13115 1000
rect 13045 940 13140 980
rect 12890 890 13140 940
rect 12890 850 12985 890
rect 12915 830 12985 850
rect 13045 850 13140 890
rect 13045 830 13115 850
rect 12830 815 12886 821
rect 12830 755 12834 815
rect 12915 805 13115 830
rect 13170 821 13200 1009
rect 13144 815 13200 821
rect 12886 755 13144 775
rect 13196 755 13200 815
rect 12830 745 13200 755
rect -370 705 0 715
rect -370 645 -366 705
rect -314 685 -56 705
rect -370 639 -314 645
rect -370 451 -340 639
rect -285 630 -85 655
rect -4 645 0 705
rect -56 639 0 645
rect -285 610 -215 630
rect -310 570 -215 610
rect -155 610 -85 630
rect -155 570 -60 610
rect -310 520 -60 570
rect -310 480 -215 520
rect -285 460 -215 480
rect -155 480 -60 520
rect -155 460 -85 480
rect -370 445 -314 451
rect -370 385 -366 445
rect -285 435 -85 460
rect -30 451 0 639
rect -56 445 0 451
rect -314 385 -56 405
rect -4 385 0 445
rect -370 375 0 385
rect 30 705 400 715
rect 30 645 34 705
rect 86 685 344 705
rect 30 639 86 645
rect 30 451 60 639
rect 115 630 315 655
rect 396 645 400 705
rect 344 639 400 645
rect 115 610 185 630
rect 90 570 185 610
rect 245 610 315 630
rect 245 570 340 610
rect 90 520 340 570
rect 90 480 185 520
rect 115 460 185 480
rect 245 480 340 520
rect 245 460 315 480
rect 30 445 86 451
rect 30 385 34 445
rect 115 435 315 460
rect 370 451 400 639
rect 344 445 400 451
rect 86 385 344 405
rect 396 385 400 445
rect 30 375 400 385
rect 430 705 800 715
rect 430 645 434 705
rect 486 685 744 705
rect 430 639 486 645
rect 430 451 460 639
rect 515 630 715 655
rect 796 645 800 705
rect 744 639 800 645
rect 515 610 585 630
rect 490 570 585 610
rect 645 610 715 630
rect 645 570 740 610
rect 490 520 740 570
rect 490 480 585 520
rect 515 460 585 480
rect 645 480 740 520
rect 645 460 715 480
rect 430 445 486 451
rect 430 385 434 445
rect 515 435 715 460
rect 770 451 800 639
rect 744 445 800 451
rect 486 385 744 405
rect 796 385 800 445
rect 430 375 800 385
rect 830 705 1200 715
rect 830 645 834 705
rect 886 685 1144 705
rect 830 639 886 645
rect 830 451 860 639
rect 915 630 1115 655
rect 1196 645 1200 705
rect 1144 639 1200 645
rect 915 610 985 630
rect 890 570 985 610
rect 1045 610 1115 630
rect 1045 570 1140 610
rect 890 520 1140 570
rect 890 480 985 520
rect 915 460 985 480
rect 1045 480 1140 520
rect 1045 460 1115 480
rect 830 445 886 451
rect 830 385 834 445
rect 915 435 1115 460
rect 1170 451 1200 639
rect 1144 445 1200 451
rect 886 385 1144 405
rect 1196 385 1200 445
rect 830 375 1200 385
rect 1230 705 1600 715
rect 1230 645 1234 705
rect 1286 685 1544 705
rect 1230 639 1286 645
rect 1230 451 1260 639
rect 1315 630 1515 655
rect 1596 645 1600 705
rect 1544 639 1600 645
rect 1315 610 1385 630
rect 1290 570 1385 610
rect 1445 610 1515 630
rect 1445 570 1540 610
rect 1290 520 1540 570
rect 1290 480 1385 520
rect 1315 460 1385 480
rect 1445 480 1540 520
rect 1445 460 1515 480
rect 1230 445 1286 451
rect 1230 385 1234 445
rect 1315 435 1515 460
rect 1570 451 1600 639
rect 1544 445 1600 451
rect 1286 385 1544 405
rect 1596 385 1600 445
rect 1230 375 1600 385
rect 1630 705 2000 715
rect 1630 645 1634 705
rect 1686 685 1944 705
rect 1630 639 1686 645
rect 1630 451 1660 639
rect 1715 630 1915 655
rect 1996 645 2000 705
rect 1944 639 2000 645
rect 1715 610 1785 630
rect 1690 570 1785 610
rect 1845 610 1915 630
rect 1845 570 1940 610
rect 1690 520 1940 570
rect 1690 480 1785 520
rect 1715 460 1785 480
rect 1845 480 1940 520
rect 1845 460 1915 480
rect 1630 445 1686 451
rect 1630 385 1634 445
rect 1715 435 1915 460
rect 1970 451 2000 639
rect 1944 445 2000 451
rect 1686 385 1944 405
rect 1996 385 2000 445
rect 1630 375 2000 385
rect 2030 705 2400 715
rect 2030 645 2034 705
rect 2086 685 2344 705
rect 2030 639 2086 645
rect 2030 451 2060 639
rect 2115 630 2315 655
rect 2396 645 2400 705
rect 2344 639 2400 645
rect 2115 610 2185 630
rect 2090 570 2185 610
rect 2245 610 2315 630
rect 2245 570 2340 610
rect 2090 520 2340 570
rect 2090 480 2185 520
rect 2115 460 2185 480
rect 2245 480 2340 520
rect 2245 460 2315 480
rect 2030 445 2086 451
rect 2030 385 2034 445
rect 2115 435 2315 460
rect 2370 451 2400 639
rect 2344 445 2400 451
rect 2086 385 2344 405
rect 2396 385 2400 445
rect 2030 375 2400 385
rect 2430 705 2800 715
rect 2430 645 2434 705
rect 2486 685 2744 705
rect 2430 639 2486 645
rect 2430 451 2460 639
rect 2515 630 2715 655
rect 2796 645 2800 705
rect 2744 639 2800 645
rect 2515 610 2585 630
rect 2490 570 2585 610
rect 2645 610 2715 630
rect 2645 570 2740 610
rect 2490 520 2740 570
rect 2490 480 2585 520
rect 2515 460 2585 480
rect 2645 480 2740 520
rect 2645 460 2715 480
rect 2430 445 2486 451
rect 2430 385 2434 445
rect 2515 435 2715 460
rect 2770 451 2800 639
rect 2744 445 2800 451
rect 2486 385 2744 405
rect 2796 385 2800 445
rect 2430 375 2800 385
rect 2830 705 3200 715
rect 2830 645 2834 705
rect 2886 685 3144 705
rect 2830 639 2886 645
rect 2830 451 2860 639
rect 2915 630 3115 655
rect 3196 645 3200 705
rect 3144 639 3200 645
rect 2915 610 2985 630
rect 2890 570 2985 610
rect 3045 610 3115 630
rect 3045 570 3140 610
rect 2890 520 3140 570
rect 2890 480 2985 520
rect 2915 460 2985 480
rect 3045 480 3140 520
rect 3045 460 3115 480
rect 2830 445 2886 451
rect 2830 385 2834 445
rect 2915 435 3115 460
rect 3170 451 3200 639
rect 3144 445 3200 451
rect 2886 385 3144 405
rect 3196 385 3200 445
rect 2830 375 3200 385
rect 3230 705 3600 715
rect 3230 645 3234 705
rect 3286 685 3544 705
rect 3230 639 3286 645
rect 3230 451 3260 639
rect 3315 630 3515 655
rect 3596 645 3600 705
rect 3544 639 3600 645
rect 3315 610 3385 630
rect 3290 570 3385 610
rect 3445 610 3515 630
rect 3445 570 3540 610
rect 3290 520 3540 570
rect 3290 480 3385 520
rect 3315 460 3385 480
rect 3445 480 3540 520
rect 3445 460 3515 480
rect 3230 445 3286 451
rect 3230 385 3234 445
rect 3315 435 3515 460
rect 3570 451 3600 639
rect 3544 445 3600 451
rect 3286 385 3544 405
rect 3596 385 3600 445
rect 3230 375 3600 385
rect 3630 705 4000 715
rect 3630 645 3634 705
rect 3686 685 3944 705
rect 3630 639 3686 645
rect 3630 451 3660 639
rect 3715 630 3915 655
rect 3996 645 4000 705
rect 3944 639 4000 645
rect 3715 610 3785 630
rect 3690 570 3785 610
rect 3845 610 3915 630
rect 3845 570 3940 610
rect 3690 520 3940 570
rect 3690 480 3785 520
rect 3715 460 3785 480
rect 3845 480 3940 520
rect 3845 460 3915 480
rect 3630 445 3686 451
rect 3630 385 3634 445
rect 3715 435 3915 460
rect 3970 451 4000 639
rect 3944 445 4000 451
rect 3686 385 3944 405
rect 3996 385 4000 445
rect 3630 375 4000 385
rect 4030 705 4400 715
rect 4030 645 4034 705
rect 4086 685 4344 705
rect 4030 639 4086 645
rect 4030 451 4060 639
rect 4115 630 4315 655
rect 4396 645 4400 705
rect 4344 639 4400 645
rect 4115 610 4185 630
rect 4090 570 4185 610
rect 4245 610 4315 630
rect 4245 570 4340 610
rect 4090 520 4340 570
rect 4090 480 4185 520
rect 4115 460 4185 480
rect 4245 480 4340 520
rect 4245 460 4315 480
rect 4030 445 4086 451
rect 4030 385 4034 445
rect 4115 435 4315 460
rect 4370 451 4400 639
rect 4344 445 4400 451
rect 4086 385 4344 405
rect 4396 385 4400 445
rect 4030 375 4400 385
rect 4430 705 4800 715
rect 4430 645 4434 705
rect 4486 685 4744 705
rect 4430 639 4486 645
rect 4430 451 4460 639
rect 4515 630 4715 655
rect 4796 645 4800 705
rect 4744 639 4800 645
rect 4515 610 4585 630
rect 4490 570 4585 610
rect 4645 610 4715 630
rect 4645 570 4740 610
rect 4490 520 4740 570
rect 4490 480 4585 520
rect 4515 460 4585 480
rect 4645 480 4740 520
rect 4645 460 4715 480
rect 4430 445 4486 451
rect 4430 385 4434 445
rect 4515 435 4715 460
rect 4770 451 4800 639
rect 4744 445 4800 451
rect 4486 385 4744 405
rect 4796 385 4800 445
rect 4430 375 4800 385
rect 4830 705 5200 715
rect 4830 645 4834 705
rect 4886 685 5144 705
rect 4830 639 4886 645
rect 4830 451 4860 639
rect 4915 630 5115 655
rect 5196 645 5200 705
rect 5144 639 5200 645
rect 4915 610 4985 630
rect 4890 570 4985 610
rect 5045 610 5115 630
rect 5045 570 5140 610
rect 4890 520 5140 570
rect 4890 480 4985 520
rect 4915 460 4985 480
rect 5045 480 5140 520
rect 5045 460 5115 480
rect 4830 445 4886 451
rect 4830 385 4834 445
rect 4915 435 5115 460
rect 5170 451 5200 639
rect 5144 445 5200 451
rect 4886 385 5144 405
rect 5196 385 5200 445
rect 4830 375 5200 385
rect 5230 705 5600 715
rect 5230 645 5234 705
rect 5286 685 5544 705
rect 5230 639 5286 645
rect 5230 451 5260 639
rect 5315 630 5515 655
rect 5596 645 5600 705
rect 5544 639 5600 645
rect 5315 610 5385 630
rect 5290 570 5385 610
rect 5445 610 5515 630
rect 5445 570 5540 610
rect 5290 520 5540 570
rect 5290 480 5385 520
rect 5315 460 5385 480
rect 5445 480 5540 520
rect 5445 460 5515 480
rect 5230 445 5286 451
rect 5230 385 5234 445
rect 5315 435 5515 460
rect 5570 451 5600 639
rect 5544 445 5600 451
rect 5286 385 5544 405
rect 5596 385 5600 445
rect 5230 375 5600 385
rect 5630 705 6000 715
rect 5630 645 5634 705
rect 5686 685 5944 705
rect 5630 639 5686 645
rect 5630 451 5660 639
rect 5715 630 5915 655
rect 5996 645 6000 705
rect 5944 639 6000 645
rect 5715 610 5785 630
rect 5690 570 5785 610
rect 5845 610 5915 630
rect 5845 570 5940 610
rect 5690 520 5940 570
rect 5690 480 5785 520
rect 5715 460 5785 480
rect 5845 480 5940 520
rect 5845 460 5915 480
rect 5630 445 5686 451
rect 5630 385 5634 445
rect 5715 435 5915 460
rect 5970 451 6000 639
rect 5944 445 6000 451
rect 5686 385 5944 405
rect 5996 385 6000 445
rect 5630 375 6000 385
rect 6030 705 6400 715
rect 6030 645 6034 705
rect 6086 685 6344 705
rect 6030 639 6086 645
rect 6030 451 6060 639
rect 6115 630 6315 655
rect 6396 645 6400 705
rect 6344 639 6400 645
rect 6115 610 6185 630
rect 6090 570 6185 610
rect 6245 610 6315 630
rect 6245 570 6340 610
rect 6090 520 6340 570
rect 6090 480 6185 520
rect 6115 460 6185 480
rect 6245 480 6340 520
rect 6245 460 6315 480
rect 6030 445 6086 451
rect 6030 385 6034 445
rect 6115 435 6315 460
rect 6370 451 6400 639
rect 6344 445 6400 451
rect 6086 385 6344 405
rect 6396 385 6400 445
rect 6030 375 6400 385
rect 6430 705 6800 715
rect 6430 645 6434 705
rect 6486 685 6744 705
rect 6430 639 6486 645
rect 6430 451 6460 639
rect 6515 630 6715 655
rect 6796 645 6800 705
rect 6744 639 6800 645
rect 6515 610 6585 630
rect 6490 570 6585 610
rect 6645 610 6715 630
rect 6645 570 6740 610
rect 6490 520 6740 570
rect 6490 480 6585 520
rect 6515 460 6585 480
rect 6645 480 6740 520
rect 6645 460 6715 480
rect 6430 445 6486 451
rect 6430 385 6434 445
rect 6515 435 6715 460
rect 6770 451 6800 639
rect 6744 445 6800 451
rect 6486 385 6744 405
rect 6796 385 6800 445
rect 6430 375 6800 385
rect 6830 705 7200 715
rect 6830 645 6834 705
rect 6886 685 7144 705
rect 6830 639 6886 645
rect 6830 451 6860 639
rect 6915 630 7115 655
rect 7196 645 7200 705
rect 7144 639 7200 645
rect 6915 610 6985 630
rect 6890 570 6985 610
rect 7045 610 7115 630
rect 7045 570 7140 610
rect 6890 520 7140 570
rect 6890 480 6985 520
rect 6915 460 6985 480
rect 7045 480 7140 520
rect 7045 460 7115 480
rect 6830 445 6886 451
rect 6830 385 6834 445
rect 6915 435 7115 460
rect 7170 451 7200 639
rect 7144 445 7200 451
rect 6886 385 7144 405
rect 7196 385 7200 445
rect 6830 375 7200 385
rect 7230 705 7600 715
rect 7230 645 7234 705
rect 7286 685 7544 705
rect 7230 639 7286 645
rect 7230 451 7260 639
rect 7315 630 7515 655
rect 7596 645 7600 705
rect 7544 639 7600 645
rect 7315 610 7385 630
rect 7290 570 7385 610
rect 7445 610 7515 630
rect 7445 570 7540 610
rect 7290 520 7540 570
rect 7290 480 7385 520
rect 7315 460 7385 480
rect 7445 480 7540 520
rect 7445 460 7515 480
rect 7230 445 7286 451
rect 7230 385 7234 445
rect 7315 435 7515 460
rect 7570 451 7600 639
rect 7544 445 7600 451
rect 7286 385 7544 405
rect 7596 385 7600 445
rect 7230 375 7600 385
rect 7630 705 8000 715
rect 7630 645 7634 705
rect 7686 685 7944 705
rect 7630 639 7686 645
rect 7630 451 7660 639
rect 7715 630 7915 655
rect 7996 645 8000 705
rect 7944 639 8000 645
rect 7715 610 7785 630
rect 7690 570 7785 610
rect 7845 610 7915 630
rect 7845 570 7940 610
rect 7690 520 7940 570
rect 7690 480 7785 520
rect 7715 460 7785 480
rect 7845 480 7940 520
rect 7845 460 7915 480
rect 7630 445 7686 451
rect 7630 385 7634 445
rect 7715 435 7915 460
rect 7970 451 8000 639
rect 7944 445 8000 451
rect 7686 385 7944 405
rect 7996 385 8000 445
rect 7630 375 8000 385
rect 8030 705 8400 715
rect 8030 645 8034 705
rect 8086 685 8344 705
rect 8030 639 8086 645
rect 8030 451 8060 639
rect 8115 630 8315 655
rect 8396 645 8400 705
rect 8344 639 8400 645
rect 8115 610 8185 630
rect 8090 570 8185 610
rect 8245 610 8315 630
rect 8245 570 8340 610
rect 8090 520 8340 570
rect 8090 480 8185 520
rect 8115 460 8185 480
rect 8245 480 8340 520
rect 8245 460 8315 480
rect 8030 445 8086 451
rect 8030 385 8034 445
rect 8115 435 8315 460
rect 8370 451 8400 639
rect 8344 445 8400 451
rect 8086 385 8344 405
rect 8396 385 8400 445
rect 8030 375 8400 385
rect 8430 705 8800 715
rect 8430 645 8434 705
rect 8486 685 8744 705
rect 8430 639 8486 645
rect 8430 451 8460 639
rect 8515 630 8715 655
rect 8796 645 8800 705
rect 8744 639 8800 645
rect 8515 610 8585 630
rect 8490 570 8585 610
rect 8645 610 8715 630
rect 8645 570 8740 610
rect 8490 520 8740 570
rect 8490 480 8585 520
rect 8515 460 8585 480
rect 8645 480 8740 520
rect 8645 460 8715 480
rect 8430 445 8486 451
rect 8430 385 8434 445
rect 8515 435 8715 460
rect 8770 451 8800 639
rect 8744 445 8800 451
rect 8486 385 8744 405
rect 8796 385 8800 445
rect 8430 375 8800 385
rect 8830 705 9200 715
rect 8830 645 8834 705
rect 8886 685 9144 705
rect 8830 639 8886 645
rect 8830 451 8860 639
rect 8915 630 9115 655
rect 9196 645 9200 705
rect 9144 639 9200 645
rect 8915 610 8985 630
rect 8890 570 8985 610
rect 9045 610 9115 630
rect 9045 570 9140 610
rect 8890 520 9140 570
rect 8890 480 8985 520
rect 8915 460 8985 480
rect 9045 480 9140 520
rect 9045 460 9115 480
rect 8830 445 8886 451
rect 8830 385 8834 445
rect 8915 435 9115 460
rect 9170 451 9200 639
rect 9144 445 9200 451
rect 8886 385 9144 405
rect 9196 385 9200 445
rect 8830 375 9200 385
rect 9230 705 9600 715
rect 9230 645 9234 705
rect 9286 685 9544 705
rect 9230 639 9286 645
rect 9230 451 9260 639
rect 9315 630 9515 655
rect 9596 645 9600 705
rect 9544 639 9600 645
rect 9315 610 9385 630
rect 9290 570 9385 610
rect 9445 610 9515 630
rect 9445 570 9540 610
rect 9290 520 9540 570
rect 9290 480 9385 520
rect 9315 460 9385 480
rect 9445 480 9540 520
rect 9445 460 9515 480
rect 9230 445 9286 451
rect 9230 385 9234 445
rect 9315 435 9515 460
rect 9570 451 9600 639
rect 9544 445 9600 451
rect 9286 385 9544 405
rect 9596 385 9600 445
rect 9230 375 9600 385
rect 9630 705 10000 715
rect 9630 645 9634 705
rect 9686 685 9944 705
rect 9630 639 9686 645
rect 9630 451 9660 639
rect 9715 630 9915 655
rect 9996 645 10000 705
rect 9944 639 10000 645
rect 9715 610 9785 630
rect 9690 570 9785 610
rect 9845 610 9915 630
rect 9845 570 9940 610
rect 9690 520 9940 570
rect 9690 480 9785 520
rect 9715 460 9785 480
rect 9845 480 9940 520
rect 9845 460 9915 480
rect 9630 445 9686 451
rect 9630 385 9634 445
rect 9715 435 9915 460
rect 9970 451 10000 639
rect 9944 445 10000 451
rect 9686 385 9944 405
rect 9996 385 10000 445
rect 9630 375 10000 385
rect 10030 705 10400 715
rect 10030 645 10034 705
rect 10086 685 10344 705
rect 10030 639 10086 645
rect 10030 451 10060 639
rect 10115 630 10315 655
rect 10396 645 10400 705
rect 10344 639 10400 645
rect 10115 610 10185 630
rect 10090 570 10185 610
rect 10245 610 10315 630
rect 10245 570 10340 610
rect 10090 520 10340 570
rect 10090 480 10185 520
rect 10115 460 10185 480
rect 10245 480 10340 520
rect 10245 460 10315 480
rect 10030 445 10086 451
rect 10030 385 10034 445
rect 10115 435 10315 460
rect 10370 451 10400 639
rect 10344 445 10400 451
rect 10086 385 10344 405
rect 10396 385 10400 445
rect 10030 375 10400 385
rect 10430 705 10800 715
rect 10430 645 10434 705
rect 10486 685 10744 705
rect 10430 639 10486 645
rect 10430 451 10460 639
rect 10515 630 10715 655
rect 10796 645 10800 705
rect 10744 639 10800 645
rect 10515 610 10585 630
rect 10490 570 10585 610
rect 10645 610 10715 630
rect 10645 570 10740 610
rect 10490 520 10740 570
rect 10490 480 10585 520
rect 10515 460 10585 480
rect 10645 480 10740 520
rect 10645 460 10715 480
rect 10430 445 10486 451
rect 10430 385 10434 445
rect 10515 435 10715 460
rect 10770 451 10800 639
rect 10744 445 10800 451
rect 10486 385 10744 405
rect 10796 385 10800 445
rect 10430 375 10800 385
rect 10830 705 11200 715
rect 10830 645 10834 705
rect 10886 685 11144 705
rect 10830 639 10886 645
rect 10830 451 10860 639
rect 10915 630 11115 655
rect 11196 645 11200 705
rect 11144 639 11200 645
rect 10915 610 10985 630
rect 10890 570 10985 610
rect 11045 610 11115 630
rect 11045 570 11140 610
rect 10890 520 11140 570
rect 10890 480 10985 520
rect 10915 460 10985 480
rect 11045 480 11140 520
rect 11045 460 11115 480
rect 10830 445 10886 451
rect 10830 385 10834 445
rect 10915 435 11115 460
rect 11170 451 11200 639
rect 11144 445 11200 451
rect 10886 385 11144 405
rect 11196 385 11200 445
rect 10830 375 11200 385
rect 11230 705 11600 715
rect 11230 645 11234 705
rect 11286 685 11544 705
rect 11230 639 11286 645
rect 11230 451 11260 639
rect 11315 630 11515 655
rect 11596 645 11600 705
rect 11544 639 11600 645
rect 11315 610 11385 630
rect 11290 570 11385 610
rect 11445 610 11515 630
rect 11445 570 11540 610
rect 11290 520 11540 570
rect 11290 480 11385 520
rect 11315 460 11385 480
rect 11445 480 11540 520
rect 11445 460 11515 480
rect 11230 445 11286 451
rect 11230 385 11234 445
rect 11315 435 11515 460
rect 11570 451 11600 639
rect 11544 445 11600 451
rect 11286 385 11544 405
rect 11596 385 11600 445
rect 11230 375 11600 385
rect 11630 705 12000 715
rect 11630 645 11634 705
rect 11686 685 11944 705
rect 11630 639 11686 645
rect 11630 451 11660 639
rect 11715 630 11915 655
rect 11996 645 12000 705
rect 11944 639 12000 645
rect 11715 610 11785 630
rect 11690 570 11785 610
rect 11845 610 11915 630
rect 11845 570 11940 610
rect 11690 520 11940 570
rect 11690 480 11785 520
rect 11715 460 11785 480
rect 11845 480 11940 520
rect 11845 460 11915 480
rect 11630 445 11686 451
rect 11630 385 11634 445
rect 11715 435 11915 460
rect 11970 451 12000 639
rect 11944 445 12000 451
rect 11686 385 11944 405
rect 11996 385 12000 445
rect 11630 375 12000 385
rect 12030 705 12400 715
rect 12030 645 12034 705
rect 12086 685 12344 705
rect 12030 639 12086 645
rect 12030 451 12060 639
rect 12115 630 12315 655
rect 12396 645 12400 705
rect 12344 639 12400 645
rect 12115 610 12185 630
rect 12090 570 12185 610
rect 12245 610 12315 630
rect 12245 570 12340 610
rect 12090 520 12340 570
rect 12090 480 12185 520
rect 12115 460 12185 480
rect 12245 480 12340 520
rect 12245 460 12315 480
rect 12030 445 12086 451
rect 12030 385 12034 445
rect 12115 435 12315 460
rect 12370 451 12400 639
rect 12344 445 12400 451
rect 12086 385 12344 405
rect 12396 385 12400 445
rect 12030 375 12400 385
rect 12430 705 12800 715
rect 12430 645 12434 705
rect 12486 685 12744 705
rect 12430 639 12486 645
rect 12430 451 12460 639
rect 12515 630 12715 655
rect 12796 645 12800 705
rect 12744 639 12800 645
rect 12515 610 12585 630
rect 12490 570 12585 610
rect 12645 610 12715 630
rect 12645 570 12740 610
rect 12490 520 12740 570
rect 12490 480 12585 520
rect 12515 460 12585 480
rect 12645 480 12740 520
rect 12645 460 12715 480
rect 12430 445 12486 451
rect 12430 385 12434 445
rect 12515 435 12715 460
rect 12770 451 12800 639
rect 12744 445 12800 451
rect 12486 385 12744 405
rect 12796 385 12800 445
rect 12430 375 12800 385
rect 12830 705 13200 715
rect 12830 645 12834 705
rect 12886 685 13144 705
rect 12830 639 12886 645
rect 12830 451 12860 639
rect 12915 630 13115 655
rect 13196 645 13200 705
rect 13144 639 13200 645
rect 12915 610 12985 630
rect 12890 570 12985 610
rect 13045 610 13115 630
rect 13045 570 13140 610
rect 12890 520 13140 570
rect 12890 480 12985 520
rect 12915 460 12985 480
rect 13045 480 13140 520
rect 13045 460 13115 480
rect 12830 445 12886 451
rect 12830 385 12834 445
rect 12915 435 13115 460
rect 13170 451 13200 639
rect 13144 445 13200 451
rect 12886 385 13144 405
rect 13196 385 13200 445
rect 12830 375 13200 385
rect -370 335 0 345
rect -370 275 -366 335
rect -314 315 -56 335
rect -370 269 -314 275
rect -370 81 -340 269
rect -285 260 -85 285
rect -4 275 0 335
rect -56 269 0 275
rect -285 240 -215 260
rect -310 200 -215 240
rect -155 240 -85 260
rect -155 200 -60 240
rect -310 150 -60 200
rect -310 110 -215 150
rect -285 90 -215 110
rect -155 110 -60 150
rect -155 90 -85 110
rect -370 75 -314 81
rect -370 15 -366 75
rect -285 65 -85 90
rect -30 81 0 269
rect -56 75 0 81
rect -314 15 -56 35
rect -4 15 0 75
rect -370 5 0 15
rect 30 335 400 345
rect 30 275 34 335
rect 86 315 344 335
rect 30 269 86 275
rect 30 81 60 269
rect 115 260 315 285
rect 396 275 400 335
rect 344 269 400 275
rect 115 240 185 260
rect 90 200 185 240
rect 245 240 315 260
rect 245 200 340 240
rect 90 150 340 200
rect 90 110 185 150
rect 115 90 185 110
rect 245 110 340 150
rect 245 90 315 110
rect 30 75 86 81
rect 30 15 34 75
rect 115 65 315 90
rect 370 81 400 269
rect 344 75 400 81
rect 86 15 344 35
rect 396 15 400 75
rect 30 5 400 15
rect 430 335 800 345
rect 430 275 434 335
rect 486 315 744 335
rect 430 269 486 275
rect 430 81 460 269
rect 515 260 715 285
rect 796 275 800 335
rect 744 269 800 275
rect 515 240 585 260
rect 490 200 585 240
rect 645 240 715 260
rect 645 200 740 240
rect 490 150 740 200
rect 490 110 585 150
rect 515 90 585 110
rect 645 110 740 150
rect 645 90 715 110
rect 430 75 486 81
rect 430 15 434 75
rect 515 65 715 90
rect 770 81 800 269
rect 744 75 800 81
rect 486 15 744 35
rect 796 15 800 75
rect 430 5 800 15
rect 830 335 1200 345
rect 830 275 834 335
rect 886 315 1144 335
rect 830 269 886 275
rect 830 81 860 269
rect 915 260 1115 285
rect 1196 275 1200 335
rect 1144 269 1200 275
rect 915 240 985 260
rect 890 200 985 240
rect 1045 240 1115 260
rect 1045 200 1140 240
rect 890 150 1140 200
rect 890 110 985 150
rect 915 90 985 110
rect 1045 110 1140 150
rect 1045 90 1115 110
rect 830 75 886 81
rect 830 15 834 75
rect 915 65 1115 90
rect 1170 81 1200 269
rect 1144 75 1200 81
rect 886 15 1144 35
rect 1196 15 1200 75
rect 830 5 1200 15
rect 1230 335 1600 345
rect 1230 275 1234 335
rect 1286 315 1544 335
rect 1230 269 1286 275
rect 1230 81 1260 269
rect 1315 260 1515 285
rect 1596 275 1600 335
rect 1544 269 1600 275
rect 1315 240 1385 260
rect 1290 200 1385 240
rect 1445 240 1515 260
rect 1445 200 1540 240
rect 1290 150 1540 200
rect 1290 110 1385 150
rect 1315 90 1385 110
rect 1445 110 1540 150
rect 1445 90 1515 110
rect 1230 75 1286 81
rect 1230 15 1234 75
rect 1315 65 1515 90
rect 1570 81 1600 269
rect 1544 75 1600 81
rect 1286 15 1544 35
rect 1596 15 1600 75
rect 1230 5 1600 15
rect 1630 335 2000 345
rect 1630 275 1634 335
rect 1686 315 1944 335
rect 1630 269 1686 275
rect 1630 81 1660 269
rect 1715 260 1915 285
rect 1996 275 2000 335
rect 1944 269 2000 275
rect 1715 240 1785 260
rect 1690 200 1785 240
rect 1845 240 1915 260
rect 1845 200 1940 240
rect 1690 150 1940 200
rect 1690 110 1785 150
rect 1715 90 1785 110
rect 1845 110 1940 150
rect 1845 90 1915 110
rect 1630 75 1686 81
rect 1630 15 1634 75
rect 1715 65 1915 90
rect 1970 81 2000 269
rect 1944 75 2000 81
rect 1686 15 1944 35
rect 1996 15 2000 75
rect 1630 5 2000 15
rect 2030 335 2400 345
rect 2030 275 2034 335
rect 2086 315 2344 335
rect 2030 269 2086 275
rect 2030 81 2060 269
rect 2115 260 2315 285
rect 2396 275 2400 335
rect 2344 269 2400 275
rect 2115 240 2185 260
rect 2090 200 2185 240
rect 2245 240 2315 260
rect 2245 200 2340 240
rect 2090 150 2340 200
rect 2090 110 2185 150
rect 2115 90 2185 110
rect 2245 110 2340 150
rect 2245 90 2315 110
rect 2030 75 2086 81
rect 2030 15 2034 75
rect 2115 65 2315 90
rect 2370 81 2400 269
rect 2344 75 2400 81
rect 2086 15 2344 35
rect 2396 15 2400 75
rect 2030 5 2400 15
rect 2430 335 2800 345
rect 2430 275 2434 335
rect 2486 315 2744 335
rect 2430 269 2486 275
rect 2430 81 2460 269
rect 2515 260 2715 285
rect 2796 275 2800 335
rect 2744 269 2800 275
rect 2515 240 2585 260
rect 2490 200 2585 240
rect 2645 240 2715 260
rect 2645 200 2740 240
rect 2490 150 2740 200
rect 2490 110 2585 150
rect 2515 90 2585 110
rect 2645 110 2740 150
rect 2645 90 2715 110
rect 2430 75 2486 81
rect 2430 15 2434 75
rect 2515 65 2715 90
rect 2770 81 2800 269
rect 2744 75 2800 81
rect 2486 15 2744 35
rect 2796 15 2800 75
rect 2430 5 2800 15
rect 2830 335 3200 345
rect 2830 275 2834 335
rect 2886 315 3144 335
rect 2830 269 2886 275
rect 2830 81 2860 269
rect 2915 260 3115 285
rect 3196 275 3200 335
rect 3144 269 3200 275
rect 2915 240 2985 260
rect 2890 200 2985 240
rect 3045 240 3115 260
rect 3045 200 3140 240
rect 2890 150 3140 200
rect 2890 110 2985 150
rect 2915 90 2985 110
rect 3045 110 3140 150
rect 3045 90 3115 110
rect 2830 75 2886 81
rect 2830 15 2834 75
rect 2915 65 3115 90
rect 3170 81 3200 269
rect 3144 75 3200 81
rect 2886 15 3144 35
rect 3196 15 3200 75
rect 2830 5 3200 15
rect 3230 335 3600 345
rect 3230 275 3234 335
rect 3286 315 3544 335
rect 3230 269 3286 275
rect 3230 81 3260 269
rect 3315 260 3515 285
rect 3596 275 3600 335
rect 3544 269 3600 275
rect 3315 240 3385 260
rect 3290 200 3385 240
rect 3445 240 3515 260
rect 3445 200 3540 240
rect 3290 150 3540 200
rect 3290 110 3385 150
rect 3315 90 3385 110
rect 3445 110 3540 150
rect 3445 90 3515 110
rect 3230 75 3286 81
rect 3230 15 3234 75
rect 3315 65 3515 90
rect 3570 81 3600 269
rect 3544 75 3600 81
rect 3286 15 3544 35
rect 3596 15 3600 75
rect 3230 5 3600 15
rect 3630 335 4000 345
rect 3630 275 3634 335
rect 3686 315 3944 335
rect 3630 269 3686 275
rect 3630 81 3660 269
rect 3715 260 3915 285
rect 3996 275 4000 335
rect 3944 269 4000 275
rect 3715 240 3785 260
rect 3690 200 3785 240
rect 3845 240 3915 260
rect 3845 200 3940 240
rect 3690 150 3940 200
rect 3690 110 3785 150
rect 3715 90 3785 110
rect 3845 110 3940 150
rect 3845 90 3915 110
rect 3630 75 3686 81
rect 3630 15 3634 75
rect 3715 65 3915 90
rect 3970 81 4000 269
rect 3944 75 4000 81
rect 3686 15 3944 35
rect 3996 15 4000 75
rect 3630 5 4000 15
rect 4030 335 4400 345
rect 4030 275 4034 335
rect 4086 315 4344 335
rect 4030 269 4086 275
rect 4030 81 4060 269
rect 4115 260 4315 285
rect 4396 275 4400 335
rect 4344 269 4400 275
rect 4115 240 4185 260
rect 4090 200 4185 240
rect 4245 240 4315 260
rect 4245 200 4340 240
rect 4090 150 4340 200
rect 4090 110 4185 150
rect 4115 90 4185 110
rect 4245 110 4340 150
rect 4245 90 4315 110
rect 4030 75 4086 81
rect 4030 15 4034 75
rect 4115 65 4315 90
rect 4370 81 4400 269
rect 4344 75 4400 81
rect 4086 15 4344 35
rect 4396 15 4400 75
rect 4030 5 4400 15
rect 4430 335 4800 345
rect 4430 275 4434 335
rect 4486 315 4744 335
rect 4430 269 4486 275
rect 4430 81 4460 269
rect 4515 260 4715 285
rect 4796 275 4800 335
rect 4744 269 4800 275
rect 4515 240 4585 260
rect 4490 200 4585 240
rect 4645 240 4715 260
rect 4645 200 4740 240
rect 4490 150 4740 200
rect 4490 110 4585 150
rect 4515 90 4585 110
rect 4645 110 4740 150
rect 4645 90 4715 110
rect 4430 75 4486 81
rect 4430 15 4434 75
rect 4515 65 4715 90
rect 4770 81 4800 269
rect 4744 75 4800 81
rect 4486 15 4744 35
rect 4796 15 4800 75
rect 4430 5 4800 15
rect 4830 335 5200 345
rect 4830 275 4834 335
rect 4886 315 5144 335
rect 4830 269 4886 275
rect 4830 81 4860 269
rect 4915 260 5115 285
rect 5196 275 5200 335
rect 5144 269 5200 275
rect 4915 240 4985 260
rect 4890 200 4985 240
rect 5045 240 5115 260
rect 5045 200 5140 240
rect 4890 150 5140 200
rect 4890 110 4985 150
rect 4915 90 4985 110
rect 5045 110 5140 150
rect 5045 90 5115 110
rect 4830 75 4886 81
rect 4830 15 4834 75
rect 4915 65 5115 90
rect 5170 81 5200 269
rect 5144 75 5200 81
rect 4886 15 5144 35
rect 5196 15 5200 75
rect 4830 5 5200 15
rect 5230 335 5600 345
rect 5230 275 5234 335
rect 5286 315 5544 335
rect 5230 269 5286 275
rect 5230 81 5260 269
rect 5315 260 5515 285
rect 5596 275 5600 335
rect 5544 269 5600 275
rect 5315 240 5385 260
rect 5290 200 5385 240
rect 5445 240 5515 260
rect 5445 200 5540 240
rect 5290 150 5540 200
rect 5290 110 5385 150
rect 5315 90 5385 110
rect 5445 110 5540 150
rect 5445 90 5515 110
rect 5230 75 5286 81
rect 5230 15 5234 75
rect 5315 65 5515 90
rect 5570 81 5600 269
rect 5544 75 5600 81
rect 5286 15 5544 35
rect 5596 15 5600 75
rect 5230 5 5600 15
rect 5630 335 6000 345
rect 5630 275 5634 335
rect 5686 315 5944 335
rect 5630 269 5686 275
rect 5630 81 5660 269
rect 5715 260 5915 285
rect 5996 275 6000 335
rect 5944 269 6000 275
rect 5715 240 5785 260
rect 5690 200 5785 240
rect 5845 240 5915 260
rect 5845 200 5940 240
rect 5690 150 5940 200
rect 5690 110 5785 150
rect 5715 90 5785 110
rect 5845 110 5940 150
rect 5845 90 5915 110
rect 5630 75 5686 81
rect 5630 15 5634 75
rect 5715 65 5915 90
rect 5970 81 6000 269
rect 5944 75 6000 81
rect 5686 15 5944 35
rect 5996 15 6000 75
rect 5630 5 6000 15
rect 6030 335 6400 345
rect 6030 275 6034 335
rect 6086 315 6344 335
rect 6030 269 6086 275
rect 6030 81 6060 269
rect 6115 260 6315 285
rect 6396 275 6400 335
rect 6344 269 6400 275
rect 6115 240 6185 260
rect 6090 200 6185 240
rect 6245 240 6315 260
rect 6245 200 6340 240
rect 6090 150 6340 200
rect 6090 110 6185 150
rect 6115 90 6185 110
rect 6245 110 6340 150
rect 6245 90 6315 110
rect 6030 75 6086 81
rect 6030 15 6034 75
rect 6115 65 6315 90
rect 6370 81 6400 269
rect 6344 75 6400 81
rect 6086 15 6344 35
rect 6396 15 6400 75
rect 6030 5 6400 15
rect 6430 335 6800 345
rect 6430 275 6434 335
rect 6486 315 6744 335
rect 6430 269 6486 275
rect 6430 81 6460 269
rect 6515 260 6715 285
rect 6796 275 6800 335
rect 6744 269 6800 275
rect 6515 240 6585 260
rect 6490 200 6585 240
rect 6645 240 6715 260
rect 6645 200 6740 240
rect 6490 150 6740 200
rect 6490 110 6585 150
rect 6515 90 6585 110
rect 6645 110 6740 150
rect 6645 90 6715 110
rect 6430 75 6486 81
rect 6430 15 6434 75
rect 6515 65 6715 90
rect 6770 81 6800 269
rect 6744 75 6800 81
rect 6486 15 6744 35
rect 6796 15 6800 75
rect 6430 5 6800 15
rect 6830 335 7200 345
rect 6830 275 6834 335
rect 6886 315 7144 335
rect 6830 269 6886 275
rect 6830 81 6860 269
rect 6915 260 7115 285
rect 7196 275 7200 335
rect 7144 269 7200 275
rect 6915 240 6985 260
rect 6890 200 6985 240
rect 7045 240 7115 260
rect 7045 200 7140 240
rect 6890 150 7140 200
rect 6890 110 6985 150
rect 6915 90 6985 110
rect 7045 110 7140 150
rect 7045 90 7115 110
rect 6830 75 6886 81
rect 6830 15 6834 75
rect 6915 65 7115 90
rect 7170 81 7200 269
rect 7144 75 7200 81
rect 6886 15 7144 35
rect 7196 15 7200 75
rect 6830 5 7200 15
rect 7230 335 7600 345
rect 7230 275 7234 335
rect 7286 315 7544 335
rect 7230 269 7286 275
rect 7230 81 7260 269
rect 7315 260 7515 285
rect 7596 275 7600 335
rect 7544 269 7600 275
rect 7315 240 7385 260
rect 7290 200 7385 240
rect 7445 240 7515 260
rect 7445 200 7540 240
rect 7290 150 7540 200
rect 7290 110 7385 150
rect 7315 90 7385 110
rect 7445 110 7540 150
rect 7445 90 7515 110
rect 7230 75 7286 81
rect 7230 15 7234 75
rect 7315 65 7515 90
rect 7570 81 7600 269
rect 7544 75 7600 81
rect 7286 15 7544 35
rect 7596 15 7600 75
rect 7230 5 7600 15
rect 7630 335 8000 345
rect 7630 275 7634 335
rect 7686 315 7944 335
rect 7630 269 7686 275
rect 7630 81 7660 269
rect 7715 260 7915 285
rect 7996 275 8000 335
rect 7944 269 8000 275
rect 7715 240 7785 260
rect 7690 200 7785 240
rect 7845 240 7915 260
rect 7845 200 7940 240
rect 7690 150 7940 200
rect 7690 110 7785 150
rect 7715 90 7785 110
rect 7845 110 7940 150
rect 7845 90 7915 110
rect 7630 75 7686 81
rect 7630 15 7634 75
rect 7715 65 7915 90
rect 7970 81 8000 269
rect 7944 75 8000 81
rect 7686 15 7944 35
rect 7996 15 8000 75
rect 7630 5 8000 15
rect 8030 335 8400 345
rect 8030 275 8034 335
rect 8086 315 8344 335
rect 8030 269 8086 275
rect 8030 81 8060 269
rect 8115 260 8315 285
rect 8396 275 8400 335
rect 8344 269 8400 275
rect 8115 240 8185 260
rect 8090 200 8185 240
rect 8245 240 8315 260
rect 8245 200 8340 240
rect 8090 150 8340 200
rect 8090 110 8185 150
rect 8115 90 8185 110
rect 8245 110 8340 150
rect 8245 90 8315 110
rect 8030 75 8086 81
rect 8030 15 8034 75
rect 8115 65 8315 90
rect 8370 81 8400 269
rect 8344 75 8400 81
rect 8086 15 8344 35
rect 8396 15 8400 75
rect 8030 5 8400 15
rect 8430 335 8800 345
rect 8430 275 8434 335
rect 8486 315 8744 335
rect 8430 269 8486 275
rect 8430 81 8460 269
rect 8515 260 8715 285
rect 8796 275 8800 335
rect 8744 269 8800 275
rect 8515 240 8585 260
rect 8490 200 8585 240
rect 8645 240 8715 260
rect 8645 200 8740 240
rect 8490 150 8740 200
rect 8490 110 8585 150
rect 8515 90 8585 110
rect 8645 110 8740 150
rect 8645 90 8715 110
rect 8430 75 8486 81
rect 8430 15 8434 75
rect 8515 65 8715 90
rect 8770 81 8800 269
rect 8744 75 8800 81
rect 8486 15 8744 35
rect 8796 15 8800 75
rect 8430 5 8800 15
rect 8830 335 9200 345
rect 8830 275 8834 335
rect 8886 315 9144 335
rect 8830 269 8886 275
rect 8830 81 8860 269
rect 8915 260 9115 285
rect 9196 275 9200 335
rect 9144 269 9200 275
rect 8915 240 8985 260
rect 8890 200 8985 240
rect 9045 240 9115 260
rect 9045 200 9140 240
rect 8890 150 9140 200
rect 8890 110 8985 150
rect 8915 90 8985 110
rect 9045 110 9140 150
rect 9045 90 9115 110
rect 8830 75 8886 81
rect 8830 15 8834 75
rect 8915 65 9115 90
rect 9170 81 9200 269
rect 9144 75 9200 81
rect 8886 15 9144 35
rect 9196 15 9200 75
rect 8830 5 9200 15
rect 9230 335 9600 345
rect 9230 275 9234 335
rect 9286 315 9544 335
rect 9230 269 9286 275
rect 9230 81 9260 269
rect 9315 260 9515 285
rect 9596 275 9600 335
rect 9544 269 9600 275
rect 9315 240 9385 260
rect 9290 200 9385 240
rect 9445 240 9515 260
rect 9445 200 9540 240
rect 9290 150 9540 200
rect 9290 110 9385 150
rect 9315 90 9385 110
rect 9445 110 9540 150
rect 9445 90 9515 110
rect 9230 75 9286 81
rect 9230 15 9234 75
rect 9315 65 9515 90
rect 9570 81 9600 269
rect 9544 75 9600 81
rect 9286 15 9544 35
rect 9596 15 9600 75
rect 9230 5 9600 15
rect 9630 335 10000 345
rect 9630 275 9634 335
rect 9686 315 9944 335
rect 9630 269 9686 275
rect 9630 81 9660 269
rect 9715 260 9915 285
rect 9996 275 10000 335
rect 9944 269 10000 275
rect 9715 240 9785 260
rect 9690 200 9785 240
rect 9845 240 9915 260
rect 9845 200 9940 240
rect 9690 150 9940 200
rect 9690 110 9785 150
rect 9715 90 9785 110
rect 9845 110 9940 150
rect 9845 90 9915 110
rect 9630 75 9686 81
rect 9630 15 9634 75
rect 9715 65 9915 90
rect 9970 81 10000 269
rect 9944 75 10000 81
rect 9686 15 9944 35
rect 9996 15 10000 75
rect 9630 5 10000 15
rect 10030 335 10400 345
rect 10030 275 10034 335
rect 10086 315 10344 335
rect 10030 269 10086 275
rect 10030 81 10060 269
rect 10115 260 10315 285
rect 10396 275 10400 335
rect 10344 269 10400 275
rect 10115 240 10185 260
rect 10090 200 10185 240
rect 10245 240 10315 260
rect 10245 200 10340 240
rect 10090 150 10340 200
rect 10090 110 10185 150
rect 10115 90 10185 110
rect 10245 110 10340 150
rect 10245 90 10315 110
rect 10030 75 10086 81
rect 10030 15 10034 75
rect 10115 65 10315 90
rect 10370 81 10400 269
rect 10344 75 10400 81
rect 10086 15 10344 35
rect 10396 15 10400 75
rect 10030 5 10400 15
rect 10430 335 10800 345
rect 10430 275 10434 335
rect 10486 315 10744 335
rect 10430 269 10486 275
rect 10430 81 10460 269
rect 10515 260 10715 285
rect 10796 275 10800 335
rect 10744 269 10800 275
rect 10515 240 10585 260
rect 10490 200 10585 240
rect 10645 240 10715 260
rect 10645 200 10740 240
rect 10490 150 10740 200
rect 10490 110 10585 150
rect 10515 90 10585 110
rect 10645 110 10740 150
rect 10645 90 10715 110
rect 10430 75 10486 81
rect 10430 15 10434 75
rect 10515 65 10715 90
rect 10770 81 10800 269
rect 10744 75 10800 81
rect 10486 15 10744 35
rect 10796 15 10800 75
rect 10430 5 10800 15
rect 10830 335 11200 345
rect 10830 275 10834 335
rect 10886 315 11144 335
rect 10830 269 10886 275
rect 10830 81 10860 269
rect 10915 260 11115 285
rect 11196 275 11200 335
rect 11144 269 11200 275
rect 10915 240 10985 260
rect 10890 200 10985 240
rect 11045 240 11115 260
rect 11045 200 11140 240
rect 10890 150 11140 200
rect 10890 110 10985 150
rect 10915 90 10985 110
rect 11045 110 11140 150
rect 11045 90 11115 110
rect 10830 75 10886 81
rect 10830 15 10834 75
rect 10915 65 11115 90
rect 11170 81 11200 269
rect 11144 75 11200 81
rect 10886 15 11144 35
rect 11196 15 11200 75
rect 10830 5 11200 15
rect 11230 335 11600 345
rect 11230 275 11234 335
rect 11286 315 11544 335
rect 11230 269 11286 275
rect 11230 81 11260 269
rect 11315 260 11515 285
rect 11596 275 11600 335
rect 11544 269 11600 275
rect 11315 240 11385 260
rect 11290 200 11385 240
rect 11445 240 11515 260
rect 11445 200 11540 240
rect 11290 150 11540 200
rect 11290 110 11385 150
rect 11315 90 11385 110
rect 11445 110 11540 150
rect 11445 90 11515 110
rect 11230 75 11286 81
rect 11230 15 11234 75
rect 11315 65 11515 90
rect 11570 81 11600 269
rect 11544 75 11600 81
rect 11286 15 11544 35
rect 11596 15 11600 75
rect 11230 5 11600 15
rect 11630 335 12000 345
rect 11630 275 11634 335
rect 11686 315 11944 335
rect 11630 269 11686 275
rect 11630 81 11660 269
rect 11715 260 11915 285
rect 11996 275 12000 335
rect 11944 269 12000 275
rect 11715 240 11785 260
rect 11690 200 11785 240
rect 11845 240 11915 260
rect 11845 200 11940 240
rect 11690 150 11940 200
rect 11690 110 11785 150
rect 11715 90 11785 110
rect 11845 110 11940 150
rect 11845 90 11915 110
rect 11630 75 11686 81
rect 11630 15 11634 75
rect 11715 65 11915 90
rect 11970 81 12000 269
rect 11944 75 12000 81
rect 11686 15 11944 35
rect 11996 15 12000 75
rect 11630 5 12000 15
rect 12030 335 12400 345
rect 12030 275 12034 335
rect 12086 315 12344 335
rect 12030 269 12086 275
rect 12030 81 12060 269
rect 12115 260 12315 285
rect 12396 275 12400 335
rect 12344 269 12400 275
rect 12115 240 12185 260
rect 12090 200 12185 240
rect 12245 240 12315 260
rect 12245 200 12340 240
rect 12090 150 12340 200
rect 12090 110 12185 150
rect 12115 90 12185 110
rect 12245 110 12340 150
rect 12245 90 12315 110
rect 12030 75 12086 81
rect 12030 15 12034 75
rect 12115 65 12315 90
rect 12370 81 12400 269
rect 12344 75 12400 81
rect 12086 15 12344 35
rect 12396 15 12400 75
rect 12030 5 12400 15
rect 12430 335 12800 345
rect 12430 275 12434 335
rect 12486 315 12744 335
rect 12430 269 12486 275
rect 12430 81 12460 269
rect 12515 260 12715 285
rect 12796 275 12800 335
rect 12744 269 12800 275
rect 12515 240 12585 260
rect 12490 200 12585 240
rect 12645 240 12715 260
rect 12645 200 12740 240
rect 12490 150 12740 200
rect 12490 110 12585 150
rect 12515 90 12585 110
rect 12645 110 12740 150
rect 12645 90 12715 110
rect 12430 75 12486 81
rect 12430 15 12434 75
rect 12515 65 12715 90
rect 12770 81 12800 269
rect 12744 75 12800 81
rect 12486 15 12744 35
rect 12796 15 12800 75
rect 12430 5 12800 15
rect 12830 335 13200 345
rect 12830 275 12834 335
rect 12886 315 13144 335
rect 12830 269 12886 275
rect 12830 81 12860 269
rect 12915 260 13115 285
rect 13196 275 13200 335
rect 13144 269 13200 275
rect 12915 240 12985 260
rect 12890 200 12985 240
rect 13045 240 13115 260
rect 13045 200 13140 240
rect 12890 150 13140 200
rect 12890 110 12985 150
rect 12915 90 12985 110
rect 13045 110 13140 150
rect 13045 90 13115 110
rect 12830 75 12886 81
rect 12830 15 12834 75
rect 12915 65 13115 90
rect 13170 81 13200 269
rect 13144 75 13200 81
rect 12886 15 13144 35
rect 13196 15 13200 75
rect 12830 5 13200 15
rect -370 -35 0 -25
rect -370 -95 -366 -35
rect -314 -55 -56 -35
rect -370 -101 -314 -95
rect -370 -289 -340 -101
rect -285 -110 -85 -85
rect -4 -95 0 -35
rect -56 -101 0 -95
rect -285 -130 -215 -110
rect -310 -170 -215 -130
rect -155 -130 -85 -110
rect -155 -170 -60 -130
rect -310 -220 -60 -170
rect -310 -260 -215 -220
rect -285 -280 -215 -260
rect -155 -260 -60 -220
rect -155 -280 -85 -260
rect -370 -295 -314 -289
rect -370 -355 -366 -295
rect -285 -305 -85 -280
rect -30 -289 0 -101
rect -56 -295 0 -289
rect -314 -355 -56 -335
rect -4 -355 0 -295
rect -370 -365 0 -355
rect 30 -35 400 -25
rect 30 -95 34 -35
rect 86 -55 344 -35
rect 30 -101 86 -95
rect 30 -289 60 -101
rect 115 -110 315 -85
rect 396 -95 400 -35
rect 344 -101 400 -95
rect 115 -130 185 -110
rect 90 -170 185 -130
rect 245 -130 315 -110
rect 245 -170 340 -130
rect 90 -220 340 -170
rect 90 -260 185 -220
rect 115 -280 185 -260
rect 245 -260 340 -220
rect 245 -280 315 -260
rect 30 -295 86 -289
rect 30 -355 34 -295
rect 115 -305 315 -280
rect 370 -289 400 -101
rect 344 -295 400 -289
rect 86 -355 344 -335
rect 396 -355 400 -295
rect 30 -365 400 -355
rect 430 -35 800 -25
rect 430 -95 434 -35
rect 486 -55 744 -35
rect 430 -101 486 -95
rect 430 -289 460 -101
rect 515 -110 715 -85
rect 796 -95 800 -35
rect 744 -101 800 -95
rect 515 -130 585 -110
rect 490 -170 585 -130
rect 645 -130 715 -110
rect 645 -170 740 -130
rect 490 -220 740 -170
rect 490 -260 585 -220
rect 515 -280 585 -260
rect 645 -260 740 -220
rect 645 -280 715 -260
rect 430 -295 486 -289
rect 430 -355 434 -295
rect 515 -305 715 -280
rect 770 -289 800 -101
rect 744 -295 800 -289
rect 486 -355 744 -335
rect 796 -355 800 -295
rect 430 -365 800 -355
rect 830 -35 1200 -25
rect 830 -95 834 -35
rect 886 -55 1144 -35
rect 830 -101 886 -95
rect 830 -289 860 -101
rect 915 -110 1115 -85
rect 1196 -95 1200 -35
rect 1144 -101 1200 -95
rect 915 -130 985 -110
rect 890 -170 985 -130
rect 1045 -130 1115 -110
rect 1045 -170 1140 -130
rect 890 -220 1140 -170
rect 890 -260 985 -220
rect 915 -280 985 -260
rect 1045 -260 1140 -220
rect 1045 -280 1115 -260
rect 830 -295 886 -289
rect 830 -355 834 -295
rect 915 -305 1115 -280
rect 1170 -289 1200 -101
rect 1144 -295 1200 -289
rect 886 -355 1144 -335
rect 1196 -355 1200 -295
rect 830 -365 1200 -355
rect 1230 -35 1600 -25
rect 1230 -95 1234 -35
rect 1286 -55 1544 -35
rect 1230 -101 1286 -95
rect 1230 -289 1260 -101
rect 1315 -110 1515 -85
rect 1596 -95 1600 -35
rect 1544 -101 1600 -95
rect 1315 -130 1385 -110
rect 1290 -170 1385 -130
rect 1445 -130 1515 -110
rect 1445 -170 1540 -130
rect 1290 -220 1540 -170
rect 1290 -260 1385 -220
rect 1315 -280 1385 -260
rect 1445 -260 1540 -220
rect 1445 -280 1515 -260
rect 1230 -295 1286 -289
rect 1230 -355 1234 -295
rect 1315 -305 1515 -280
rect 1570 -289 1600 -101
rect 1544 -295 1600 -289
rect 1286 -355 1544 -335
rect 1596 -355 1600 -295
rect 1230 -365 1600 -355
rect 1630 -35 2000 -25
rect 1630 -95 1634 -35
rect 1686 -55 1944 -35
rect 1630 -101 1686 -95
rect 1630 -289 1660 -101
rect 1715 -110 1915 -85
rect 1996 -95 2000 -35
rect 1944 -101 2000 -95
rect 1715 -130 1785 -110
rect 1690 -170 1785 -130
rect 1845 -130 1915 -110
rect 1845 -170 1940 -130
rect 1690 -220 1940 -170
rect 1690 -260 1785 -220
rect 1715 -280 1785 -260
rect 1845 -260 1940 -220
rect 1845 -280 1915 -260
rect 1630 -295 1686 -289
rect 1630 -355 1634 -295
rect 1715 -305 1915 -280
rect 1970 -289 2000 -101
rect 1944 -295 2000 -289
rect 1686 -355 1944 -335
rect 1996 -355 2000 -295
rect 1630 -365 2000 -355
rect 2030 -35 2400 -25
rect 2030 -95 2034 -35
rect 2086 -55 2344 -35
rect 2030 -101 2086 -95
rect 2030 -289 2060 -101
rect 2115 -110 2315 -85
rect 2396 -95 2400 -35
rect 2344 -101 2400 -95
rect 2115 -130 2185 -110
rect 2090 -170 2185 -130
rect 2245 -130 2315 -110
rect 2245 -170 2340 -130
rect 2090 -220 2340 -170
rect 2090 -260 2185 -220
rect 2115 -280 2185 -260
rect 2245 -260 2340 -220
rect 2245 -280 2315 -260
rect 2030 -295 2086 -289
rect 2030 -355 2034 -295
rect 2115 -305 2315 -280
rect 2370 -289 2400 -101
rect 2344 -295 2400 -289
rect 2086 -355 2344 -335
rect 2396 -355 2400 -295
rect 2030 -365 2400 -355
rect 2430 -35 2800 -25
rect 2430 -95 2434 -35
rect 2486 -55 2744 -35
rect 2430 -101 2486 -95
rect 2430 -289 2460 -101
rect 2515 -110 2715 -85
rect 2796 -95 2800 -35
rect 2744 -101 2800 -95
rect 2515 -130 2585 -110
rect 2490 -170 2585 -130
rect 2645 -130 2715 -110
rect 2645 -170 2740 -130
rect 2490 -220 2740 -170
rect 2490 -260 2585 -220
rect 2515 -280 2585 -260
rect 2645 -260 2740 -220
rect 2645 -280 2715 -260
rect 2430 -295 2486 -289
rect 2430 -355 2434 -295
rect 2515 -305 2715 -280
rect 2770 -289 2800 -101
rect 2744 -295 2800 -289
rect 2486 -355 2744 -335
rect 2796 -355 2800 -295
rect 2430 -365 2800 -355
rect 2830 -35 3200 -25
rect 2830 -95 2834 -35
rect 2886 -55 3144 -35
rect 2830 -101 2886 -95
rect 2830 -289 2860 -101
rect 2915 -110 3115 -85
rect 3196 -95 3200 -35
rect 3144 -101 3200 -95
rect 2915 -130 2985 -110
rect 2890 -170 2985 -130
rect 3045 -130 3115 -110
rect 3045 -170 3140 -130
rect 2890 -220 3140 -170
rect 2890 -260 2985 -220
rect 2915 -280 2985 -260
rect 3045 -260 3140 -220
rect 3045 -280 3115 -260
rect 2830 -295 2886 -289
rect 2830 -355 2834 -295
rect 2915 -305 3115 -280
rect 3170 -289 3200 -101
rect 3144 -295 3200 -289
rect 2886 -355 3144 -335
rect 3196 -355 3200 -295
rect 2830 -365 3200 -355
rect 3230 -35 3600 -25
rect 3230 -95 3234 -35
rect 3286 -55 3544 -35
rect 3230 -101 3286 -95
rect 3230 -289 3260 -101
rect 3315 -110 3515 -85
rect 3596 -95 3600 -35
rect 3544 -101 3600 -95
rect 3315 -130 3385 -110
rect 3290 -170 3385 -130
rect 3445 -130 3515 -110
rect 3445 -170 3540 -130
rect 3290 -220 3540 -170
rect 3290 -260 3385 -220
rect 3315 -280 3385 -260
rect 3445 -260 3540 -220
rect 3445 -280 3515 -260
rect 3230 -295 3286 -289
rect 3230 -355 3234 -295
rect 3315 -305 3515 -280
rect 3570 -289 3600 -101
rect 3544 -295 3600 -289
rect 3286 -355 3544 -335
rect 3596 -355 3600 -295
rect 3230 -365 3600 -355
rect 3630 -35 4000 -25
rect 3630 -95 3634 -35
rect 3686 -55 3944 -35
rect 3630 -101 3686 -95
rect 3630 -289 3660 -101
rect 3715 -110 3915 -85
rect 3996 -95 4000 -35
rect 3944 -101 4000 -95
rect 3715 -130 3785 -110
rect 3690 -170 3785 -130
rect 3845 -130 3915 -110
rect 3845 -170 3940 -130
rect 3690 -220 3940 -170
rect 3690 -260 3785 -220
rect 3715 -280 3785 -260
rect 3845 -260 3940 -220
rect 3845 -280 3915 -260
rect 3630 -295 3686 -289
rect 3630 -355 3634 -295
rect 3715 -305 3915 -280
rect 3970 -289 4000 -101
rect 3944 -295 4000 -289
rect 3686 -355 3944 -335
rect 3996 -355 4000 -295
rect 3630 -365 4000 -355
rect 4030 -35 4400 -25
rect 4030 -95 4034 -35
rect 4086 -55 4344 -35
rect 4030 -101 4086 -95
rect 4030 -289 4060 -101
rect 4115 -110 4315 -85
rect 4396 -95 4400 -35
rect 4344 -101 4400 -95
rect 4115 -130 4185 -110
rect 4090 -170 4185 -130
rect 4245 -130 4315 -110
rect 4245 -170 4340 -130
rect 4090 -220 4340 -170
rect 4090 -260 4185 -220
rect 4115 -280 4185 -260
rect 4245 -260 4340 -220
rect 4245 -280 4315 -260
rect 4030 -295 4086 -289
rect 4030 -355 4034 -295
rect 4115 -305 4315 -280
rect 4370 -289 4400 -101
rect 4344 -295 4400 -289
rect 4086 -355 4344 -335
rect 4396 -355 4400 -295
rect 4030 -365 4400 -355
rect 4430 -35 4800 -25
rect 4430 -95 4434 -35
rect 4486 -55 4744 -35
rect 4430 -101 4486 -95
rect 4430 -289 4460 -101
rect 4515 -110 4715 -85
rect 4796 -95 4800 -35
rect 4744 -101 4800 -95
rect 4515 -130 4585 -110
rect 4490 -170 4585 -130
rect 4645 -130 4715 -110
rect 4645 -170 4740 -130
rect 4490 -220 4740 -170
rect 4490 -260 4585 -220
rect 4515 -280 4585 -260
rect 4645 -260 4740 -220
rect 4645 -280 4715 -260
rect 4430 -295 4486 -289
rect 4430 -355 4434 -295
rect 4515 -305 4715 -280
rect 4770 -289 4800 -101
rect 4744 -295 4800 -289
rect 4486 -355 4744 -335
rect 4796 -355 4800 -295
rect 4430 -365 4800 -355
rect 4830 -35 5200 -25
rect 4830 -95 4834 -35
rect 4886 -55 5144 -35
rect 4830 -101 4886 -95
rect 4830 -289 4860 -101
rect 4915 -110 5115 -85
rect 5196 -95 5200 -35
rect 5144 -101 5200 -95
rect 4915 -130 4985 -110
rect 4890 -170 4985 -130
rect 5045 -130 5115 -110
rect 5045 -170 5140 -130
rect 4890 -220 5140 -170
rect 4890 -260 4985 -220
rect 4915 -280 4985 -260
rect 5045 -260 5140 -220
rect 5045 -280 5115 -260
rect 4830 -295 4886 -289
rect 4830 -355 4834 -295
rect 4915 -305 5115 -280
rect 5170 -289 5200 -101
rect 5144 -295 5200 -289
rect 4886 -355 5144 -335
rect 5196 -355 5200 -295
rect 4830 -365 5200 -355
rect 5230 -35 5600 -25
rect 5230 -95 5234 -35
rect 5286 -55 5544 -35
rect 5230 -101 5286 -95
rect 5230 -289 5260 -101
rect 5315 -110 5515 -85
rect 5596 -95 5600 -35
rect 5544 -101 5600 -95
rect 5315 -130 5385 -110
rect 5290 -170 5385 -130
rect 5445 -130 5515 -110
rect 5445 -170 5540 -130
rect 5290 -220 5540 -170
rect 5290 -260 5385 -220
rect 5315 -280 5385 -260
rect 5445 -260 5540 -220
rect 5445 -280 5515 -260
rect 5230 -295 5286 -289
rect 5230 -355 5234 -295
rect 5315 -305 5515 -280
rect 5570 -289 5600 -101
rect 5544 -295 5600 -289
rect 5286 -355 5544 -335
rect 5596 -355 5600 -295
rect 5230 -365 5600 -355
rect 5630 -35 6000 -25
rect 5630 -95 5634 -35
rect 5686 -55 5944 -35
rect 5630 -101 5686 -95
rect 5630 -289 5660 -101
rect 5715 -110 5915 -85
rect 5996 -95 6000 -35
rect 5944 -101 6000 -95
rect 5715 -130 5785 -110
rect 5690 -170 5785 -130
rect 5845 -130 5915 -110
rect 5845 -170 5940 -130
rect 5690 -220 5940 -170
rect 5690 -260 5785 -220
rect 5715 -280 5785 -260
rect 5845 -260 5940 -220
rect 5845 -280 5915 -260
rect 5630 -295 5686 -289
rect 5630 -355 5634 -295
rect 5715 -305 5915 -280
rect 5970 -289 6000 -101
rect 5944 -295 6000 -289
rect 5686 -355 5944 -335
rect 5996 -355 6000 -295
rect 5630 -365 6000 -355
rect 6030 -35 6400 -25
rect 6030 -95 6034 -35
rect 6086 -55 6344 -35
rect 6030 -101 6086 -95
rect 6030 -289 6060 -101
rect 6115 -110 6315 -85
rect 6396 -95 6400 -35
rect 6344 -101 6400 -95
rect 6115 -130 6185 -110
rect 6090 -170 6185 -130
rect 6245 -130 6315 -110
rect 6245 -170 6340 -130
rect 6090 -220 6340 -170
rect 6090 -260 6185 -220
rect 6115 -280 6185 -260
rect 6245 -260 6340 -220
rect 6245 -280 6315 -260
rect 6030 -295 6086 -289
rect 6030 -355 6034 -295
rect 6115 -305 6315 -280
rect 6370 -289 6400 -101
rect 6344 -295 6400 -289
rect 6086 -355 6344 -335
rect 6396 -355 6400 -295
rect 6030 -365 6400 -355
rect 6430 -35 6800 -25
rect 6430 -95 6434 -35
rect 6486 -55 6744 -35
rect 6430 -101 6486 -95
rect 6430 -289 6460 -101
rect 6515 -110 6715 -85
rect 6796 -95 6800 -35
rect 6744 -101 6800 -95
rect 6515 -130 6585 -110
rect 6490 -170 6585 -130
rect 6645 -130 6715 -110
rect 6645 -170 6740 -130
rect 6490 -220 6740 -170
rect 6490 -260 6585 -220
rect 6515 -280 6585 -260
rect 6645 -260 6740 -220
rect 6645 -280 6715 -260
rect 6430 -295 6486 -289
rect 6430 -355 6434 -295
rect 6515 -305 6715 -280
rect 6770 -289 6800 -101
rect 6744 -295 6800 -289
rect 6486 -355 6744 -335
rect 6796 -355 6800 -295
rect 6430 -365 6800 -355
rect 6830 -35 7200 -25
rect 6830 -95 6834 -35
rect 6886 -55 7144 -35
rect 6830 -101 6886 -95
rect 6830 -289 6860 -101
rect 6915 -110 7115 -85
rect 7196 -95 7200 -35
rect 7144 -101 7200 -95
rect 6915 -130 6985 -110
rect 6890 -170 6985 -130
rect 7045 -130 7115 -110
rect 7045 -170 7140 -130
rect 6890 -220 7140 -170
rect 6890 -260 6985 -220
rect 6915 -280 6985 -260
rect 7045 -260 7140 -220
rect 7045 -280 7115 -260
rect 6830 -295 6886 -289
rect 6830 -355 6834 -295
rect 6915 -305 7115 -280
rect 7170 -289 7200 -101
rect 7144 -295 7200 -289
rect 6886 -355 7144 -335
rect 7196 -355 7200 -295
rect 6830 -365 7200 -355
rect 7230 -35 7600 -25
rect 7230 -95 7234 -35
rect 7286 -55 7544 -35
rect 7230 -101 7286 -95
rect 7230 -289 7260 -101
rect 7315 -110 7515 -85
rect 7596 -95 7600 -35
rect 7544 -101 7600 -95
rect 7315 -130 7385 -110
rect 7290 -170 7385 -130
rect 7445 -130 7515 -110
rect 7445 -170 7540 -130
rect 7290 -220 7540 -170
rect 7290 -260 7385 -220
rect 7315 -280 7385 -260
rect 7445 -260 7540 -220
rect 7445 -280 7515 -260
rect 7230 -295 7286 -289
rect 7230 -355 7234 -295
rect 7315 -305 7515 -280
rect 7570 -289 7600 -101
rect 7544 -295 7600 -289
rect 7286 -355 7544 -335
rect 7596 -355 7600 -295
rect 7230 -365 7600 -355
rect 7630 -35 8000 -25
rect 7630 -95 7634 -35
rect 7686 -55 7944 -35
rect 7630 -101 7686 -95
rect 7630 -289 7660 -101
rect 7715 -110 7915 -85
rect 7996 -95 8000 -35
rect 7944 -101 8000 -95
rect 7715 -130 7785 -110
rect 7690 -170 7785 -130
rect 7845 -130 7915 -110
rect 7845 -170 7940 -130
rect 7690 -220 7940 -170
rect 7690 -260 7785 -220
rect 7715 -280 7785 -260
rect 7845 -260 7940 -220
rect 7845 -280 7915 -260
rect 7630 -295 7686 -289
rect 7630 -355 7634 -295
rect 7715 -305 7915 -280
rect 7970 -289 8000 -101
rect 7944 -295 8000 -289
rect 7686 -355 7944 -335
rect 7996 -355 8000 -295
rect 7630 -365 8000 -355
rect 8030 -35 8400 -25
rect 8030 -95 8034 -35
rect 8086 -55 8344 -35
rect 8030 -101 8086 -95
rect 8030 -289 8060 -101
rect 8115 -110 8315 -85
rect 8396 -95 8400 -35
rect 8344 -101 8400 -95
rect 8115 -130 8185 -110
rect 8090 -170 8185 -130
rect 8245 -130 8315 -110
rect 8245 -170 8340 -130
rect 8090 -220 8340 -170
rect 8090 -260 8185 -220
rect 8115 -280 8185 -260
rect 8245 -260 8340 -220
rect 8245 -280 8315 -260
rect 8030 -295 8086 -289
rect 8030 -355 8034 -295
rect 8115 -305 8315 -280
rect 8370 -289 8400 -101
rect 8344 -295 8400 -289
rect 8086 -355 8344 -335
rect 8396 -355 8400 -295
rect 8030 -365 8400 -355
rect 8430 -35 8800 -25
rect 8430 -95 8434 -35
rect 8486 -55 8744 -35
rect 8430 -101 8486 -95
rect 8430 -289 8460 -101
rect 8515 -110 8715 -85
rect 8796 -95 8800 -35
rect 8744 -101 8800 -95
rect 8515 -130 8585 -110
rect 8490 -170 8585 -130
rect 8645 -130 8715 -110
rect 8645 -170 8740 -130
rect 8490 -220 8740 -170
rect 8490 -260 8585 -220
rect 8515 -280 8585 -260
rect 8645 -260 8740 -220
rect 8645 -280 8715 -260
rect 8430 -295 8486 -289
rect 8430 -355 8434 -295
rect 8515 -305 8715 -280
rect 8770 -289 8800 -101
rect 8744 -295 8800 -289
rect 8486 -355 8744 -335
rect 8796 -355 8800 -295
rect 8430 -365 8800 -355
rect 8830 -35 9200 -25
rect 8830 -95 8834 -35
rect 8886 -55 9144 -35
rect 8830 -101 8886 -95
rect 8830 -289 8860 -101
rect 8915 -110 9115 -85
rect 9196 -95 9200 -35
rect 9144 -101 9200 -95
rect 8915 -130 8985 -110
rect 8890 -170 8985 -130
rect 9045 -130 9115 -110
rect 9045 -170 9140 -130
rect 8890 -220 9140 -170
rect 8890 -260 8985 -220
rect 8915 -280 8985 -260
rect 9045 -260 9140 -220
rect 9045 -280 9115 -260
rect 8830 -295 8886 -289
rect 8830 -355 8834 -295
rect 8915 -305 9115 -280
rect 9170 -289 9200 -101
rect 9144 -295 9200 -289
rect 8886 -355 9144 -335
rect 9196 -355 9200 -295
rect 8830 -365 9200 -355
rect 9230 -35 9600 -25
rect 9230 -95 9234 -35
rect 9286 -55 9544 -35
rect 9230 -101 9286 -95
rect 9230 -289 9260 -101
rect 9315 -110 9515 -85
rect 9596 -95 9600 -35
rect 9544 -101 9600 -95
rect 9315 -130 9385 -110
rect 9290 -170 9385 -130
rect 9445 -130 9515 -110
rect 9445 -170 9540 -130
rect 9290 -220 9540 -170
rect 9290 -260 9385 -220
rect 9315 -280 9385 -260
rect 9445 -260 9540 -220
rect 9445 -280 9515 -260
rect 9230 -295 9286 -289
rect 9230 -355 9234 -295
rect 9315 -305 9515 -280
rect 9570 -289 9600 -101
rect 9544 -295 9600 -289
rect 9286 -355 9544 -335
rect 9596 -355 9600 -295
rect 9230 -365 9600 -355
rect 9630 -35 10000 -25
rect 9630 -95 9634 -35
rect 9686 -55 9944 -35
rect 9630 -101 9686 -95
rect 9630 -289 9660 -101
rect 9715 -110 9915 -85
rect 9996 -95 10000 -35
rect 9944 -101 10000 -95
rect 9715 -130 9785 -110
rect 9690 -170 9785 -130
rect 9845 -130 9915 -110
rect 9845 -170 9940 -130
rect 9690 -220 9940 -170
rect 9690 -260 9785 -220
rect 9715 -280 9785 -260
rect 9845 -260 9940 -220
rect 9845 -280 9915 -260
rect 9630 -295 9686 -289
rect 9630 -355 9634 -295
rect 9715 -305 9915 -280
rect 9970 -289 10000 -101
rect 9944 -295 10000 -289
rect 9686 -355 9944 -335
rect 9996 -355 10000 -295
rect 9630 -365 10000 -355
rect 10030 -35 10400 -25
rect 10030 -95 10034 -35
rect 10086 -55 10344 -35
rect 10030 -101 10086 -95
rect 10030 -289 10060 -101
rect 10115 -110 10315 -85
rect 10396 -95 10400 -35
rect 10344 -101 10400 -95
rect 10115 -130 10185 -110
rect 10090 -170 10185 -130
rect 10245 -130 10315 -110
rect 10245 -170 10340 -130
rect 10090 -220 10340 -170
rect 10090 -260 10185 -220
rect 10115 -280 10185 -260
rect 10245 -260 10340 -220
rect 10245 -280 10315 -260
rect 10030 -295 10086 -289
rect 10030 -355 10034 -295
rect 10115 -305 10315 -280
rect 10370 -289 10400 -101
rect 10344 -295 10400 -289
rect 10086 -355 10344 -335
rect 10396 -355 10400 -295
rect 10030 -365 10400 -355
rect 10430 -35 10800 -25
rect 10430 -95 10434 -35
rect 10486 -55 10744 -35
rect 10430 -101 10486 -95
rect 10430 -289 10460 -101
rect 10515 -110 10715 -85
rect 10796 -95 10800 -35
rect 10744 -101 10800 -95
rect 10515 -130 10585 -110
rect 10490 -170 10585 -130
rect 10645 -130 10715 -110
rect 10645 -170 10740 -130
rect 10490 -220 10740 -170
rect 10490 -260 10585 -220
rect 10515 -280 10585 -260
rect 10645 -260 10740 -220
rect 10645 -280 10715 -260
rect 10430 -295 10486 -289
rect 10430 -355 10434 -295
rect 10515 -305 10715 -280
rect 10770 -289 10800 -101
rect 10744 -295 10800 -289
rect 10486 -355 10744 -335
rect 10796 -355 10800 -295
rect 10430 -365 10800 -355
rect 10830 -35 11200 -25
rect 10830 -95 10834 -35
rect 10886 -55 11144 -35
rect 10830 -101 10886 -95
rect 10830 -289 10860 -101
rect 10915 -110 11115 -85
rect 11196 -95 11200 -35
rect 11144 -101 11200 -95
rect 10915 -130 10985 -110
rect 10890 -170 10985 -130
rect 11045 -130 11115 -110
rect 11045 -170 11140 -130
rect 10890 -220 11140 -170
rect 10890 -260 10985 -220
rect 10915 -280 10985 -260
rect 11045 -260 11140 -220
rect 11045 -280 11115 -260
rect 10830 -295 10886 -289
rect 10830 -355 10834 -295
rect 10915 -305 11115 -280
rect 11170 -289 11200 -101
rect 11144 -295 11200 -289
rect 10886 -355 11144 -335
rect 11196 -355 11200 -295
rect 10830 -365 11200 -355
rect 11230 -35 11600 -25
rect 11230 -95 11234 -35
rect 11286 -55 11544 -35
rect 11230 -101 11286 -95
rect 11230 -289 11260 -101
rect 11315 -110 11515 -85
rect 11596 -95 11600 -35
rect 11544 -101 11600 -95
rect 11315 -130 11385 -110
rect 11290 -170 11385 -130
rect 11445 -130 11515 -110
rect 11445 -170 11540 -130
rect 11290 -220 11540 -170
rect 11290 -260 11385 -220
rect 11315 -280 11385 -260
rect 11445 -260 11540 -220
rect 11445 -280 11515 -260
rect 11230 -295 11286 -289
rect 11230 -355 11234 -295
rect 11315 -305 11515 -280
rect 11570 -289 11600 -101
rect 11544 -295 11600 -289
rect 11286 -355 11544 -335
rect 11596 -355 11600 -295
rect 11230 -365 11600 -355
rect 11630 -35 12000 -25
rect 11630 -95 11634 -35
rect 11686 -55 11944 -35
rect 11630 -101 11686 -95
rect 11630 -289 11660 -101
rect 11715 -110 11915 -85
rect 11996 -95 12000 -35
rect 11944 -101 12000 -95
rect 11715 -130 11785 -110
rect 11690 -170 11785 -130
rect 11845 -130 11915 -110
rect 11845 -170 11940 -130
rect 11690 -220 11940 -170
rect 11690 -260 11785 -220
rect 11715 -280 11785 -260
rect 11845 -260 11940 -220
rect 11845 -280 11915 -260
rect 11630 -295 11686 -289
rect 11630 -355 11634 -295
rect 11715 -305 11915 -280
rect 11970 -289 12000 -101
rect 11944 -295 12000 -289
rect 11686 -355 11944 -335
rect 11996 -355 12000 -295
rect 11630 -365 12000 -355
rect 12030 -35 12400 -25
rect 12030 -95 12034 -35
rect 12086 -55 12344 -35
rect 12030 -101 12086 -95
rect 12030 -289 12060 -101
rect 12115 -110 12315 -85
rect 12396 -95 12400 -35
rect 12344 -101 12400 -95
rect 12115 -130 12185 -110
rect 12090 -170 12185 -130
rect 12245 -130 12315 -110
rect 12245 -170 12340 -130
rect 12090 -220 12340 -170
rect 12090 -260 12185 -220
rect 12115 -280 12185 -260
rect 12245 -260 12340 -220
rect 12245 -280 12315 -260
rect 12030 -295 12086 -289
rect 12030 -355 12034 -295
rect 12115 -305 12315 -280
rect 12370 -289 12400 -101
rect 12344 -295 12400 -289
rect 12086 -355 12344 -335
rect 12396 -355 12400 -295
rect 12030 -365 12400 -355
rect 12430 -35 12800 -25
rect 12430 -95 12434 -35
rect 12486 -55 12744 -35
rect 12430 -101 12486 -95
rect 12430 -289 12460 -101
rect 12515 -110 12715 -85
rect 12796 -95 12800 -35
rect 12744 -101 12800 -95
rect 12515 -130 12585 -110
rect 12490 -170 12585 -130
rect 12645 -130 12715 -110
rect 12645 -170 12740 -130
rect 12490 -220 12740 -170
rect 12490 -260 12585 -220
rect 12515 -280 12585 -260
rect 12645 -260 12740 -220
rect 12645 -280 12715 -260
rect 12430 -295 12486 -289
rect 12430 -355 12434 -295
rect 12515 -305 12715 -280
rect 12770 -289 12800 -101
rect 12744 -295 12800 -289
rect 12486 -355 12744 -335
rect 12796 -355 12800 -295
rect 12430 -365 12800 -355
rect 12830 -35 13200 -25
rect 12830 -95 12834 -35
rect 12886 -55 13144 -35
rect 12830 -101 12886 -95
rect 12830 -289 12860 -101
rect 12915 -110 13115 -85
rect 13196 -95 13200 -35
rect 13144 -101 13200 -95
rect 12915 -130 12985 -110
rect 12890 -170 12985 -130
rect 13045 -130 13115 -110
rect 13045 -170 13140 -130
rect 12890 -220 13140 -170
rect 12890 -260 12985 -220
rect 12915 -280 12985 -260
rect 13045 -260 13140 -220
rect 13045 -280 13115 -260
rect 12830 -295 12886 -289
rect 12830 -355 12834 -295
rect 12915 -305 13115 -280
rect 13170 -289 13200 -101
rect 13144 -295 13200 -289
rect 12886 -355 13144 -335
rect 13196 -355 13200 -295
rect 12830 -365 13200 -355
<< via2 >>
rect -265 24120 -205 24180
rect -165 24120 -105 24180
rect 12915 24065 12930 24125
rect 12930 24065 12975 24125
rect 13045 24065 13090 24125
rect 13090 24065 13105 24125
rect -215 23880 -155 23940
rect -215 23770 -155 23830
rect 185 23880 245 23940
rect 185 23770 245 23830
rect 585 23880 645 23940
rect 585 23770 645 23830
rect 985 23880 1045 23940
rect 985 23770 1045 23830
rect 1385 23880 1445 23940
rect 1385 23770 1445 23830
rect 1785 23880 1845 23940
rect 1785 23770 1845 23830
rect 2185 23880 2245 23940
rect 2185 23770 2245 23830
rect 2585 23880 2645 23940
rect 2585 23770 2645 23830
rect 2985 23880 3045 23940
rect 2985 23770 3045 23830
rect 3385 23880 3445 23940
rect 3385 23770 3445 23830
rect 3785 23880 3845 23940
rect 3785 23770 3845 23830
rect 4185 23880 4245 23940
rect 4185 23770 4245 23830
rect 4585 23880 4645 23940
rect 4585 23770 4645 23830
rect 4985 23880 5045 23940
rect 4985 23770 5045 23830
rect 5385 23880 5445 23940
rect 5385 23770 5445 23830
rect 5785 23880 5845 23940
rect 5785 23770 5845 23830
rect 6185 23880 6245 23940
rect 6185 23770 6245 23830
rect 6585 23880 6645 23940
rect 6585 23770 6645 23830
rect 6985 23880 7045 23940
rect 6985 23770 7045 23830
rect 7385 23880 7445 23940
rect 7385 23770 7445 23830
rect 7785 23880 7845 23940
rect 7785 23770 7845 23830
rect 8185 23880 8245 23940
rect 8185 23770 8245 23830
rect 8585 23880 8645 23940
rect 8585 23770 8645 23830
rect 8985 23880 9045 23940
rect 8985 23770 9045 23830
rect 9385 23880 9445 23940
rect 9385 23770 9445 23830
rect 9785 23880 9845 23940
rect 9785 23770 9845 23830
rect 10185 23880 10245 23940
rect 10185 23770 10245 23830
rect 10585 23880 10645 23940
rect 10585 23770 10645 23830
rect 10985 23880 11045 23940
rect 10985 23770 11045 23830
rect 11385 23880 11445 23940
rect 11385 23770 11445 23830
rect 11785 23880 11845 23940
rect 11785 23770 11845 23830
rect 12185 23880 12245 23940
rect 12185 23770 12245 23830
rect 12585 23880 12645 23940
rect 12585 23770 12645 23830
rect 12985 23880 13045 23940
rect 12985 23770 13045 23830
rect -215 23510 -155 23570
rect -215 23400 -155 23460
rect 185 23510 245 23570
rect 185 23400 245 23460
rect 585 23510 645 23570
rect 585 23400 645 23460
rect 985 23510 1045 23570
rect 985 23400 1045 23460
rect 1385 23510 1445 23570
rect 1385 23400 1445 23460
rect 1785 23510 1845 23570
rect 1785 23400 1845 23460
rect 2185 23510 2245 23570
rect 2185 23400 2245 23460
rect 2585 23510 2645 23570
rect 2585 23400 2645 23460
rect 2985 23510 3045 23570
rect 2985 23400 3045 23460
rect 3385 23510 3445 23570
rect 3385 23400 3445 23460
rect 3785 23510 3845 23570
rect 3785 23400 3845 23460
rect 4185 23510 4245 23570
rect 4185 23400 4245 23460
rect 4585 23510 4645 23570
rect 4585 23400 4645 23460
rect 4985 23510 5045 23570
rect 4985 23400 5045 23460
rect 5385 23510 5445 23570
rect 5385 23400 5445 23460
rect 5785 23510 5845 23570
rect 5785 23400 5845 23460
rect 6185 23510 6245 23570
rect 6185 23400 6245 23460
rect 6585 23510 6645 23570
rect 6585 23400 6645 23460
rect 6985 23510 7045 23570
rect 6985 23400 7045 23460
rect 7385 23510 7445 23570
rect 7385 23400 7445 23460
rect 7785 23510 7845 23570
rect 7785 23400 7845 23460
rect 8185 23510 8245 23570
rect 8185 23400 8245 23460
rect 8585 23510 8645 23570
rect 8585 23400 8645 23460
rect 8985 23510 9045 23570
rect 8985 23400 9045 23460
rect 9385 23510 9445 23570
rect 9385 23400 9445 23460
rect 9785 23510 9845 23570
rect 9785 23400 9845 23460
rect 10185 23510 10245 23570
rect 10185 23400 10245 23460
rect 10585 23510 10645 23570
rect 10585 23400 10645 23460
rect 10985 23510 11045 23570
rect 10985 23400 11045 23460
rect 11385 23510 11445 23570
rect 11385 23400 11445 23460
rect 11785 23510 11845 23570
rect 11785 23400 11845 23460
rect 12185 23510 12245 23570
rect 12185 23400 12245 23460
rect 12585 23510 12645 23570
rect 12585 23400 12645 23460
rect 12985 23510 13045 23570
rect 12985 23400 13045 23460
rect -215 23140 -155 23200
rect -215 23030 -155 23090
rect 185 23140 245 23200
rect 185 23030 245 23090
rect 585 23140 645 23200
rect 585 23030 645 23090
rect 985 23140 1045 23200
rect 985 23030 1045 23090
rect 1385 23140 1445 23200
rect 1385 23030 1445 23090
rect 1785 23140 1845 23200
rect 1785 23030 1845 23090
rect 2185 23140 2245 23200
rect 2185 23030 2245 23090
rect 2585 23140 2645 23200
rect 2585 23030 2645 23090
rect 2985 23140 3045 23200
rect 2985 23030 3045 23090
rect 3385 23140 3445 23200
rect 3385 23030 3445 23090
rect 3785 23140 3845 23200
rect 3785 23030 3845 23090
rect 4185 23140 4245 23200
rect 4185 23030 4245 23090
rect 4585 23140 4645 23200
rect 4585 23030 4645 23090
rect 4985 23140 5045 23200
rect 4985 23030 5045 23090
rect 5385 23140 5445 23200
rect 5385 23030 5445 23090
rect 5785 23140 5845 23200
rect 5785 23030 5845 23090
rect 6185 23140 6245 23200
rect 6185 23030 6245 23090
rect 6585 23140 6645 23200
rect 6585 23030 6645 23090
rect 6985 23140 7045 23200
rect 6985 23030 7045 23090
rect 7385 23140 7445 23200
rect 7385 23030 7445 23090
rect 7785 23140 7845 23200
rect 7785 23030 7845 23090
rect 8185 23140 8245 23200
rect 8185 23030 8245 23090
rect 8585 23140 8645 23200
rect 8585 23030 8645 23090
rect 8985 23140 9045 23200
rect 8985 23030 9045 23090
rect 9385 23140 9445 23200
rect 9385 23030 9445 23090
rect 9785 23140 9845 23200
rect 9785 23030 9845 23090
rect 10185 23140 10245 23200
rect 10185 23030 10245 23090
rect 10585 23140 10645 23200
rect 10585 23030 10645 23090
rect 10985 23140 11045 23200
rect 10985 23030 11045 23090
rect 11385 23140 11445 23200
rect 11385 23030 11445 23090
rect 11785 23140 11845 23200
rect 11785 23030 11845 23090
rect 12185 23140 12245 23200
rect 12185 23030 12245 23090
rect 12585 23140 12645 23200
rect 12585 23030 12645 23090
rect 12985 23140 13045 23200
rect 12985 23030 13045 23090
rect -215 22770 -155 22830
rect -215 22660 -155 22720
rect 185 22770 245 22830
rect 185 22660 245 22720
rect 585 22770 645 22830
rect 585 22660 645 22720
rect 985 22770 1045 22830
rect 985 22660 1045 22720
rect 1385 22770 1445 22830
rect 1385 22660 1445 22720
rect 1785 22770 1845 22830
rect 1785 22660 1845 22720
rect 2185 22770 2245 22830
rect 2185 22660 2245 22720
rect 2585 22770 2645 22830
rect 2585 22660 2645 22720
rect 2985 22770 3045 22830
rect 2985 22660 3045 22720
rect 3385 22770 3445 22830
rect 3385 22660 3445 22720
rect 3785 22770 3845 22830
rect 3785 22660 3845 22720
rect 4185 22770 4245 22830
rect 4185 22660 4245 22720
rect 4585 22770 4645 22830
rect 4585 22660 4645 22720
rect 4985 22770 5045 22830
rect 4985 22660 5045 22720
rect 5385 22770 5445 22830
rect 5385 22660 5445 22720
rect 5785 22770 5845 22830
rect 5785 22660 5845 22720
rect 6185 22770 6245 22830
rect 6185 22660 6245 22720
rect 6585 22770 6645 22830
rect 6585 22660 6645 22720
rect 6985 22770 7045 22830
rect 6985 22660 7045 22720
rect 7385 22770 7445 22830
rect 7385 22660 7445 22720
rect 7785 22770 7845 22830
rect 7785 22660 7845 22720
rect 8185 22770 8245 22830
rect 8185 22660 8245 22720
rect 8585 22770 8645 22830
rect 8585 22660 8645 22720
rect 8985 22770 9045 22830
rect 8985 22660 9045 22720
rect 9385 22770 9445 22830
rect 9385 22660 9445 22720
rect 9785 22770 9845 22830
rect 9785 22660 9845 22720
rect 10185 22770 10245 22830
rect 10185 22660 10245 22720
rect 10585 22770 10645 22830
rect 10585 22660 10645 22720
rect 10985 22770 11045 22830
rect 10985 22660 11045 22720
rect 11385 22770 11445 22830
rect 11385 22660 11445 22720
rect 11785 22770 11845 22830
rect 11785 22660 11845 22720
rect 12185 22770 12245 22830
rect 12185 22660 12245 22720
rect 12585 22770 12645 22830
rect 12585 22660 12645 22720
rect 12985 22770 13045 22830
rect 12985 22660 13045 22720
rect -215 22400 -155 22460
rect -215 22290 -155 22350
rect 185 22400 245 22460
rect 185 22290 245 22350
rect 585 22400 645 22460
rect 585 22290 645 22350
rect 985 22400 1045 22460
rect 985 22290 1045 22350
rect 1385 22400 1445 22460
rect 1385 22290 1445 22350
rect 1785 22400 1845 22460
rect 1785 22290 1845 22350
rect 2185 22400 2245 22460
rect 2185 22290 2245 22350
rect 2585 22400 2645 22460
rect 2585 22290 2645 22350
rect 2985 22400 3045 22460
rect 2985 22290 3045 22350
rect 3385 22400 3445 22460
rect 3385 22290 3445 22350
rect 3785 22400 3845 22460
rect 3785 22290 3845 22350
rect 4185 22400 4245 22460
rect 4185 22290 4245 22350
rect 4585 22400 4645 22460
rect 4585 22290 4645 22350
rect 4985 22400 5045 22460
rect 4985 22290 5045 22350
rect 5385 22400 5445 22460
rect 5385 22290 5445 22350
rect 5785 22400 5845 22460
rect 5785 22290 5845 22350
rect 6185 22400 6245 22460
rect 6185 22290 6245 22350
rect 6585 22400 6645 22460
rect 6585 22290 6645 22350
rect 6985 22400 7045 22460
rect 6985 22290 7045 22350
rect 7385 22400 7445 22460
rect 7385 22290 7445 22350
rect 7785 22400 7845 22460
rect 7785 22290 7845 22350
rect 8185 22400 8245 22460
rect 8185 22290 8245 22350
rect 8585 22400 8645 22460
rect 8585 22290 8645 22350
rect 8985 22400 9045 22460
rect 8985 22290 9045 22350
rect 9385 22400 9445 22460
rect 9385 22290 9445 22350
rect 9785 22400 9845 22460
rect 9785 22290 9845 22350
rect 10185 22400 10245 22460
rect 10185 22290 10245 22350
rect 10585 22400 10645 22460
rect 10585 22290 10645 22350
rect 10985 22400 11045 22460
rect 10985 22290 11045 22350
rect 11385 22400 11445 22460
rect 11385 22290 11445 22350
rect 11785 22400 11845 22460
rect 11785 22290 11845 22350
rect 12185 22400 12245 22460
rect 12185 22290 12245 22350
rect 12585 22400 12645 22460
rect 12585 22290 12645 22350
rect 12985 22400 13045 22460
rect 12985 22290 13045 22350
rect -215 22030 -155 22090
rect -215 21920 -155 21980
rect 185 22030 245 22090
rect 185 21920 245 21980
rect 585 22030 645 22090
rect 585 21920 645 21980
rect 985 22030 1045 22090
rect 985 21920 1045 21980
rect 1385 22030 1445 22090
rect 1385 21920 1445 21980
rect 1785 22030 1845 22090
rect 1785 21920 1845 21980
rect 2185 22030 2245 22090
rect 2185 21920 2245 21980
rect 2585 22030 2645 22090
rect 2585 21920 2645 21980
rect 2985 22030 3045 22090
rect 2985 21920 3045 21980
rect 3385 22030 3445 22090
rect 3385 21920 3445 21980
rect 3785 22030 3845 22090
rect 3785 21920 3845 21980
rect 4185 22030 4245 22090
rect 4185 21920 4245 21980
rect 4585 22030 4645 22090
rect 4585 21920 4645 21980
rect 4985 22030 5045 22090
rect 4985 21920 5045 21980
rect 5385 22030 5445 22090
rect 5385 21920 5445 21980
rect 5785 22030 5845 22090
rect 5785 21920 5845 21980
rect 6185 22030 6245 22090
rect 6185 21920 6245 21980
rect 6585 22030 6645 22090
rect 6585 21920 6645 21980
rect 6985 22030 7045 22090
rect 6985 21920 7045 21980
rect 7385 22030 7445 22090
rect 7385 21920 7445 21980
rect 7785 22030 7845 22090
rect 7785 21920 7845 21980
rect 8185 22030 8245 22090
rect 8185 21920 8245 21980
rect 8585 22030 8645 22090
rect 8585 21920 8645 21980
rect 8985 22030 9045 22090
rect 8985 21920 9045 21980
rect 9385 22030 9445 22090
rect 9385 21920 9445 21980
rect 9785 22030 9845 22090
rect 9785 21920 9845 21980
rect 10185 22030 10245 22090
rect 10185 21920 10245 21980
rect 10585 22030 10645 22090
rect 10585 21920 10645 21980
rect 10985 22030 11045 22090
rect 10985 21920 11045 21980
rect 11385 22030 11445 22090
rect 11385 21920 11445 21980
rect 11785 22030 11845 22090
rect 11785 21920 11845 21980
rect 12185 22030 12245 22090
rect 12185 21920 12245 21980
rect 12585 22030 12645 22090
rect 12585 21920 12645 21980
rect 12985 22030 13045 22090
rect 12985 21920 13045 21980
rect -215 21660 -155 21720
rect -215 21550 -155 21610
rect 185 21660 245 21720
rect 185 21550 245 21610
rect 585 21660 645 21720
rect 585 21550 645 21610
rect 985 21660 1045 21720
rect 985 21550 1045 21610
rect 1385 21660 1445 21720
rect 1385 21550 1445 21610
rect 1785 21660 1845 21720
rect 1785 21550 1845 21610
rect 2185 21660 2245 21720
rect 2185 21550 2245 21610
rect 2585 21660 2645 21720
rect 2585 21550 2645 21610
rect 2985 21660 3045 21720
rect 2985 21550 3045 21610
rect 3385 21660 3445 21720
rect 3385 21550 3445 21610
rect 3785 21660 3845 21720
rect 3785 21550 3845 21610
rect 4185 21660 4245 21720
rect 4185 21550 4245 21610
rect 4585 21660 4645 21720
rect 4585 21550 4645 21610
rect 4985 21660 5045 21720
rect 4985 21550 5045 21610
rect 5385 21660 5445 21720
rect 5385 21550 5445 21610
rect 5785 21660 5845 21720
rect 5785 21550 5845 21610
rect 6185 21660 6245 21720
rect 6185 21550 6245 21610
rect 6585 21660 6645 21720
rect 6585 21550 6645 21610
rect 6985 21660 7045 21720
rect 6985 21550 7045 21610
rect 7385 21660 7445 21720
rect 7385 21550 7445 21610
rect 7785 21660 7845 21720
rect 7785 21550 7845 21610
rect 8185 21660 8245 21720
rect 8185 21550 8245 21610
rect 8585 21660 8645 21720
rect 8585 21550 8645 21610
rect 8985 21660 9045 21720
rect 8985 21550 9045 21610
rect 9385 21660 9445 21720
rect 9385 21550 9445 21610
rect 9785 21660 9845 21720
rect 9785 21550 9845 21610
rect 10185 21660 10245 21720
rect 10185 21550 10245 21610
rect 10585 21660 10645 21720
rect 10585 21550 10645 21610
rect 10985 21660 11045 21720
rect 10985 21550 11045 21610
rect 11385 21660 11445 21720
rect 11385 21550 11445 21610
rect 11785 21660 11845 21720
rect 11785 21550 11845 21610
rect 12185 21660 12245 21720
rect 12185 21550 12245 21610
rect 12585 21660 12645 21720
rect 12585 21550 12645 21610
rect 12985 21660 13045 21720
rect 12985 21550 13045 21610
rect -215 21290 -155 21350
rect -215 21180 -155 21240
rect 185 21290 245 21350
rect 185 21180 245 21240
rect 585 21290 645 21350
rect 585 21180 645 21240
rect 985 21290 1045 21350
rect 985 21180 1045 21240
rect 1385 21290 1445 21350
rect 1385 21180 1445 21240
rect 1785 21290 1845 21350
rect 1785 21180 1845 21240
rect 2185 21290 2245 21350
rect 2185 21180 2245 21240
rect 2585 21290 2645 21350
rect 2585 21180 2645 21240
rect 2985 21290 3045 21350
rect 2985 21180 3045 21240
rect 3385 21290 3445 21350
rect 3385 21180 3445 21240
rect 3785 21290 3845 21350
rect 3785 21180 3845 21240
rect 4185 21290 4245 21350
rect 4185 21180 4245 21240
rect 4585 21290 4645 21350
rect 4585 21180 4645 21240
rect 4985 21290 5045 21350
rect 4985 21180 5045 21240
rect 5385 21290 5445 21350
rect 5385 21180 5445 21240
rect 5785 21290 5845 21350
rect 5785 21180 5845 21240
rect 6185 21290 6245 21350
rect 6185 21180 6245 21240
rect 6585 21290 6645 21350
rect 6585 21180 6645 21240
rect 6985 21290 7045 21350
rect 6985 21180 7045 21240
rect 7385 21290 7445 21350
rect 7385 21180 7445 21240
rect 7785 21290 7845 21350
rect 7785 21180 7845 21240
rect 8185 21290 8245 21350
rect 8185 21180 8245 21240
rect 8585 21290 8645 21350
rect 8585 21180 8645 21240
rect 8985 21290 9045 21350
rect 8985 21180 9045 21240
rect 9385 21290 9445 21350
rect 9385 21180 9445 21240
rect 9785 21290 9845 21350
rect 9785 21180 9845 21240
rect 10185 21290 10245 21350
rect 10185 21180 10245 21240
rect 10585 21290 10645 21350
rect 10585 21180 10645 21240
rect 10985 21290 11045 21350
rect 10985 21180 11045 21240
rect 11385 21290 11445 21350
rect 11385 21180 11445 21240
rect 11785 21290 11845 21350
rect 11785 21180 11845 21240
rect 12185 21290 12245 21350
rect 12185 21180 12245 21240
rect 12585 21290 12645 21350
rect 12585 21180 12645 21240
rect 12985 21290 13045 21350
rect 12985 21180 13045 21240
rect -215 20920 -155 20980
rect -215 20810 -155 20870
rect 185 20920 245 20980
rect 185 20810 245 20870
rect 585 20920 645 20980
rect 585 20810 645 20870
rect 985 20920 1045 20980
rect 985 20810 1045 20870
rect 1385 20920 1445 20980
rect 1385 20810 1445 20870
rect 1785 20920 1845 20980
rect 1785 20810 1845 20870
rect 2185 20920 2245 20980
rect 2185 20810 2245 20870
rect 2585 20920 2645 20980
rect 2585 20810 2645 20870
rect 2985 20920 3045 20980
rect 2985 20810 3045 20870
rect 3385 20920 3445 20980
rect 3385 20810 3445 20870
rect 3785 20920 3845 20980
rect 3785 20810 3845 20870
rect 4185 20920 4245 20980
rect 4185 20810 4245 20870
rect 4585 20920 4645 20980
rect 4585 20810 4645 20870
rect 4985 20920 5045 20980
rect 4985 20810 5045 20870
rect 5385 20920 5445 20980
rect 5385 20810 5445 20870
rect 5785 20920 5845 20980
rect 5785 20810 5845 20870
rect 6185 20920 6245 20980
rect 6185 20810 6245 20870
rect 6585 20920 6645 20980
rect 6585 20810 6645 20870
rect 6985 20920 7045 20980
rect 6985 20810 7045 20870
rect 7385 20920 7445 20980
rect 7385 20810 7445 20870
rect 7785 20920 7845 20980
rect 7785 20810 7845 20870
rect 8185 20920 8245 20980
rect 8185 20810 8245 20870
rect 8585 20920 8645 20980
rect 8585 20810 8645 20870
rect 8985 20920 9045 20980
rect 8985 20810 9045 20870
rect 9385 20920 9445 20980
rect 9385 20810 9445 20870
rect 9785 20920 9845 20980
rect 9785 20810 9845 20870
rect 10185 20920 10245 20980
rect 10185 20810 10245 20870
rect 10585 20920 10645 20980
rect 10585 20810 10645 20870
rect 10985 20920 11045 20980
rect 10985 20810 11045 20870
rect 11385 20920 11445 20980
rect 11385 20810 11445 20870
rect 11785 20920 11845 20980
rect 11785 20810 11845 20870
rect 12185 20920 12245 20980
rect 12185 20810 12245 20870
rect 12585 20920 12645 20980
rect 12585 20810 12645 20870
rect 12985 20920 13045 20980
rect 12985 20810 13045 20870
rect -215 20550 -155 20610
rect -215 20440 -155 20500
rect 185 20550 245 20610
rect 185 20440 245 20500
rect 585 20550 645 20610
rect 585 20440 645 20500
rect 985 20550 1045 20610
rect 985 20440 1045 20500
rect 1385 20550 1445 20610
rect 1385 20440 1445 20500
rect 1785 20550 1845 20610
rect 1785 20440 1845 20500
rect 2185 20550 2245 20610
rect 2185 20440 2245 20500
rect 2585 20550 2645 20610
rect 2585 20440 2645 20500
rect 2985 20550 3045 20610
rect 2985 20440 3045 20500
rect 3385 20550 3445 20610
rect 3385 20440 3445 20500
rect 3785 20550 3845 20610
rect 3785 20440 3845 20500
rect 4185 20550 4245 20610
rect 4185 20440 4245 20500
rect 4585 20550 4645 20610
rect 4585 20440 4645 20500
rect 4985 20550 5045 20610
rect 4985 20440 5045 20500
rect 5385 20550 5445 20610
rect 5385 20440 5445 20500
rect 5785 20550 5845 20610
rect 5785 20440 5845 20500
rect 6185 20550 6245 20610
rect 6185 20440 6245 20500
rect 6585 20550 6645 20610
rect 6585 20440 6645 20500
rect 6985 20550 7045 20610
rect 6985 20440 7045 20500
rect 7385 20550 7445 20610
rect 7385 20440 7445 20500
rect 7785 20550 7845 20610
rect 7785 20440 7845 20500
rect 8185 20550 8245 20610
rect 8185 20440 8245 20500
rect 8585 20550 8645 20610
rect 8585 20440 8645 20500
rect 8985 20550 9045 20610
rect 8985 20440 9045 20500
rect 9385 20550 9445 20610
rect 9385 20440 9445 20500
rect 9785 20550 9845 20610
rect 9785 20440 9845 20500
rect 10185 20550 10245 20610
rect 10185 20440 10245 20500
rect 10585 20550 10645 20610
rect 10585 20440 10645 20500
rect 10985 20550 11045 20610
rect 10985 20440 11045 20500
rect 11385 20550 11445 20610
rect 11385 20440 11445 20500
rect 11785 20550 11845 20610
rect 11785 20440 11845 20500
rect 12185 20550 12245 20610
rect 12185 20440 12245 20500
rect 12585 20550 12645 20610
rect 12585 20440 12645 20500
rect 12985 20550 13045 20610
rect 12985 20440 13045 20500
rect -215 20180 -155 20240
rect -215 20070 -155 20130
rect 185 20180 245 20240
rect 185 20070 245 20130
rect 585 20180 645 20240
rect 585 20070 645 20130
rect 985 20180 1045 20240
rect 985 20070 1045 20130
rect 1385 20180 1445 20240
rect 1385 20070 1445 20130
rect 1785 20180 1845 20240
rect 1785 20070 1845 20130
rect 2185 20180 2245 20240
rect 2185 20070 2245 20130
rect 2585 20180 2645 20240
rect 2585 20070 2645 20130
rect 2985 20180 3045 20240
rect 2985 20070 3045 20130
rect 3385 20180 3445 20240
rect 3385 20070 3445 20130
rect 3785 20180 3845 20240
rect 3785 20070 3845 20130
rect 4185 20180 4245 20240
rect 4185 20070 4245 20130
rect 4585 20180 4645 20240
rect 4585 20070 4645 20130
rect 4985 20180 5045 20240
rect 4985 20070 5045 20130
rect 5385 20180 5445 20240
rect 5385 20070 5445 20130
rect 5785 20180 5845 20240
rect 5785 20070 5845 20130
rect 6185 20180 6245 20240
rect 6185 20070 6245 20130
rect 6585 20180 6645 20240
rect 6585 20070 6645 20130
rect 6985 20180 7045 20240
rect 6985 20070 7045 20130
rect 7385 20180 7445 20240
rect 7385 20070 7445 20130
rect 7785 20180 7845 20240
rect 7785 20070 7845 20130
rect 8185 20180 8245 20240
rect 8185 20070 8245 20130
rect 8585 20180 8645 20240
rect 8585 20070 8645 20130
rect 8985 20180 9045 20240
rect 8985 20070 9045 20130
rect 9385 20180 9445 20240
rect 9385 20070 9445 20130
rect 9785 20180 9845 20240
rect 9785 20070 9845 20130
rect 10185 20180 10245 20240
rect 10185 20070 10245 20130
rect 10585 20180 10645 20240
rect 10585 20070 10645 20130
rect 10985 20180 11045 20240
rect 10985 20070 11045 20130
rect 11385 20180 11445 20240
rect 11385 20070 11445 20130
rect 11785 20180 11845 20240
rect 11785 20070 11845 20130
rect 12185 20180 12245 20240
rect 12185 20070 12245 20130
rect 12585 20180 12645 20240
rect 12585 20070 12645 20130
rect 12985 20180 13045 20240
rect 12985 20070 13045 20130
rect -215 19810 -155 19870
rect -215 19700 -155 19760
rect 185 19810 245 19870
rect 185 19700 245 19760
rect 585 19810 645 19870
rect 585 19700 645 19760
rect 985 19810 1045 19870
rect 985 19700 1045 19760
rect 1385 19810 1445 19870
rect 1385 19700 1445 19760
rect 1785 19810 1845 19870
rect 1785 19700 1845 19760
rect 2185 19810 2245 19870
rect 2185 19700 2245 19760
rect 2585 19810 2645 19870
rect 2585 19700 2645 19760
rect 2985 19810 3045 19870
rect 2985 19700 3045 19760
rect 3385 19810 3445 19870
rect 3385 19700 3445 19760
rect 3785 19810 3845 19870
rect 3785 19700 3845 19760
rect 4185 19810 4245 19870
rect 4185 19700 4245 19760
rect 4585 19810 4645 19870
rect 4585 19700 4645 19760
rect 4985 19810 5045 19870
rect 4985 19700 5045 19760
rect 5385 19810 5445 19870
rect 5385 19700 5445 19760
rect 5785 19810 5845 19870
rect 5785 19700 5845 19760
rect 6185 19810 6245 19870
rect 6185 19700 6245 19760
rect 6585 19810 6645 19870
rect 6585 19700 6645 19760
rect 6985 19810 7045 19870
rect 6985 19700 7045 19760
rect 7385 19810 7445 19870
rect 7385 19700 7445 19760
rect 7785 19810 7845 19870
rect 7785 19700 7845 19760
rect 8185 19810 8245 19870
rect 8185 19700 8245 19760
rect 8585 19810 8645 19870
rect 8585 19700 8645 19760
rect 8985 19810 9045 19870
rect 8985 19700 9045 19760
rect 9385 19810 9445 19870
rect 9385 19700 9445 19760
rect 9785 19810 9845 19870
rect 9785 19700 9845 19760
rect 10185 19810 10245 19870
rect 10185 19700 10245 19760
rect 10585 19810 10645 19870
rect 10585 19700 10645 19760
rect 10985 19810 11045 19870
rect 10985 19700 11045 19760
rect 11385 19810 11445 19870
rect 11385 19700 11445 19760
rect 11785 19810 11845 19870
rect 11785 19700 11845 19760
rect 12185 19810 12245 19870
rect 12185 19700 12245 19760
rect 12585 19810 12645 19870
rect 12585 19700 12645 19760
rect 12985 19810 13045 19870
rect 12985 19700 13045 19760
rect -215 19440 -155 19500
rect -215 19330 -155 19390
rect 185 19440 245 19500
rect 185 19330 245 19390
rect 585 19440 645 19500
rect 585 19330 645 19390
rect 985 19440 1045 19500
rect 985 19330 1045 19390
rect 1385 19440 1445 19500
rect 1385 19330 1445 19390
rect 1785 19440 1845 19500
rect 1785 19330 1845 19390
rect 2185 19440 2245 19500
rect 2185 19330 2245 19390
rect 2585 19440 2645 19500
rect 2585 19330 2645 19390
rect 2985 19440 3045 19500
rect 2985 19330 3045 19390
rect 3385 19440 3445 19500
rect 3385 19330 3445 19390
rect 3785 19440 3845 19500
rect 3785 19330 3845 19390
rect 4185 19440 4245 19500
rect 4185 19330 4245 19390
rect 4585 19440 4645 19500
rect 4585 19330 4645 19390
rect 4985 19440 5045 19500
rect 4985 19330 5045 19390
rect 5385 19440 5445 19500
rect 5385 19330 5445 19390
rect 5785 19440 5845 19500
rect 5785 19330 5845 19390
rect 6185 19440 6245 19500
rect 6185 19330 6245 19390
rect 6585 19440 6645 19500
rect 6585 19330 6645 19390
rect 6985 19440 7045 19500
rect 6985 19330 7045 19390
rect 7385 19440 7445 19500
rect 7385 19330 7445 19390
rect 7785 19440 7845 19500
rect 7785 19330 7845 19390
rect 8185 19440 8245 19500
rect 8185 19330 8245 19390
rect 8585 19440 8645 19500
rect 8585 19330 8645 19390
rect 8985 19440 9045 19500
rect 8985 19330 9045 19390
rect 9385 19440 9445 19500
rect 9385 19330 9445 19390
rect 9785 19440 9845 19500
rect 9785 19330 9845 19390
rect 10185 19440 10245 19500
rect 10185 19330 10245 19390
rect 10585 19440 10645 19500
rect 10585 19330 10645 19390
rect 10985 19440 11045 19500
rect 10985 19330 11045 19390
rect 11385 19440 11445 19500
rect 11385 19330 11445 19390
rect 11785 19440 11845 19500
rect 11785 19330 11845 19390
rect 12185 19440 12245 19500
rect 12185 19330 12245 19390
rect 12585 19440 12645 19500
rect 12585 19330 12645 19390
rect 12985 19440 13045 19500
rect 12985 19330 13045 19390
rect -215 19070 -155 19130
rect -215 18960 -155 19020
rect 185 19070 245 19130
rect 185 18960 245 19020
rect 585 19070 645 19130
rect 585 18960 645 19020
rect 985 19070 1045 19130
rect 985 18960 1045 19020
rect 1385 19070 1445 19130
rect 1385 18960 1445 19020
rect 1785 19070 1845 19130
rect 1785 18960 1845 19020
rect 2185 19070 2245 19130
rect 2185 18960 2245 19020
rect 2585 19070 2645 19130
rect 2585 18960 2645 19020
rect 2985 19070 3045 19130
rect 2985 18960 3045 19020
rect 3385 19070 3445 19130
rect 3385 18960 3445 19020
rect 3785 19070 3845 19130
rect 3785 18960 3845 19020
rect 4185 19070 4245 19130
rect 4185 18960 4245 19020
rect 4585 19070 4645 19130
rect 4585 18960 4645 19020
rect 4985 19070 5045 19130
rect 4985 18960 5045 19020
rect 5385 19070 5445 19130
rect 5385 18960 5445 19020
rect 5785 19070 5845 19130
rect 5785 18960 5845 19020
rect 6185 19070 6245 19130
rect 6185 18960 6245 19020
rect 6585 19070 6645 19130
rect 6585 18960 6645 19020
rect 6985 19070 7045 19130
rect 6985 18960 7045 19020
rect 7385 19070 7445 19130
rect 7385 18960 7445 19020
rect 7785 19070 7845 19130
rect 7785 18960 7845 19020
rect 8185 19070 8245 19130
rect 8185 18960 8245 19020
rect 8585 19070 8645 19130
rect 8585 18960 8645 19020
rect 8985 19070 9045 19130
rect 8985 18960 9045 19020
rect 9385 19070 9445 19130
rect 9385 18960 9445 19020
rect 9785 19070 9845 19130
rect 9785 18960 9845 19020
rect 10185 19070 10245 19130
rect 10185 18960 10245 19020
rect 10585 19070 10645 19130
rect 10585 18960 10645 19020
rect 10985 19070 11045 19130
rect 10985 18960 11045 19020
rect 11385 19070 11445 19130
rect 11385 18960 11445 19020
rect 11785 19070 11845 19130
rect 11785 18960 11845 19020
rect 12185 19070 12245 19130
rect 12185 18960 12245 19020
rect 12585 19070 12645 19130
rect 12585 18960 12645 19020
rect 12985 19070 13045 19130
rect 12985 18960 13045 19020
rect -215 18700 -155 18760
rect -215 18590 -155 18650
rect 185 18700 245 18760
rect 185 18590 245 18650
rect 585 18700 645 18760
rect 585 18590 645 18650
rect 985 18700 1045 18760
rect 985 18590 1045 18650
rect 1385 18700 1445 18760
rect 1385 18590 1445 18650
rect 1785 18700 1845 18760
rect 1785 18590 1845 18650
rect 2185 18700 2245 18760
rect 2185 18590 2245 18650
rect 2585 18700 2645 18760
rect 2585 18590 2645 18650
rect 2985 18700 3045 18760
rect 2985 18590 3045 18650
rect 3385 18700 3445 18760
rect 3385 18590 3445 18650
rect 3785 18700 3845 18760
rect 3785 18590 3845 18650
rect 4185 18700 4245 18760
rect 4185 18590 4245 18650
rect 4585 18700 4645 18760
rect 4585 18590 4645 18650
rect 4985 18700 5045 18760
rect 4985 18590 5045 18650
rect 5385 18700 5445 18760
rect 5385 18590 5445 18650
rect 5785 18700 5845 18760
rect 5785 18590 5845 18650
rect 6185 18700 6245 18760
rect 6185 18590 6245 18650
rect 6585 18700 6645 18760
rect 6585 18590 6645 18650
rect 6985 18700 7045 18760
rect 6985 18590 7045 18650
rect 7385 18700 7445 18760
rect 7385 18590 7445 18650
rect 7785 18700 7845 18760
rect 7785 18590 7845 18650
rect 8185 18700 8245 18760
rect 8185 18590 8245 18650
rect 8585 18700 8645 18760
rect 8585 18590 8645 18650
rect 8985 18700 9045 18760
rect 8985 18590 9045 18650
rect 9385 18700 9445 18760
rect 9385 18590 9445 18650
rect 9785 18700 9845 18760
rect 9785 18590 9845 18650
rect 10185 18700 10245 18760
rect 10185 18590 10245 18650
rect 10585 18700 10645 18760
rect 10585 18590 10645 18650
rect 10985 18700 11045 18760
rect 10985 18590 11045 18650
rect 11385 18700 11445 18760
rect 11385 18590 11445 18650
rect 11785 18700 11845 18760
rect 11785 18590 11845 18650
rect 12185 18700 12245 18760
rect 12185 18590 12245 18650
rect 12585 18700 12645 18760
rect 12585 18590 12645 18650
rect 12985 18700 13045 18760
rect 12985 18590 13045 18650
rect -215 18330 -155 18390
rect -215 18220 -155 18280
rect 185 18330 245 18390
rect 185 18220 245 18280
rect 585 18330 645 18390
rect 585 18220 645 18280
rect 985 18330 1045 18390
rect 985 18220 1045 18280
rect 1385 18330 1445 18390
rect 1385 18220 1445 18280
rect 1785 18330 1845 18390
rect 1785 18220 1845 18280
rect 2185 18330 2245 18390
rect 2185 18220 2245 18280
rect 2585 18330 2645 18390
rect 2585 18220 2645 18280
rect 2985 18330 3045 18390
rect 2985 18220 3045 18280
rect 3385 18330 3445 18390
rect 3385 18220 3445 18280
rect 3785 18330 3845 18390
rect 3785 18220 3845 18280
rect 4185 18330 4245 18390
rect 4185 18220 4245 18280
rect 4585 18330 4645 18390
rect 4585 18220 4645 18280
rect 4985 18330 5045 18390
rect 4985 18220 5045 18280
rect 5385 18330 5445 18390
rect 5385 18220 5445 18280
rect 5785 18330 5845 18390
rect 5785 18220 5845 18280
rect 6185 18330 6245 18390
rect 6185 18220 6245 18280
rect 6585 18330 6645 18390
rect 6585 18220 6645 18280
rect 6985 18330 7045 18390
rect 6985 18220 7045 18280
rect 7385 18330 7445 18390
rect 7385 18220 7445 18280
rect 7785 18330 7845 18390
rect 7785 18220 7845 18280
rect 8185 18330 8245 18390
rect 8185 18220 8245 18280
rect 8585 18330 8645 18390
rect 8585 18220 8645 18280
rect 8985 18330 9045 18390
rect 8985 18220 9045 18280
rect 9385 18330 9445 18390
rect 9385 18220 9445 18280
rect 9785 18330 9845 18390
rect 9785 18220 9845 18280
rect 10185 18330 10245 18390
rect 10185 18220 10245 18280
rect 10585 18330 10645 18390
rect 10585 18220 10645 18280
rect 10985 18330 11045 18390
rect 10985 18220 11045 18280
rect 11385 18330 11445 18390
rect 11385 18220 11445 18280
rect 11785 18330 11845 18390
rect 11785 18220 11845 18280
rect 12185 18330 12245 18390
rect 12185 18220 12245 18280
rect 12585 18330 12645 18390
rect 12585 18220 12645 18280
rect 12985 18330 13045 18390
rect 12985 18220 13045 18280
rect -215 17960 -155 18020
rect -215 17850 -155 17910
rect 185 17960 245 18020
rect 185 17850 245 17910
rect 585 17960 645 18020
rect 585 17850 645 17910
rect 985 17960 1045 18020
rect 985 17850 1045 17910
rect 1385 17960 1445 18020
rect 1385 17850 1445 17910
rect 1785 17960 1845 18020
rect 1785 17850 1845 17910
rect 2185 17960 2245 18020
rect 2185 17850 2245 17910
rect 2585 17960 2645 18020
rect 2585 17850 2645 17910
rect 2985 17960 3045 18020
rect 2985 17850 3045 17910
rect 3385 17960 3445 18020
rect 3385 17850 3445 17910
rect 3785 17960 3845 18020
rect 3785 17850 3845 17910
rect 4185 17960 4245 18020
rect 4185 17850 4245 17910
rect 4585 17960 4645 18020
rect 4585 17850 4645 17910
rect 4985 17960 5045 18020
rect 4985 17850 5045 17910
rect 5385 17960 5445 18020
rect 5385 17850 5445 17910
rect 5785 17960 5845 18020
rect 5785 17850 5845 17910
rect 6185 17960 6245 18020
rect 6185 17850 6245 17910
rect 6585 17960 6645 18020
rect 6585 17850 6645 17910
rect 6985 17960 7045 18020
rect 6985 17850 7045 17910
rect 7385 17960 7445 18020
rect 7385 17850 7445 17910
rect 7785 17960 7845 18020
rect 7785 17850 7845 17910
rect 8185 17960 8245 18020
rect 8185 17850 8245 17910
rect 8585 17960 8645 18020
rect 8585 17850 8645 17910
rect 8985 17960 9045 18020
rect 8985 17850 9045 17910
rect 9385 17960 9445 18020
rect 9385 17850 9445 17910
rect 9785 17960 9845 18020
rect 9785 17850 9845 17910
rect 10185 17960 10245 18020
rect 10185 17850 10245 17910
rect 10585 17960 10645 18020
rect 10585 17850 10645 17910
rect 10985 17960 11045 18020
rect 10985 17850 11045 17910
rect 11385 17960 11445 18020
rect 11385 17850 11445 17910
rect 11785 17960 11845 18020
rect 11785 17850 11845 17910
rect 12185 17960 12245 18020
rect 12185 17850 12245 17910
rect 12585 17960 12645 18020
rect 12585 17850 12645 17910
rect 12985 17960 13045 18020
rect 12985 17850 13045 17910
rect -215 17590 -155 17650
rect -215 17480 -155 17540
rect 185 17590 245 17650
rect 185 17480 245 17540
rect 585 17590 645 17650
rect 585 17480 645 17540
rect 985 17590 1045 17650
rect 985 17480 1045 17540
rect 1385 17590 1445 17650
rect 1385 17480 1445 17540
rect 1785 17590 1845 17650
rect 1785 17480 1845 17540
rect 2185 17590 2245 17650
rect 2185 17480 2245 17540
rect 2585 17590 2645 17650
rect 2585 17480 2645 17540
rect 2985 17590 3045 17650
rect 2985 17480 3045 17540
rect 3385 17590 3445 17650
rect 3385 17480 3445 17540
rect 3785 17590 3845 17650
rect 3785 17480 3845 17540
rect 4185 17590 4245 17650
rect 4185 17480 4245 17540
rect 4585 17590 4645 17650
rect 4585 17480 4645 17540
rect 4985 17590 5045 17650
rect 4985 17480 5045 17540
rect 5385 17590 5445 17650
rect 5385 17480 5445 17540
rect 5785 17590 5845 17650
rect 5785 17480 5845 17540
rect 6185 17590 6245 17650
rect 6185 17480 6245 17540
rect 6585 17590 6645 17650
rect 6585 17480 6645 17540
rect 6985 17590 7045 17650
rect 6985 17480 7045 17540
rect 7385 17590 7445 17650
rect 7385 17480 7445 17540
rect 7785 17590 7845 17650
rect 7785 17480 7845 17540
rect 8185 17590 8245 17650
rect 8185 17480 8245 17540
rect 8585 17590 8645 17650
rect 8585 17480 8645 17540
rect 8985 17590 9045 17650
rect 8985 17480 9045 17540
rect 9385 17590 9445 17650
rect 9385 17480 9445 17540
rect 9785 17590 9845 17650
rect 9785 17480 9845 17540
rect 10185 17590 10245 17650
rect 10185 17480 10245 17540
rect 10585 17590 10645 17650
rect 10585 17480 10645 17540
rect 10985 17590 11045 17650
rect 10985 17480 11045 17540
rect 11385 17590 11445 17650
rect 11385 17480 11445 17540
rect 11785 17590 11845 17650
rect 11785 17480 11845 17540
rect 12185 17590 12245 17650
rect 12185 17480 12245 17540
rect 12585 17590 12645 17650
rect 12585 17480 12645 17540
rect 12985 17590 13045 17650
rect 12985 17480 13045 17540
rect -215 17220 -155 17280
rect -215 17110 -155 17170
rect 185 17220 245 17280
rect 185 17110 245 17170
rect 585 17220 645 17280
rect 585 17110 645 17170
rect 985 17220 1045 17280
rect 985 17110 1045 17170
rect 1385 17220 1445 17280
rect 1385 17110 1445 17170
rect 1785 17220 1845 17280
rect 1785 17110 1845 17170
rect 2185 17220 2245 17280
rect 2185 17110 2245 17170
rect 2585 17220 2645 17280
rect 2585 17110 2645 17170
rect 2985 17220 3045 17280
rect 2985 17110 3045 17170
rect 3385 17220 3445 17280
rect 3385 17110 3445 17170
rect 3785 17220 3845 17280
rect 3785 17110 3845 17170
rect 4185 17220 4245 17280
rect 4185 17110 4245 17170
rect 4585 17220 4645 17280
rect 4585 17110 4645 17170
rect 4985 17220 5045 17280
rect 4985 17110 5045 17170
rect 5385 17220 5445 17280
rect 5385 17110 5445 17170
rect 5785 17220 5845 17280
rect 5785 17110 5845 17170
rect 6185 17220 6245 17280
rect 6185 17110 6245 17170
rect 6585 17220 6645 17280
rect 6585 17110 6645 17170
rect 6985 17220 7045 17280
rect 6985 17110 7045 17170
rect 7385 17220 7445 17280
rect 7385 17110 7445 17170
rect 7785 17220 7845 17280
rect 7785 17110 7845 17170
rect 8185 17220 8245 17280
rect 8185 17110 8245 17170
rect 8585 17220 8645 17280
rect 8585 17110 8645 17170
rect 8985 17220 9045 17280
rect 8985 17110 9045 17170
rect 9385 17220 9445 17280
rect 9385 17110 9445 17170
rect 9785 17220 9845 17280
rect 9785 17110 9845 17170
rect 10185 17220 10245 17280
rect 10185 17110 10245 17170
rect 10585 17220 10645 17280
rect 10585 17110 10645 17170
rect 10985 17220 11045 17280
rect 10985 17110 11045 17170
rect 11385 17220 11445 17280
rect 11385 17110 11445 17170
rect 11785 17220 11845 17280
rect 11785 17110 11845 17170
rect 12185 17220 12245 17280
rect 12185 17110 12245 17170
rect 12585 17220 12645 17280
rect 12585 17110 12645 17170
rect 12985 17220 13045 17280
rect 12985 17110 13045 17170
rect -215 16850 -155 16910
rect -215 16740 -155 16800
rect 185 16850 245 16910
rect 185 16740 245 16800
rect 585 16850 645 16910
rect 585 16740 645 16800
rect 985 16850 1045 16910
rect 985 16740 1045 16800
rect 1385 16850 1445 16910
rect 1385 16740 1445 16800
rect 1785 16850 1845 16910
rect 1785 16740 1845 16800
rect 2185 16850 2245 16910
rect 2185 16740 2245 16800
rect 2585 16850 2645 16910
rect 2585 16740 2645 16800
rect 2985 16850 3045 16910
rect 2985 16740 3045 16800
rect 3385 16850 3445 16910
rect 3385 16740 3445 16800
rect 3785 16850 3845 16910
rect 3785 16740 3845 16800
rect 4185 16850 4245 16910
rect 4185 16740 4245 16800
rect 4585 16850 4645 16910
rect 4585 16740 4645 16800
rect 4985 16850 5045 16910
rect 4985 16740 5045 16800
rect 5385 16850 5445 16910
rect 5385 16740 5445 16800
rect 5785 16850 5845 16910
rect 5785 16740 5845 16800
rect 6185 16850 6245 16910
rect 6185 16740 6245 16800
rect 6585 16850 6645 16910
rect 6585 16740 6645 16800
rect 6985 16850 7045 16910
rect 6985 16740 7045 16800
rect 7385 16850 7445 16910
rect 7385 16740 7445 16800
rect 7785 16850 7845 16910
rect 7785 16740 7845 16800
rect 8185 16850 8245 16910
rect 8185 16740 8245 16800
rect 8585 16850 8645 16910
rect 8585 16740 8645 16800
rect 8985 16850 9045 16910
rect 8985 16740 9045 16800
rect 9385 16850 9445 16910
rect 9385 16740 9445 16800
rect 9785 16850 9845 16910
rect 9785 16740 9845 16800
rect 10185 16850 10245 16910
rect 10185 16740 10245 16800
rect 10585 16850 10645 16910
rect 10585 16740 10645 16800
rect 10985 16850 11045 16910
rect 10985 16740 11045 16800
rect 11385 16850 11445 16910
rect 11385 16740 11445 16800
rect 11785 16850 11845 16910
rect 11785 16740 11845 16800
rect 12185 16850 12245 16910
rect 12185 16740 12245 16800
rect 12585 16850 12645 16910
rect 12585 16740 12645 16800
rect 12985 16850 13045 16910
rect 12985 16740 13045 16800
rect -215 16480 -155 16540
rect -215 16370 -155 16430
rect 185 16480 245 16540
rect 185 16370 245 16430
rect 585 16480 645 16540
rect 585 16370 645 16430
rect 985 16480 1045 16540
rect 985 16370 1045 16430
rect 1385 16480 1445 16540
rect 1385 16370 1445 16430
rect 1785 16480 1845 16540
rect 1785 16370 1845 16430
rect 2185 16480 2245 16540
rect 2185 16370 2245 16430
rect 2585 16480 2645 16540
rect 2585 16370 2645 16430
rect 2985 16480 3045 16540
rect 2985 16370 3045 16430
rect 3385 16480 3445 16540
rect 3385 16370 3445 16430
rect 3785 16480 3845 16540
rect 3785 16370 3845 16430
rect 4185 16480 4245 16540
rect 4185 16370 4245 16430
rect 4585 16480 4645 16540
rect 4585 16370 4645 16430
rect 4985 16480 5045 16540
rect 4985 16370 5045 16430
rect 5385 16480 5445 16540
rect 5385 16370 5445 16430
rect 5785 16480 5845 16540
rect 5785 16370 5845 16430
rect 6185 16480 6245 16540
rect 6185 16370 6245 16430
rect 6585 16480 6645 16540
rect 6585 16370 6645 16430
rect 6985 16480 7045 16540
rect 6985 16370 7045 16430
rect 7385 16480 7445 16540
rect 7385 16370 7445 16430
rect 7785 16480 7845 16540
rect 7785 16370 7845 16430
rect 8185 16480 8245 16540
rect 8185 16370 8245 16430
rect 8585 16480 8645 16540
rect 8585 16370 8645 16430
rect 8985 16480 9045 16540
rect 8985 16370 9045 16430
rect 9385 16480 9445 16540
rect 9385 16370 9445 16430
rect 9785 16480 9845 16540
rect 9785 16370 9845 16430
rect 10185 16480 10245 16540
rect 10185 16370 10245 16430
rect 10585 16480 10645 16540
rect 10585 16370 10645 16430
rect 10985 16480 11045 16540
rect 10985 16370 11045 16430
rect 11385 16480 11445 16540
rect 11385 16370 11445 16430
rect 11785 16480 11845 16540
rect 11785 16370 11845 16430
rect 12185 16480 12245 16540
rect 12185 16370 12245 16430
rect 12585 16480 12645 16540
rect 12585 16370 12645 16430
rect 12985 16480 13045 16540
rect 12985 16370 13045 16430
rect -215 16110 -155 16170
rect -215 16000 -155 16060
rect 185 16110 245 16170
rect 185 16000 245 16060
rect 585 16110 645 16170
rect 585 16000 645 16060
rect 985 16110 1045 16170
rect 985 16000 1045 16060
rect 1385 16110 1445 16170
rect 1385 16000 1445 16060
rect 1785 16110 1845 16170
rect 1785 16000 1845 16060
rect 2185 16110 2245 16170
rect 2185 16000 2245 16060
rect 2585 16110 2645 16170
rect 2585 16000 2645 16060
rect 2985 16110 3045 16170
rect 2985 16000 3045 16060
rect 3385 16110 3445 16170
rect 3385 16000 3445 16060
rect 3785 16110 3845 16170
rect 3785 16000 3845 16060
rect 4185 16110 4245 16170
rect 4185 16000 4245 16060
rect 4585 16110 4645 16170
rect 4585 16000 4645 16060
rect 4985 16110 5045 16170
rect 4985 16000 5045 16060
rect 5385 16110 5445 16170
rect 5385 16000 5445 16060
rect 5785 16110 5845 16170
rect 5785 16000 5845 16060
rect 6185 16110 6245 16170
rect 6185 16000 6245 16060
rect 6585 16110 6645 16170
rect 6585 16000 6645 16060
rect 6985 16110 7045 16170
rect 6985 16000 7045 16060
rect 7385 16110 7445 16170
rect 7385 16000 7445 16060
rect 7785 16110 7845 16170
rect 7785 16000 7845 16060
rect 8185 16110 8245 16170
rect 8185 16000 8245 16060
rect 8585 16110 8645 16170
rect 8585 16000 8645 16060
rect 8985 16110 9045 16170
rect 8985 16000 9045 16060
rect 9385 16110 9445 16170
rect 9385 16000 9445 16060
rect 9785 16110 9845 16170
rect 9785 16000 9845 16060
rect 10185 16110 10245 16170
rect 10185 16000 10245 16060
rect 10585 16110 10645 16170
rect 10585 16000 10645 16060
rect 10985 16110 11045 16170
rect 10985 16000 11045 16060
rect 11385 16110 11445 16170
rect 11385 16000 11445 16060
rect 11785 16110 11845 16170
rect 11785 16000 11845 16060
rect 12185 16110 12245 16170
rect 12185 16000 12245 16060
rect 12585 16110 12645 16170
rect 12585 16000 12645 16060
rect 12985 16110 13045 16170
rect 12985 16000 13045 16060
rect -215 15740 -155 15800
rect -215 15630 -155 15690
rect 185 15740 245 15800
rect 185 15630 245 15690
rect 585 15740 645 15800
rect 585 15630 645 15690
rect 985 15740 1045 15800
rect 985 15630 1045 15690
rect 1385 15740 1445 15800
rect 1385 15630 1445 15690
rect 1785 15740 1845 15800
rect 1785 15630 1845 15690
rect 2185 15740 2245 15800
rect 2185 15630 2245 15690
rect 2585 15740 2645 15800
rect 2585 15630 2645 15690
rect 2985 15740 3045 15800
rect 2985 15630 3045 15690
rect 3385 15740 3445 15800
rect 3385 15630 3445 15690
rect 3785 15740 3845 15800
rect 3785 15630 3845 15690
rect 4185 15740 4245 15800
rect 4185 15630 4245 15690
rect 4585 15740 4645 15800
rect 4585 15630 4645 15690
rect 4985 15740 5045 15800
rect 4985 15630 5045 15690
rect 5385 15740 5445 15800
rect 5385 15630 5445 15690
rect 5785 15740 5845 15800
rect 5785 15630 5845 15690
rect 6185 15740 6245 15800
rect 6185 15630 6245 15690
rect 6585 15740 6645 15800
rect 6585 15630 6645 15690
rect 6985 15740 7045 15800
rect 6985 15630 7045 15690
rect 7385 15740 7445 15800
rect 7385 15630 7445 15690
rect 7785 15740 7845 15800
rect 7785 15630 7845 15690
rect 8185 15740 8245 15800
rect 8185 15630 8245 15690
rect 8585 15740 8645 15800
rect 8585 15630 8645 15690
rect 8985 15740 9045 15800
rect 8985 15630 9045 15690
rect 9385 15740 9445 15800
rect 9385 15630 9445 15690
rect 9785 15740 9845 15800
rect 9785 15630 9845 15690
rect 10185 15740 10245 15800
rect 10185 15630 10245 15690
rect 10585 15740 10645 15800
rect 10585 15630 10645 15690
rect 10985 15740 11045 15800
rect 10985 15630 11045 15690
rect 11385 15740 11445 15800
rect 11385 15630 11445 15690
rect 11785 15740 11845 15800
rect 11785 15630 11845 15690
rect 12185 15740 12245 15800
rect 12185 15630 12245 15690
rect 12585 15740 12645 15800
rect 12585 15630 12645 15690
rect 12985 15740 13045 15800
rect 12985 15630 13045 15690
rect -215 15370 -155 15430
rect -215 15260 -155 15320
rect 185 15370 245 15430
rect 185 15260 245 15320
rect 585 15370 645 15430
rect 585 15260 645 15320
rect 985 15370 1045 15430
rect 985 15260 1045 15320
rect 1385 15370 1445 15430
rect 1385 15260 1445 15320
rect 1785 15370 1845 15430
rect 1785 15260 1845 15320
rect 2185 15370 2245 15430
rect 2185 15260 2245 15320
rect 2585 15370 2645 15430
rect 2585 15260 2645 15320
rect 2985 15370 3045 15430
rect 2985 15260 3045 15320
rect 3385 15370 3445 15430
rect 3385 15260 3445 15320
rect 3785 15370 3845 15430
rect 3785 15260 3845 15320
rect 4185 15370 4245 15430
rect 4185 15260 4245 15320
rect 4585 15370 4645 15430
rect 4585 15260 4645 15320
rect 4985 15370 5045 15430
rect 4985 15260 5045 15320
rect 5385 15370 5445 15430
rect 5385 15260 5445 15320
rect 5785 15370 5845 15430
rect 5785 15260 5845 15320
rect 6185 15370 6245 15430
rect 6185 15260 6245 15320
rect 6585 15370 6645 15430
rect 6585 15260 6645 15320
rect 6985 15370 7045 15430
rect 6985 15260 7045 15320
rect 7385 15370 7445 15430
rect 7385 15260 7445 15320
rect 7785 15370 7845 15430
rect 7785 15260 7845 15320
rect 8185 15370 8245 15430
rect 8185 15260 8245 15320
rect 8585 15370 8645 15430
rect 8585 15260 8645 15320
rect 8985 15370 9045 15430
rect 8985 15260 9045 15320
rect 9385 15370 9445 15430
rect 9385 15260 9445 15320
rect 9785 15370 9845 15430
rect 9785 15260 9845 15320
rect 10185 15370 10245 15430
rect 10185 15260 10245 15320
rect 10585 15370 10645 15430
rect 10585 15260 10645 15320
rect 10985 15370 11045 15430
rect 10985 15260 11045 15320
rect 11385 15370 11445 15430
rect 11385 15260 11445 15320
rect 11785 15370 11845 15430
rect 11785 15260 11845 15320
rect 12185 15370 12245 15430
rect 12185 15260 12245 15320
rect 12585 15370 12645 15430
rect 12585 15260 12645 15320
rect 12985 15370 13045 15430
rect 12985 15260 13045 15320
rect -215 15000 -155 15060
rect -215 14890 -155 14950
rect 185 15000 245 15060
rect 185 14890 245 14950
rect 585 15000 645 15060
rect 585 14890 645 14950
rect 985 15000 1045 15060
rect 985 14890 1045 14950
rect 1385 15000 1445 15060
rect 1385 14890 1445 14950
rect 1785 15000 1845 15060
rect 1785 14890 1845 14950
rect 2185 15000 2245 15060
rect 2185 14890 2245 14950
rect 2585 15000 2645 15060
rect 2585 14890 2645 14950
rect 2985 15000 3045 15060
rect 2985 14890 3045 14950
rect 3385 15000 3445 15060
rect 3385 14890 3445 14950
rect 3785 15000 3845 15060
rect 3785 14890 3845 14950
rect 4185 15000 4245 15060
rect 4185 14890 4245 14950
rect 4585 15000 4645 15060
rect 4585 14890 4645 14950
rect 4985 15000 5045 15060
rect 4985 14890 5045 14950
rect 5385 15000 5445 15060
rect 5385 14890 5445 14950
rect 5785 15000 5845 15060
rect 5785 14890 5845 14950
rect 6185 15000 6245 15060
rect 6185 14890 6245 14950
rect 6585 15000 6645 15060
rect 6585 14890 6645 14950
rect 6985 15000 7045 15060
rect 6985 14890 7045 14950
rect 7385 15000 7445 15060
rect 7385 14890 7445 14950
rect 7785 15000 7845 15060
rect 7785 14890 7845 14950
rect 8185 15000 8245 15060
rect 8185 14890 8245 14950
rect 8585 15000 8645 15060
rect 8585 14890 8645 14950
rect 8985 15000 9045 15060
rect 8985 14890 9045 14950
rect 9385 15000 9445 15060
rect 9385 14890 9445 14950
rect 9785 15000 9845 15060
rect 9785 14890 9845 14950
rect 10185 15000 10245 15060
rect 10185 14890 10245 14950
rect 10585 15000 10645 15060
rect 10585 14890 10645 14950
rect 10985 15000 11045 15060
rect 10985 14890 11045 14950
rect 11385 15000 11445 15060
rect 11385 14890 11445 14950
rect 11785 15000 11845 15060
rect 11785 14890 11845 14950
rect 12185 15000 12245 15060
rect 12185 14890 12245 14950
rect 12585 15000 12645 15060
rect 12585 14890 12645 14950
rect 12985 15000 13045 15060
rect 12985 14890 13045 14950
rect -215 14630 -155 14690
rect -215 14520 -155 14580
rect 185 14630 245 14690
rect 185 14520 245 14580
rect 585 14630 645 14690
rect 585 14520 645 14580
rect 985 14630 1045 14690
rect 985 14520 1045 14580
rect 1385 14630 1445 14690
rect 1385 14520 1445 14580
rect 1785 14630 1845 14690
rect 1785 14520 1845 14580
rect 2185 14630 2245 14690
rect 2185 14520 2245 14580
rect 2585 14630 2645 14690
rect 2585 14520 2645 14580
rect 2985 14630 3045 14690
rect 2985 14520 3045 14580
rect 3385 14630 3445 14690
rect 3385 14520 3445 14580
rect 3785 14630 3845 14690
rect 3785 14520 3845 14580
rect 4185 14630 4245 14690
rect 4185 14520 4245 14580
rect 4585 14630 4645 14690
rect 4585 14520 4645 14580
rect 4985 14630 5045 14690
rect 4985 14520 5045 14580
rect 5385 14630 5445 14690
rect 5385 14520 5445 14580
rect 5785 14630 5845 14690
rect 5785 14520 5845 14580
rect 6185 14630 6245 14690
rect 6185 14520 6245 14580
rect 6585 14630 6645 14690
rect 6585 14520 6645 14580
rect 6985 14630 7045 14690
rect 6985 14520 7045 14580
rect 7385 14630 7445 14690
rect 7385 14520 7445 14580
rect 7785 14630 7845 14690
rect 7785 14520 7845 14580
rect 8185 14630 8245 14690
rect 8185 14520 8245 14580
rect 8585 14630 8645 14690
rect 8585 14520 8645 14580
rect 8985 14630 9045 14690
rect 8985 14520 9045 14580
rect 9385 14630 9445 14690
rect 9385 14520 9445 14580
rect 9785 14630 9845 14690
rect 9785 14520 9845 14580
rect 10185 14630 10245 14690
rect 10185 14520 10245 14580
rect 10585 14630 10645 14690
rect 10585 14520 10645 14580
rect 10985 14630 11045 14690
rect 10985 14520 11045 14580
rect 11385 14630 11445 14690
rect 11385 14520 11445 14580
rect 11785 14630 11845 14690
rect 11785 14520 11845 14580
rect 12185 14630 12245 14690
rect 12185 14520 12245 14580
rect 12585 14630 12645 14690
rect 12585 14520 12645 14580
rect 12985 14630 13045 14690
rect 12985 14520 13045 14580
rect -215 14260 -155 14320
rect -215 14150 -155 14210
rect 185 14260 245 14320
rect 185 14150 245 14210
rect 585 14260 645 14320
rect 585 14150 645 14210
rect 985 14260 1045 14320
rect 985 14150 1045 14210
rect 1385 14260 1445 14320
rect 1385 14150 1445 14210
rect 1785 14260 1845 14320
rect 1785 14150 1845 14210
rect 2185 14260 2245 14320
rect 2185 14150 2245 14210
rect 2585 14260 2645 14320
rect 2585 14150 2645 14210
rect 2985 14260 3045 14320
rect 2985 14150 3045 14210
rect 3385 14260 3445 14320
rect 3385 14150 3445 14210
rect 3785 14260 3845 14320
rect 3785 14150 3845 14210
rect 4185 14260 4245 14320
rect 4185 14150 4245 14210
rect 4585 14260 4645 14320
rect 4585 14150 4645 14210
rect 4985 14260 5045 14320
rect 4985 14150 5045 14210
rect 5385 14260 5445 14320
rect 5385 14150 5445 14210
rect 5785 14260 5845 14320
rect 5785 14150 5845 14210
rect 6185 14260 6245 14320
rect 6185 14150 6245 14210
rect 6585 14260 6645 14320
rect 6585 14150 6645 14210
rect 6985 14260 7045 14320
rect 6985 14150 7045 14210
rect 7385 14260 7445 14320
rect 7385 14150 7445 14210
rect 7785 14260 7845 14320
rect 7785 14150 7845 14210
rect 8185 14260 8245 14320
rect 8185 14150 8245 14210
rect 8585 14260 8645 14320
rect 8585 14150 8645 14210
rect 8985 14260 9045 14320
rect 8985 14150 9045 14210
rect 9385 14260 9445 14320
rect 9385 14150 9445 14210
rect 9785 14260 9845 14320
rect 9785 14150 9845 14210
rect 10185 14260 10245 14320
rect 10185 14150 10245 14210
rect 10585 14260 10645 14320
rect 10585 14150 10645 14210
rect 10985 14260 11045 14320
rect 10985 14150 11045 14210
rect 11385 14260 11445 14320
rect 11385 14150 11445 14210
rect 11785 14260 11845 14320
rect 11785 14150 11845 14210
rect 12185 14260 12245 14320
rect 12185 14150 12245 14210
rect 12585 14260 12645 14320
rect 12585 14150 12645 14210
rect 12985 14260 13045 14320
rect 12985 14150 13045 14210
rect -215 13890 -155 13950
rect -215 13780 -155 13840
rect 185 13890 245 13950
rect 185 13780 245 13840
rect 585 13890 645 13950
rect 585 13780 645 13840
rect 985 13890 1045 13950
rect 985 13780 1045 13840
rect 1385 13890 1445 13950
rect 1385 13780 1445 13840
rect 1785 13890 1845 13950
rect 1785 13780 1845 13840
rect 2185 13890 2245 13950
rect 2185 13780 2245 13840
rect 2585 13890 2645 13950
rect 2585 13780 2645 13840
rect 2985 13890 3045 13950
rect 2985 13780 3045 13840
rect 3385 13890 3445 13950
rect 3385 13780 3445 13840
rect 3785 13890 3845 13950
rect 3785 13780 3845 13840
rect 4185 13890 4245 13950
rect 4185 13780 4245 13840
rect 4585 13890 4645 13950
rect 4585 13780 4645 13840
rect 4985 13890 5045 13950
rect 4985 13780 5045 13840
rect 5385 13890 5445 13950
rect 5385 13780 5445 13840
rect 5785 13890 5845 13950
rect 5785 13780 5845 13840
rect 6185 13890 6245 13950
rect 6185 13780 6245 13840
rect 6585 13890 6645 13950
rect 6585 13780 6645 13840
rect 6985 13890 7045 13950
rect 6985 13780 7045 13840
rect 7385 13890 7445 13950
rect 7385 13780 7445 13840
rect 7785 13890 7845 13950
rect 7785 13780 7845 13840
rect 8185 13890 8245 13950
rect 8185 13780 8245 13840
rect 8585 13890 8645 13950
rect 8585 13780 8645 13840
rect 8985 13890 9045 13950
rect 8985 13780 9045 13840
rect 9385 13890 9445 13950
rect 9385 13780 9445 13840
rect 9785 13890 9845 13950
rect 9785 13780 9845 13840
rect 10185 13890 10245 13950
rect 10185 13780 10245 13840
rect 10585 13890 10645 13950
rect 10585 13780 10645 13840
rect 10985 13890 11045 13950
rect 10985 13780 11045 13840
rect 11385 13890 11445 13950
rect 11385 13780 11445 13840
rect 11785 13890 11845 13950
rect 11785 13780 11845 13840
rect 12185 13890 12245 13950
rect 12185 13780 12245 13840
rect 12585 13890 12645 13950
rect 12585 13780 12645 13840
rect 12985 13890 13045 13950
rect 12985 13780 13045 13840
rect -215 13520 -155 13580
rect -215 13410 -155 13470
rect 185 13520 245 13580
rect 185 13410 245 13470
rect 585 13520 645 13580
rect 585 13410 645 13470
rect 985 13520 1045 13580
rect 985 13410 1045 13470
rect 1385 13520 1445 13580
rect 1385 13410 1445 13470
rect 1785 13520 1845 13580
rect 1785 13410 1845 13470
rect 2185 13520 2245 13580
rect 2185 13410 2245 13470
rect 2585 13520 2645 13580
rect 2585 13410 2645 13470
rect 2985 13520 3045 13580
rect 2985 13410 3045 13470
rect 3385 13520 3445 13580
rect 3385 13410 3445 13470
rect 3785 13520 3845 13580
rect 3785 13410 3845 13470
rect 4185 13520 4245 13580
rect 4185 13410 4245 13470
rect 4585 13520 4645 13580
rect 4585 13410 4645 13470
rect 4985 13520 5045 13580
rect 4985 13410 5045 13470
rect 5385 13520 5445 13580
rect 5385 13410 5445 13470
rect 5785 13520 5845 13580
rect 5785 13410 5845 13470
rect 6185 13520 6245 13580
rect 6185 13410 6245 13470
rect 6585 13520 6645 13580
rect 6585 13410 6645 13470
rect 6985 13520 7045 13580
rect 6985 13410 7045 13470
rect 7385 13520 7445 13580
rect 7385 13410 7445 13470
rect 7785 13520 7845 13580
rect 7785 13410 7845 13470
rect 8185 13520 8245 13580
rect 8185 13410 8245 13470
rect 8585 13520 8645 13580
rect 8585 13410 8645 13470
rect 8985 13520 9045 13580
rect 8985 13410 9045 13470
rect 9385 13520 9445 13580
rect 9385 13410 9445 13470
rect 9785 13520 9845 13580
rect 9785 13410 9845 13470
rect 10185 13520 10245 13580
rect 10185 13410 10245 13470
rect 10585 13520 10645 13580
rect 10585 13410 10645 13470
rect 10985 13520 11045 13580
rect 10985 13410 11045 13470
rect 11385 13520 11445 13580
rect 11385 13410 11445 13470
rect 11785 13520 11845 13580
rect 11785 13410 11845 13470
rect 12185 13520 12245 13580
rect 12185 13410 12245 13470
rect 12585 13520 12645 13580
rect 12585 13410 12645 13470
rect 12985 13520 13045 13580
rect 12985 13410 13045 13470
rect -215 13150 -155 13210
rect -215 13040 -155 13100
rect 185 13150 245 13210
rect 185 13040 245 13100
rect 585 13150 645 13210
rect 585 13040 645 13100
rect 985 13150 1045 13210
rect 985 13040 1045 13100
rect 1385 13150 1445 13210
rect 1385 13040 1445 13100
rect 1785 13150 1845 13210
rect 1785 13040 1845 13100
rect 2185 13150 2245 13210
rect 2185 13040 2245 13100
rect 2585 13150 2645 13210
rect 2585 13040 2645 13100
rect 2985 13150 3045 13210
rect 2985 13040 3045 13100
rect 3385 13150 3445 13210
rect 3385 13040 3445 13100
rect 3785 13150 3845 13210
rect 3785 13040 3845 13100
rect 4185 13150 4245 13210
rect 4185 13040 4245 13100
rect 4585 13150 4645 13210
rect 4585 13040 4645 13100
rect 4985 13150 5045 13210
rect 4985 13040 5045 13100
rect 5385 13150 5445 13210
rect 5385 13040 5445 13100
rect 5785 13150 5845 13210
rect 5785 13040 5845 13100
rect 6185 13150 6245 13210
rect 6185 13040 6245 13100
rect 6585 13150 6645 13210
rect 6585 13040 6645 13100
rect 6985 13150 7045 13210
rect 6985 13040 7045 13100
rect 7385 13150 7445 13210
rect 7385 13040 7445 13100
rect 7785 13150 7845 13210
rect 7785 13040 7845 13100
rect 8185 13150 8245 13210
rect 8185 13040 8245 13100
rect 8585 13150 8645 13210
rect 8585 13040 8645 13100
rect 8985 13150 9045 13210
rect 8985 13040 9045 13100
rect 9385 13150 9445 13210
rect 9385 13040 9445 13100
rect 9785 13150 9845 13210
rect 9785 13040 9845 13100
rect 10185 13150 10245 13210
rect 10185 13040 10245 13100
rect 10585 13150 10645 13210
rect 10585 13040 10645 13100
rect 10985 13150 11045 13210
rect 10985 13040 11045 13100
rect 11385 13150 11445 13210
rect 11385 13040 11445 13100
rect 11785 13150 11845 13210
rect 11785 13040 11845 13100
rect 12185 13150 12245 13210
rect 12185 13040 12245 13100
rect 12585 13150 12645 13210
rect 12585 13040 12645 13100
rect 12985 13150 13045 13210
rect 12985 13040 13045 13100
rect -215 12780 -155 12840
rect -215 12670 -155 12730
rect 185 12780 245 12840
rect 185 12670 245 12730
rect 585 12780 645 12840
rect 585 12670 645 12730
rect 985 12780 1045 12840
rect 985 12670 1045 12730
rect 1385 12780 1445 12840
rect 1385 12670 1445 12730
rect 1785 12780 1845 12840
rect 1785 12670 1845 12730
rect 2185 12780 2245 12840
rect 2185 12670 2245 12730
rect 2585 12780 2645 12840
rect 2585 12670 2645 12730
rect 2985 12780 3045 12840
rect 2985 12670 3045 12730
rect 3385 12780 3445 12840
rect 3385 12670 3445 12730
rect 3785 12780 3845 12840
rect 3785 12670 3845 12730
rect 4185 12780 4245 12840
rect 4185 12670 4245 12730
rect 4585 12780 4645 12840
rect 4585 12670 4645 12730
rect 4985 12780 5045 12840
rect 4985 12670 5045 12730
rect 5385 12780 5445 12840
rect 5385 12670 5445 12730
rect 5785 12780 5845 12840
rect 5785 12670 5845 12730
rect 6185 12780 6245 12840
rect 6185 12670 6245 12730
rect 6585 12780 6645 12840
rect 6585 12670 6645 12730
rect 6985 12780 7045 12840
rect 6985 12670 7045 12730
rect 7385 12780 7445 12840
rect 7385 12670 7445 12730
rect 7785 12780 7845 12840
rect 7785 12670 7845 12730
rect 8185 12780 8245 12840
rect 8185 12670 8245 12730
rect 8585 12780 8645 12840
rect 8585 12670 8645 12730
rect 8985 12780 9045 12840
rect 8985 12670 9045 12730
rect 9385 12780 9445 12840
rect 9385 12670 9445 12730
rect 9785 12780 9845 12840
rect 9785 12670 9845 12730
rect 10185 12780 10245 12840
rect 10185 12670 10245 12730
rect 10585 12780 10645 12840
rect 10585 12670 10645 12730
rect 10985 12780 11045 12840
rect 10985 12670 11045 12730
rect 11385 12780 11445 12840
rect 11385 12670 11445 12730
rect 11785 12780 11845 12840
rect 11785 12670 11845 12730
rect 12185 12780 12245 12840
rect 12185 12670 12245 12730
rect 12585 12780 12645 12840
rect 12585 12670 12645 12730
rect 12985 12780 13045 12840
rect 12985 12670 13045 12730
rect -215 12410 -155 12470
rect -215 12300 -155 12360
rect 185 12410 245 12470
rect 185 12300 245 12360
rect 585 12410 645 12470
rect 585 12300 645 12360
rect 985 12410 1045 12470
rect 985 12300 1045 12360
rect 1385 12410 1445 12470
rect 1385 12300 1445 12360
rect 1785 12410 1845 12470
rect 1785 12300 1845 12360
rect 2185 12410 2245 12470
rect 2185 12300 2245 12360
rect 2585 12410 2645 12470
rect 2585 12300 2645 12360
rect 2985 12410 3045 12470
rect 2985 12300 3045 12360
rect 3385 12410 3445 12470
rect 3385 12300 3445 12360
rect 3785 12410 3845 12470
rect 3785 12300 3845 12360
rect 4185 12410 4245 12470
rect 4185 12300 4245 12360
rect 4585 12410 4645 12470
rect 4585 12300 4645 12360
rect 4985 12410 5045 12470
rect 4985 12300 5045 12360
rect 5385 12410 5445 12470
rect 5385 12300 5445 12360
rect 5785 12410 5845 12470
rect 5785 12300 5845 12360
rect 6185 12410 6245 12470
rect 6185 12300 6245 12360
rect 6585 12410 6645 12470
rect 6585 12300 6645 12360
rect 6985 12410 7045 12470
rect 6985 12300 7045 12360
rect 7385 12410 7445 12470
rect 7385 12300 7445 12360
rect 7785 12410 7845 12470
rect 7785 12300 7845 12360
rect 8185 12410 8245 12470
rect 8185 12300 8245 12360
rect 8585 12410 8645 12470
rect 8585 12300 8645 12360
rect 8985 12410 9045 12470
rect 8985 12300 9045 12360
rect 9385 12410 9445 12470
rect 9385 12300 9445 12360
rect 9785 12410 9845 12470
rect 9785 12300 9845 12360
rect 10185 12410 10245 12470
rect 10185 12300 10245 12360
rect 10585 12410 10645 12470
rect 10585 12300 10645 12360
rect 10985 12410 11045 12470
rect 10985 12300 11045 12360
rect 11385 12410 11445 12470
rect 11385 12300 11445 12360
rect 11785 12410 11845 12470
rect 11785 12300 11845 12360
rect 12185 12410 12245 12470
rect 12185 12300 12245 12360
rect 12585 12410 12645 12470
rect 12585 12300 12645 12360
rect 12985 12410 13045 12470
rect 12985 12300 13045 12360
rect -215 12040 -155 12100
rect -215 11930 -155 11990
rect 185 12040 245 12100
rect 185 11930 245 11990
rect 585 12040 645 12100
rect 585 11930 645 11990
rect 985 12040 1045 12100
rect 985 11930 1045 11990
rect 1385 12040 1445 12100
rect 1385 11930 1445 11990
rect 1785 12040 1845 12100
rect 1785 11930 1845 11990
rect 2185 12040 2245 12100
rect 2185 11930 2245 11990
rect 2585 12040 2645 12100
rect 2585 11930 2645 11990
rect 2985 12040 3045 12100
rect 2985 11930 3045 11990
rect 3385 12040 3445 12100
rect 3385 11930 3445 11990
rect 3785 12040 3845 12100
rect 3785 11930 3845 11990
rect 4185 12040 4245 12100
rect 4185 11930 4245 11990
rect 4585 12040 4645 12100
rect 4585 11930 4645 11990
rect 4985 12040 5045 12100
rect 4985 11930 5045 11990
rect 5385 12040 5445 12100
rect 5385 11930 5445 11990
rect 5785 12040 5845 12100
rect 5785 11930 5845 11990
rect 6185 12040 6245 12100
rect 6185 11930 6245 11990
rect 6585 12040 6645 12100
rect 6585 11930 6645 11990
rect 6985 12040 7045 12100
rect 6985 11930 7045 11990
rect 7385 12040 7445 12100
rect 7385 11930 7445 11990
rect 7785 12040 7845 12100
rect 7785 11930 7845 11990
rect 8185 12040 8245 12100
rect 8185 11930 8245 11990
rect 8585 12040 8645 12100
rect 8585 11930 8645 11990
rect 8985 12040 9045 12100
rect 8985 11930 9045 11990
rect 9385 12040 9445 12100
rect 9385 11930 9445 11990
rect 9785 12040 9845 12100
rect 9785 11930 9845 11990
rect 10185 12040 10245 12100
rect 10185 11930 10245 11990
rect 10585 12040 10645 12100
rect 10585 11930 10645 11990
rect 10985 12040 11045 12100
rect 10985 11930 11045 11990
rect 11385 12040 11445 12100
rect 11385 11930 11445 11990
rect 11785 12040 11845 12100
rect 11785 11930 11845 11990
rect 12185 12040 12245 12100
rect 12185 11930 12245 11990
rect 12585 12040 12645 12100
rect 12585 11930 12645 11990
rect 12985 12040 13045 12100
rect 12985 11930 13045 11990
rect -215 11670 -155 11730
rect -215 11560 -155 11620
rect 185 11670 245 11730
rect 185 11560 245 11620
rect 585 11670 645 11730
rect 585 11560 645 11620
rect 985 11670 1045 11730
rect 985 11560 1045 11620
rect 1385 11670 1445 11730
rect 1385 11560 1445 11620
rect 1785 11670 1845 11730
rect 1785 11560 1845 11620
rect 2185 11670 2245 11730
rect 2185 11560 2245 11620
rect 2585 11670 2645 11730
rect 2585 11560 2645 11620
rect 2985 11670 3045 11730
rect 2985 11560 3045 11620
rect 3385 11670 3445 11730
rect 3385 11560 3445 11620
rect 3785 11670 3845 11730
rect 3785 11560 3845 11620
rect 4185 11670 4245 11730
rect 4185 11560 4245 11620
rect 4585 11670 4645 11730
rect 4585 11560 4645 11620
rect 4985 11670 5045 11730
rect 4985 11560 5045 11620
rect 5385 11670 5445 11730
rect 5385 11560 5445 11620
rect 5785 11670 5845 11730
rect 5785 11560 5845 11620
rect 6185 11670 6245 11730
rect 6185 11560 6245 11620
rect 6585 11670 6645 11730
rect 6585 11560 6645 11620
rect 6985 11670 7045 11730
rect 6985 11560 7045 11620
rect 7385 11670 7445 11730
rect 7385 11560 7445 11620
rect 7785 11670 7845 11730
rect 7785 11560 7845 11620
rect 8185 11670 8245 11730
rect 8185 11560 8245 11620
rect 8585 11670 8645 11730
rect 8585 11560 8645 11620
rect 8985 11670 9045 11730
rect 8985 11560 9045 11620
rect 9385 11670 9445 11730
rect 9385 11560 9445 11620
rect 9785 11670 9845 11730
rect 9785 11560 9845 11620
rect 10185 11670 10245 11730
rect 10185 11560 10245 11620
rect 10585 11670 10645 11730
rect 10585 11560 10645 11620
rect 10985 11670 11045 11730
rect 10985 11560 11045 11620
rect 11385 11670 11445 11730
rect 11385 11560 11445 11620
rect 11785 11670 11845 11730
rect 11785 11560 11845 11620
rect 12185 11670 12245 11730
rect 12185 11560 12245 11620
rect 12585 11670 12645 11730
rect 12585 11560 12645 11620
rect 12985 11670 13045 11730
rect 12985 11560 13045 11620
rect -215 11300 -155 11360
rect -215 11190 -155 11250
rect 185 11300 245 11360
rect 185 11190 245 11250
rect 585 11300 645 11360
rect 585 11190 645 11250
rect 985 11300 1045 11360
rect 985 11190 1045 11250
rect 1385 11300 1445 11360
rect 1385 11190 1445 11250
rect 1785 11300 1845 11360
rect 1785 11190 1845 11250
rect 2185 11300 2245 11360
rect 2185 11190 2245 11250
rect 2585 11300 2645 11360
rect 2585 11190 2645 11250
rect 2985 11300 3045 11360
rect 2985 11190 3045 11250
rect 3385 11300 3445 11360
rect 3385 11190 3445 11250
rect 3785 11300 3845 11360
rect 3785 11190 3845 11250
rect 4185 11300 4245 11360
rect 4185 11190 4245 11250
rect 4585 11300 4645 11360
rect 4585 11190 4645 11250
rect 4985 11300 5045 11360
rect 4985 11190 5045 11250
rect 5385 11300 5445 11360
rect 5385 11190 5445 11250
rect 5785 11300 5845 11360
rect 5785 11190 5845 11250
rect 6185 11300 6245 11360
rect 6185 11190 6245 11250
rect 6585 11300 6645 11360
rect 6585 11190 6645 11250
rect 6985 11300 7045 11360
rect 6985 11190 7045 11250
rect 7385 11300 7445 11360
rect 7385 11190 7445 11250
rect 7785 11300 7845 11360
rect 7785 11190 7845 11250
rect 8185 11300 8245 11360
rect 8185 11190 8245 11250
rect 8585 11300 8645 11360
rect 8585 11190 8645 11250
rect 8985 11300 9045 11360
rect 8985 11190 9045 11250
rect 9385 11300 9445 11360
rect 9385 11190 9445 11250
rect 9785 11300 9845 11360
rect 9785 11190 9845 11250
rect 10185 11300 10245 11360
rect 10185 11190 10245 11250
rect 10585 11300 10645 11360
rect 10585 11190 10645 11250
rect 10985 11300 11045 11360
rect 10985 11190 11045 11250
rect 11385 11300 11445 11360
rect 11385 11190 11445 11250
rect 11785 11300 11845 11360
rect 11785 11190 11845 11250
rect 12185 11300 12245 11360
rect 12185 11190 12245 11250
rect 12585 11300 12645 11360
rect 12585 11190 12645 11250
rect 12985 11300 13045 11360
rect 12985 11190 13045 11250
rect -215 10930 -155 10990
rect -215 10820 -155 10880
rect 185 10930 245 10990
rect 185 10820 245 10880
rect 585 10930 645 10990
rect 585 10820 645 10880
rect 985 10930 1045 10990
rect 985 10820 1045 10880
rect 1385 10930 1445 10990
rect 1385 10820 1445 10880
rect 1785 10930 1845 10990
rect 1785 10820 1845 10880
rect 2185 10930 2245 10990
rect 2185 10820 2245 10880
rect 2585 10930 2645 10990
rect 2585 10820 2645 10880
rect 2985 10930 3045 10990
rect 2985 10820 3045 10880
rect 3385 10930 3445 10990
rect 3385 10820 3445 10880
rect 3785 10930 3845 10990
rect 3785 10820 3845 10880
rect 4185 10930 4245 10990
rect 4185 10820 4245 10880
rect 4585 10930 4645 10990
rect 4585 10820 4645 10880
rect 4985 10930 5045 10990
rect 4985 10820 5045 10880
rect 5385 10930 5445 10990
rect 5385 10820 5445 10880
rect 5785 10930 5845 10990
rect 5785 10820 5845 10880
rect 6185 10930 6245 10990
rect 6185 10820 6245 10880
rect 6585 10930 6645 10990
rect 6585 10820 6645 10880
rect 6985 10930 7045 10990
rect 6985 10820 7045 10880
rect 7385 10930 7445 10990
rect 7385 10820 7445 10880
rect 7785 10930 7845 10990
rect 7785 10820 7845 10880
rect 8185 10930 8245 10990
rect 8185 10820 8245 10880
rect 8585 10930 8645 10990
rect 8585 10820 8645 10880
rect 8985 10930 9045 10990
rect 8985 10820 9045 10880
rect 9385 10930 9445 10990
rect 9385 10820 9445 10880
rect 9785 10930 9845 10990
rect 9785 10820 9845 10880
rect 10185 10930 10245 10990
rect 10185 10820 10245 10880
rect 10585 10930 10645 10990
rect 10585 10820 10645 10880
rect 10985 10930 11045 10990
rect 10985 10820 11045 10880
rect 11385 10930 11445 10990
rect 11385 10820 11445 10880
rect 11785 10930 11845 10990
rect 11785 10820 11845 10880
rect 12185 10930 12245 10990
rect 12185 10820 12245 10880
rect 12585 10930 12645 10990
rect 12585 10820 12645 10880
rect 12985 10930 13045 10990
rect 12985 10820 13045 10880
rect -215 10560 -155 10620
rect -215 10450 -155 10510
rect 185 10560 245 10620
rect 185 10450 245 10510
rect 585 10560 645 10620
rect 585 10450 645 10510
rect 985 10560 1045 10620
rect 985 10450 1045 10510
rect 1385 10560 1445 10620
rect 1385 10450 1445 10510
rect 1785 10560 1845 10620
rect 1785 10450 1845 10510
rect 2185 10560 2245 10620
rect 2185 10450 2245 10510
rect 2585 10560 2645 10620
rect 2585 10450 2645 10510
rect 2985 10560 3045 10620
rect 2985 10450 3045 10510
rect 3385 10560 3445 10620
rect 3385 10450 3445 10510
rect 3785 10560 3845 10620
rect 3785 10450 3845 10510
rect 4185 10560 4245 10620
rect 4185 10450 4245 10510
rect 4585 10560 4645 10620
rect 4585 10450 4645 10510
rect 4985 10560 5045 10620
rect 4985 10450 5045 10510
rect 5385 10560 5445 10620
rect 5385 10450 5445 10510
rect 5785 10560 5845 10620
rect 5785 10450 5845 10510
rect 6185 10560 6245 10620
rect 6185 10450 6245 10510
rect 6585 10560 6645 10620
rect 6585 10450 6645 10510
rect 6985 10560 7045 10620
rect 6985 10450 7045 10510
rect 7385 10560 7445 10620
rect 7385 10450 7445 10510
rect 7785 10560 7845 10620
rect 7785 10450 7845 10510
rect 8185 10560 8245 10620
rect 8185 10450 8245 10510
rect 8585 10560 8645 10620
rect 8585 10450 8645 10510
rect 8985 10560 9045 10620
rect 8985 10450 9045 10510
rect 9385 10560 9445 10620
rect 9385 10450 9445 10510
rect 9785 10560 9845 10620
rect 9785 10450 9845 10510
rect 10185 10560 10245 10620
rect 10185 10450 10245 10510
rect 10585 10560 10645 10620
rect 10585 10450 10645 10510
rect 10985 10560 11045 10620
rect 10985 10450 11045 10510
rect 11385 10560 11445 10620
rect 11385 10450 11445 10510
rect 11785 10560 11845 10620
rect 11785 10450 11845 10510
rect 12185 10560 12245 10620
rect 12185 10450 12245 10510
rect 12585 10560 12645 10620
rect 12585 10450 12645 10510
rect 12985 10560 13045 10620
rect 12985 10450 13045 10510
rect -215 10190 -155 10250
rect -215 10080 -155 10140
rect 185 10190 245 10250
rect 185 10080 245 10140
rect 585 10190 645 10250
rect 585 10080 645 10140
rect 985 10190 1045 10250
rect 985 10080 1045 10140
rect 1385 10190 1445 10250
rect 1385 10080 1445 10140
rect 1785 10190 1845 10250
rect 1785 10080 1845 10140
rect 2185 10190 2245 10250
rect 2185 10080 2245 10140
rect 2585 10190 2645 10250
rect 2585 10080 2645 10140
rect 2985 10190 3045 10250
rect 2985 10080 3045 10140
rect 3385 10190 3445 10250
rect 3385 10080 3445 10140
rect 3785 10190 3845 10250
rect 3785 10080 3845 10140
rect 4185 10190 4245 10250
rect 4185 10080 4245 10140
rect 4585 10190 4645 10250
rect 4585 10080 4645 10140
rect 4985 10190 5045 10250
rect 4985 10080 5045 10140
rect 5385 10190 5445 10250
rect 5385 10080 5445 10140
rect 5785 10190 5845 10250
rect 5785 10080 5845 10140
rect 6185 10190 6245 10250
rect 6185 10080 6245 10140
rect 6585 10190 6645 10250
rect 6585 10080 6645 10140
rect 6985 10190 7045 10250
rect 6985 10080 7045 10140
rect 7385 10190 7445 10250
rect 7385 10080 7445 10140
rect 7785 10190 7845 10250
rect 7785 10080 7845 10140
rect 8185 10190 8245 10250
rect 8185 10080 8245 10140
rect 8585 10190 8645 10250
rect 8585 10080 8645 10140
rect 8985 10190 9045 10250
rect 8985 10080 9045 10140
rect 9385 10190 9445 10250
rect 9385 10080 9445 10140
rect 9785 10190 9845 10250
rect 9785 10080 9845 10140
rect 10185 10190 10245 10250
rect 10185 10080 10245 10140
rect 10585 10190 10645 10250
rect 10585 10080 10645 10140
rect 10985 10190 11045 10250
rect 10985 10080 11045 10140
rect 11385 10190 11445 10250
rect 11385 10080 11445 10140
rect 11785 10190 11845 10250
rect 11785 10080 11845 10140
rect 12185 10190 12245 10250
rect 12185 10080 12245 10140
rect 12585 10190 12645 10250
rect 12585 10080 12645 10140
rect 12985 10190 13045 10250
rect 12985 10080 13045 10140
rect -215 9820 -155 9880
rect -215 9710 -155 9770
rect 185 9820 245 9880
rect 185 9710 245 9770
rect 585 9820 645 9880
rect 585 9710 645 9770
rect 985 9820 1045 9880
rect 985 9710 1045 9770
rect 1385 9820 1445 9880
rect 1385 9710 1445 9770
rect 1785 9820 1845 9880
rect 1785 9710 1845 9770
rect 2185 9820 2245 9880
rect 2185 9710 2245 9770
rect 2585 9820 2645 9880
rect 2585 9710 2645 9770
rect 2985 9820 3045 9880
rect 2985 9710 3045 9770
rect 3385 9820 3445 9880
rect 3385 9710 3445 9770
rect 3785 9820 3845 9880
rect 3785 9710 3845 9770
rect 4185 9820 4245 9880
rect 4185 9710 4245 9770
rect 4585 9820 4645 9880
rect 4585 9710 4645 9770
rect 4985 9820 5045 9880
rect 4985 9710 5045 9770
rect 5385 9820 5445 9880
rect 5385 9710 5445 9770
rect 5785 9820 5845 9880
rect 5785 9710 5845 9770
rect 6185 9820 6245 9880
rect 6185 9710 6245 9770
rect 6585 9820 6645 9880
rect 6585 9710 6645 9770
rect 6985 9820 7045 9880
rect 6985 9710 7045 9770
rect 7385 9820 7445 9880
rect 7385 9710 7445 9770
rect 7785 9820 7845 9880
rect 7785 9710 7845 9770
rect 8185 9820 8245 9880
rect 8185 9710 8245 9770
rect 8585 9820 8645 9880
rect 8585 9710 8645 9770
rect 8985 9820 9045 9880
rect 8985 9710 9045 9770
rect 9385 9820 9445 9880
rect 9385 9710 9445 9770
rect 9785 9820 9845 9880
rect 9785 9710 9845 9770
rect 10185 9820 10245 9880
rect 10185 9710 10245 9770
rect 10585 9820 10645 9880
rect 10585 9710 10645 9770
rect 10985 9820 11045 9880
rect 10985 9710 11045 9770
rect 11385 9820 11445 9880
rect 11385 9710 11445 9770
rect 11785 9820 11845 9880
rect 11785 9710 11845 9770
rect 12185 9820 12245 9880
rect 12185 9710 12245 9770
rect 12585 9820 12645 9880
rect 12585 9710 12645 9770
rect 12985 9820 13045 9880
rect 12985 9710 13045 9770
rect -215 9450 -155 9510
rect -215 9340 -155 9400
rect 185 9450 245 9510
rect 185 9340 245 9400
rect 585 9450 645 9510
rect 585 9340 645 9400
rect 985 9450 1045 9510
rect 985 9340 1045 9400
rect 1385 9450 1445 9510
rect 1385 9340 1445 9400
rect 1785 9450 1845 9510
rect 1785 9340 1845 9400
rect 2185 9450 2245 9510
rect 2185 9340 2245 9400
rect 2585 9450 2645 9510
rect 2585 9340 2645 9400
rect 2985 9450 3045 9510
rect 2985 9340 3045 9400
rect 3385 9450 3445 9510
rect 3385 9340 3445 9400
rect 3785 9450 3845 9510
rect 3785 9340 3845 9400
rect 4185 9450 4245 9510
rect 4185 9340 4245 9400
rect 4585 9450 4645 9510
rect 4585 9340 4645 9400
rect 4985 9450 5045 9510
rect 4985 9340 5045 9400
rect 5385 9450 5445 9510
rect 5385 9340 5445 9400
rect 5785 9450 5845 9510
rect 5785 9340 5845 9400
rect 6185 9450 6245 9510
rect 6185 9340 6245 9400
rect 6585 9450 6645 9510
rect 6585 9340 6645 9400
rect 6985 9450 7045 9510
rect 6985 9340 7045 9400
rect 7385 9450 7445 9510
rect 7385 9340 7445 9400
rect 7785 9450 7845 9510
rect 7785 9340 7845 9400
rect 8185 9450 8245 9510
rect 8185 9340 8245 9400
rect 8585 9450 8645 9510
rect 8585 9340 8645 9400
rect 8985 9450 9045 9510
rect 8985 9340 9045 9400
rect 9385 9450 9445 9510
rect 9385 9340 9445 9400
rect 9785 9450 9845 9510
rect 9785 9340 9845 9400
rect 10185 9450 10245 9510
rect 10185 9340 10245 9400
rect 10585 9450 10645 9510
rect 10585 9340 10645 9400
rect 10985 9450 11045 9510
rect 10985 9340 11045 9400
rect 11385 9450 11445 9510
rect 11385 9340 11445 9400
rect 11785 9450 11845 9510
rect 11785 9340 11845 9400
rect 12185 9450 12245 9510
rect 12185 9340 12245 9400
rect 12585 9450 12645 9510
rect 12585 9340 12645 9400
rect 12985 9450 13045 9510
rect 12985 9340 13045 9400
rect -215 9080 -155 9140
rect -215 8970 -155 9030
rect 185 9080 245 9140
rect 185 8970 245 9030
rect 585 9080 645 9140
rect 585 8970 645 9030
rect 985 9080 1045 9140
rect 985 8970 1045 9030
rect 1385 9080 1445 9140
rect 1385 8970 1445 9030
rect 1785 9080 1845 9140
rect 1785 8970 1845 9030
rect 2185 9080 2245 9140
rect 2185 8970 2245 9030
rect 2585 9080 2645 9140
rect 2585 8970 2645 9030
rect 2985 9080 3045 9140
rect 2985 8970 3045 9030
rect 3385 9080 3445 9140
rect 3385 8970 3445 9030
rect 3785 9080 3845 9140
rect 3785 8970 3845 9030
rect 4185 9080 4245 9140
rect 4185 8970 4245 9030
rect 4585 9080 4645 9140
rect 4585 8970 4645 9030
rect 4985 9080 5045 9140
rect 4985 8970 5045 9030
rect 5385 9080 5445 9140
rect 5385 8970 5445 9030
rect 5785 9080 5845 9140
rect 5785 8970 5845 9030
rect 6185 9080 6245 9140
rect 6185 8970 6245 9030
rect 6585 9080 6645 9140
rect 6585 8970 6645 9030
rect 6985 9080 7045 9140
rect 6985 8970 7045 9030
rect 7385 9080 7445 9140
rect 7385 8970 7445 9030
rect 7785 9080 7845 9140
rect 7785 8970 7845 9030
rect 8185 9080 8245 9140
rect 8185 8970 8245 9030
rect 8585 9080 8645 9140
rect 8585 8970 8645 9030
rect 8985 9080 9045 9140
rect 8985 8970 9045 9030
rect 9385 9080 9445 9140
rect 9385 8970 9445 9030
rect 9785 9080 9845 9140
rect 9785 8970 9845 9030
rect 10185 9080 10245 9140
rect 10185 8970 10245 9030
rect 10585 9080 10645 9140
rect 10585 8970 10645 9030
rect 10985 9080 11045 9140
rect 10985 8970 11045 9030
rect 11385 9080 11445 9140
rect 11385 8970 11445 9030
rect 11785 9080 11845 9140
rect 11785 8970 11845 9030
rect 12185 9080 12245 9140
rect 12185 8970 12245 9030
rect 12585 9080 12645 9140
rect 12585 8970 12645 9030
rect 12985 9080 13045 9140
rect 12985 8970 13045 9030
rect -215 8710 -155 8770
rect -215 8600 -155 8660
rect 185 8710 245 8770
rect 185 8600 245 8660
rect 585 8710 645 8770
rect 585 8600 645 8660
rect 985 8710 1045 8770
rect 985 8600 1045 8660
rect 1385 8710 1445 8770
rect 1385 8600 1445 8660
rect 1785 8710 1845 8770
rect 1785 8600 1845 8660
rect 2185 8710 2245 8770
rect 2185 8600 2245 8660
rect 2585 8710 2645 8770
rect 2585 8600 2645 8660
rect 2985 8710 3045 8770
rect 2985 8600 3045 8660
rect 3385 8710 3445 8770
rect 3385 8600 3445 8660
rect 3785 8710 3845 8770
rect 3785 8600 3845 8660
rect 4185 8710 4245 8770
rect 4185 8600 4245 8660
rect 4585 8710 4645 8770
rect 4585 8600 4645 8660
rect 4985 8710 5045 8770
rect 4985 8600 5045 8660
rect 5385 8710 5445 8770
rect 5385 8600 5445 8660
rect 5785 8710 5845 8770
rect 5785 8600 5845 8660
rect 6185 8710 6245 8770
rect 6185 8600 6245 8660
rect 6585 8710 6645 8770
rect 6585 8600 6645 8660
rect 6985 8710 7045 8770
rect 6985 8600 7045 8660
rect 7385 8710 7445 8770
rect 7385 8600 7445 8660
rect 7785 8710 7845 8770
rect 7785 8600 7845 8660
rect 8185 8710 8245 8770
rect 8185 8600 8245 8660
rect 8585 8710 8645 8770
rect 8585 8600 8645 8660
rect 8985 8710 9045 8770
rect 8985 8600 9045 8660
rect 9385 8710 9445 8770
rect 9385 8600 9445 8660
rect 9785 8710 9845 8770
rect 9785 8600 9845 8660
rect 10185 8710 10245 8770
rect 10185 8600 10245 8660
rect 10585 8710 10645 8770
rect 10585 8600 10645 8660
rect 10985 8710 11045 8770
rect 10985 8600 11045 8660
rect 11385 8710 11445 8770
rect 11385 8600 11445 8660
rect 11785 8710 11845 8770
rect 11785 8600 11845 8660
rect 12185 8710 12245 8770
rect 12185 8600 12245 8660
rect 12585 8710 12645 8770
rect 12585 8600 12645 8660
rect 12985 8710 13045 8770
rect 12985 8600 13045 8660
rect -215 8340 -155 8400
rect -215 8230 -155 8290
rect 185 8340 245 8400
rect 185 8230 245 8290
rect 585 8340 645 8400
rect 585 8230 645 8290
rect 985 8340 1045 8400
rect 985 8230 1045 8290
rect 1385 8340 1445 8400
rect 1385 8230 1445 8290
rect 1785 8340 1845 8400
rect 1785 8230 1845 8290
rect 2185 8340 2245 8400
rect 2185 8230 2245 8290
rect 2585 8340 2645 8400
rect 2585 8230 2645 8290
rect 2985 8340 3045 8400
rect 2985 8230 3045 8290
rect 3385 8340 3445 8400
rect 3385 8230 3445 8290
rect 3785 8340 3845 8400
rect 3785 8230 3845 8290
rect 4185 8340 4245 8400
rect 4185 8230 4245 8290
rect 4585 8340 4645 8400
rect 4585 8230 4645 8290
rect 4985 8340 5045 8400
rect 4985 8230 5045 8290
rect 5385 8340 5445 8400
rect 5385 8230 5445 8290
rect 5785 8340 5845 8400
rect 5785 8230 5845 8290
rect 6185 8340 6245 8400
rect 6185 8230 6245 8290
rect 6585 8340 6645 8400
rect 6585 8230 6645 8290
rect 6985 8340 7045 8400
rect 6985 8230 7045 8290
rect 7385 8340 7445 8400
rect 7385 8230 7445 8290
rect 7785 8340 7845 8400
rect 7785 8230 7845 8290
rect 8185 8340 8245 8400
rect 8185 8230 8245 8290
rect 8585 8340 8645 8400
rect 8585 8230 8645 8290
rect 8985 8340 9045 8400
rect 8985 8230 9045 8290
rect 9385 8340 9445 8400
rect 9385 8230 9445 8290
rect 9785 8340 9845 8400
rect 9785 8230 9845 8290
rect 10185 8340 10245 8400
rect 10185 8230 10245 8290
rect 10585 8340 10645 8400
rect 10585 8230 10645 8290
rect 10985 8340 11045 8400
rect 10985 8230 11045 8290
rect 11385 8340 11445 8400
rect 11385 8230 11445 8290
rect 11785 8340 11845 8400
rect 11785 8230 11845 8290
rect 12185 8340 12245 8400
rect 12185 8230 12245 8290
rect 12585 8340 12645 8400
rect 12585 8230 12645 8290
rect 12985 8340 13045 8400
rect 12985 8230 13045 8290
rect -215 7970 -155 8030
rect -215 7860 -155 7920
rect 185 7970 245 8030
rect 185 7860 245 7920
rect 585 7970 645 8030
rect 585 7860 645 7920
rect 985 7970 1045 8030
rect 985 7860 1045 7920
rect 1385 7970 1445 8030
rect 1385 7860 1445 7920
rect 1785 7970 1845 8030
rect 1785 7860 1845 7920
rect 2185 7970 2245 8030
rect 2185 7860 2245 7920
rect 2585 7970 2645 8030
rect 2585 7860 2645 7920
rect 2985 7970 3045 8030
rect 2985 7860 3045 7920
rect 3385 7970 3445 8030
rect 3385 7860 3445 7920
rect 3785 7970 3845 8030
rect 3785 7860 3845 7920
rect 4185 7970 4245 8030
rect 4185 7860 4245 7920
rect 4585 7970 4645 8030
rect 4585 7860 4645 7920
rect 4985 7970 5045 8030
rect 4985 7860 5045 7920
rect 5385 7970 5445 8030
rect 5385 7860 5445 7920
rect 5785 7970 5845 8030
rect 5785 7860 5845 7920
rect 6185 7970 6245 8030
rect 6185 7860 6245 7920
rect 6585 7970 6645 8030
rect 6585 7860 6645 7920
rect 6985 7970 7045 8030
rect 6985 7860 7045 7920
rect 7385 7970 7445 8030
rect 7385 7860 7445 7920
rect 7785 7970 7845 8030
rect 7785 7860 7845 7920
rect 8185 7970 8245 8030
rect 8185 7860 8245 7920
rect 8585 7970 8645 8030
rect 8585 7860 8645 7920
rect 8985 7970 9045 8030
rect 8985 7860 9045 7920
rect 9385 7970 9445 8030
rect 9385 7860 9445 7920
rect 9785 7970 9845 8030
rect 9785 7860 9845 7920
rect 10185 7970 10245 8030
rect 10185 7860 10245 7920
rect 10585 7970 10645 8030
rect 10585 7860 10645 7920
rect 10985 7970 11045 8030
rect 10985 7860 11045 7920
rect 11385 7970 11445 8030
rect 11385 7860 11445 7920
rect 11785 7970 11845 8030
rect 11785 7860 11845 7920
rect 12185 7970 12245 8030
rect 12185 7860 12245 7920
rect 12585 7970 12645 8030
rect 12585 7860 12645 7920
rect 12985 7970 13045 8030
rect 12985 7860 13045 7920
rect -215 7600 -155 7660
rect -215 7490 -155 7550
rect 185 7600 245 7660
rect 185 7490 245 7550
rect 585 7600 645 7660
rect 585 7490 645 7550
rect 985 7600 1045 7660
rect 985 7490 1045 7550
rect 1385 7600 1445 7660
rect 1385 7490 1445 7550
rect 1785 7600 1845 7660
rect 1785 7490 1845 7550
rect 2185 7600 2245 7660
rect 2185 7490 2245 7550
rect 2585 7600 2645 7660
rect 2585 7490 2645 7550
rect 2985 7600 3045 7660
rect 2985 7490 3045 7550
rect 3385 7600 3445 7660
rect 3385 7490 3445 7550
rect 3785 7600 3845 7660
rect 3785 7490 3845 7550
rect 4185 7600 4245 7660
rect 4185 7490 4245 7550
rect 4585 7600 4645 7660
rect 4585 7490 4645 7550
rect 4985 7600 5045 7660
rect 4985 7490 5045 7550
rect 5385 7600 5445 7660
rect 5385 7490 5445 7550
rect 5785 7600 5845 7660
rect 5785 7490 5845 7550
rect 6185 7600 6245 7660
rect 6185 7490 6245 7550
rect 6585 7600 6645 7660
rect 6585 7490 6645 7550
rect 6985 7600 7045 7660
rect 6985 7490 7045 7550
rect 7385 7600 7445 7660
rect 7385 7490 7445 7550
rect 7785 7600 7845 7660
rect 7785 7490 7845 7550
rect 8185 7600 8245 7660
rect 8185 7490 8245 7550
rect 8585 7600 8645 7660
rect 8585 7490 8645 7550
rect 8985 7600 9045 7660
rect 8985 7490 9045 7550
rect 9385 7600 9445 7660
rect 9385 7490 9445 7550
rect 9785 7600 9845 7660
rect 9785 7490 9845 7550
rect 10185 7600 10245 7660
rect 10185 7490 10245 7550
rect 10585 7600 10645 7660
rect 10585 7490 10645 7550
rect 10985 7600 11045 7660
rect 10985 7490 11045 7550
rect 11385 7600 11445 7660
rect 11385 7490 11445 7550
rect 11785 7600 11845 7660
rect 11785 7490 11845 7550
rect 12185 7600 12245 7660
rect 12185 7490 12245 7550
rect 12585 7600 12645 7660
rect 12585 7490 12645 7550
rect 12985 7600 13045 7660
rect 12985 7490 13045 7550
rect -215 7230 -155 7290
rect -215 7120 -155 7180
rect 185 7230 245 7290
rect 185 7120 245 7180
rect 585 7230 645 7290
rect 585 7120 645 7180
rect 985 7230 1045 7290
rect 985 7120 1045 7180
rect 1385 7230 1445 7290
rect 1385 7120 1445 7180
rect 1785 7230 1845 7290
rect 1785 7120 1845 7180
rect 2185 7230 2245 7290
rect 2185 7120 2245 7180
rect 2585 7230 2645 7290
rect 2585 7120 2645 7180
rect 2985 7230 3045 7290
rect 2985 7120 3045 7180
rect 3385 7230 3445 7290
rect 3385 7120 3445 7180
rect 3785 7230 3845 7290
rect 3785 7120 3845 7180
rect 4185 7230 4245 7290
rect 4185 7120 4245 7180
rect 4585 7230 4645 7290
rect 4585 7120 4645 7180
rect 4985 7230 5045 7290
rect 4985 7120 5045 7180
rect 5385 7230 5445 7290
rect 5385 7120 5445 7180
rect 5785 7230 5845 7290
rect 5785 7120 5845 7180
rect 6185 7230 6245 7290
rect 6185 7120 6245 7180
rect 6585 7230 6645 7290
rect 6585 7120 6645 7180
rect 6985 7230 7045 7290
rect 6985 7120 7045 7180
rect 7385 7230 7445 7290
rect 7385 7120 7445 7180
rect 7785 7230 7845 7290
rect 7785 7120 7845 7180
rect 8185 7230 8245 7290
rect 8185 7120 8245 7180
rect 8585 7230 8645 7290
rect 8585 7120 8645 7180
rect 8985 7230 9045 7290
rect 8985 7120 9045 7180
rect 9385 7230 9445 7290
rect 9385 7120 9445 7180
rect 9785 7230 9845 7290
rect 9785 7120 9845 7180
rect 10185 7230 10245 7290
rect 10185 7120 10245 7180
rect 10585 7230 10645 7290
rect 10585 7120 10645 7180
rect 10985 7230 11045 7290
rect 10985 7120 11045 7180
rect 11385 7230 11445 7290
rect 11385 7120 11445 7180
rect 11785 7230 11845 7290
rect 11785 7120 11845 7180
rect 12185 7230 12245 7290
rect 12185 7120 12245 7180
rect 12585 7230 12645 7290
rect 12585 7120 12645 7180
rect 12985 7230 13045 7290
rect 12985 7120 13045 7180
rect -215 6860 -155 6920
rect -215 6750 -155 6810
rect 185 6860 245 6920
rect 185 6750 245 6810
rect 585 6860 645 6920
rect 585 6750 645 6810
rect 985 6860 1045 6920
rect 985 6750 1045 6810
rect 1385 6860 1445 6920
rect 1385 6750 1445 6810
rect 1785 6860 1845 6920
rect 1785 6750 1845 6810
rect 2185 6860 2245 6920
rect 2185 6750 2245 6810
rect 2585 6860 2645 6920
rect 2585 6750 2645 6810
rect 2985 6860 3045 6920
rect 2985 6750 3045 6810
rect 3385 6860 3445 6920
rect 3385 6750 3445 6810
rect 3785 6860 3845 6920
rect 3785 6750 3845 6810
rect 4185 6860 4245 6920
rect 4185 6750 4245 6810
rect 4585 6860 4645 6920
rect 4585 6750 4645 6810
rect 4985 6860 5045 6920
rect 4985 6750 5045 6810
rect 5385 6860 5445 6920
rect 5385 6750 5445 6810
rect 5785 6860 5845 6920
rect 5785 6750 5845 6810
rect 6185 6860 6245 6920
rect 6185 6750 6245 6810
rect 6585 6860 6645 6920
rect 6585 6750 6645 6810
rect 6985 6860 7045 6920
rect 6985 6750 7045 6810
rect 7385 6860 7445 6920
rect 7385 6750 7445 6810
rect 7785 6860 7845 6920
rect 7785 6750 7845 6810
rect 8185 6860 8245 6920
rect 8185 6750 8245 6810
rect 8585 6860 8645 6920
rect 8585 6750 8645 6810
rect 8985 6860 9045 6920
rect 8985 6750 9045 6810
rect 9385 6860 9445 6920
rect 9385 6750 9445 6810
rect 9785 6860 9845 6920
rect 9785 6750 9845 6810
rect 10185 6860 10245 6920
rect 10185 6750 10245 6810
rect 10585 6860 10645 6920
rect 10585 6750 10645 6810
rect 10985 6860 11045 6920
rect 10985 6750 11045 6810
rect 11385 6860 11445 6920
rect 11385 6750 11445 6810
rect 11785 6860 11845 6920
rect 11785 6750 11845 6810
rect 12185 6860 12245 6920
rect 12185 6750 12245 6810
rect 12585 6860 12645 6920
rect 12585 6750 12645 6810
rect 12985 6860 13045 6920
rect 12985 6750 13045 6810
rect -215 6490 -155 6550
rect -215 6380 -155 6440
rect 185 6490 245 6550
rect 185 6380 245 6440
rect 585 6490 645 6550
rect 585 6380 645 6440
rect 985 6490 1045 6550
rect 985 6380 1045 6440
rect 1385 6490 1445 6550
rect 1385 6380 1445 6440
rect 1785 6490 1845 6550
rect 1785 6380 1845 6440
rect 2185 6490 2245 6550
rect 2185 6380 2245 6440
rect 2585 6490 2645 6550
rect 2585 6380 2645 6440
rect 2985 6490 3045 6550
rect 2985 6380 3045 6440
rect 3385 6490 3445 6550
rect 3385 6380 3445 6440
rect 3785 6490 3845 6550
rect 3785 6380 3845 6440
rect 4185 6490 4245 6550
rect 4185 6380 4245 6440
rect 4585 6490 4645 6550
rect 4585 6380 4645 6440
rect 4985 6490 5045 6550
rect 4985 6380 5045 6440
rect 5385 6490 5445 6550
rect 5385 6380 5445 6440
rect 5785 6490 5845 6550
rect 5785 6380 5845 6440
rect 6185 6490 6245 6550
rect 6185 6380 6245 6440
rect 6585 6490 6645 6550
rect 6585 6380 6645 6440
rect 6985 6490 7045 6550
rect 6985 6380 7045 6440
rect 7385 6490 7445 6550
rect 7385 6380 7445 6440
rect 7785 6490 7845 6550
rect 7785 6380 7845 6440
rect 8185 6490 8245 6550
rect 8185 6380 8245 6440
rect 8585 6490 8645 6550
rect 8585 6380 8645 6440
rect 8985 6490 9045 6550
rect 8985 6380 9045 6440
rect 9385 6490 9445 6550
rect 9385 6380 9445 6440
rect 9785 6490 9845 6550
rect 9785 6380 9845 6440
rect 10185 6490 10245 6550
rect 10185 6380 10245 6440
rect 10585 6490 10645 6550
rect 10585 6380 10645 6440
rect 10985 6490 11045 6550
rect 10985 6380 11045 6440
rect 11385 6490 11445 6550
rect 11385 6380 11445 6440
rect 11785 6490 11845 6550
rect 11785 6380 11845 6440
rect 12185 6490 12245 6550
rect 12185 6380 12245 6440
rect 12585 6490 12645 6550
rect 12585 6380 12645 6440
rect 12985 6490 13045 6550
rect 12985 6380 13045 6440
rect -215 6120 -155 6180
rect -215 6010 -155 6070
rect 185 6120 245 6180
rect 185 6010 245 6070
rect 585 6120 645 6180
rect 585 6010 645 6070
rect 985 6120 1045 6180
rect 985 6010 1045 6070
rect 1385 6120 1445 6180
rect 1385 6010 1445 6070
rect 1785 6120 1845 6180
rect 1785 6010 1845 6070
rect 2185 6120 2245 6180
rect 2185 6010 2245 6070
rect 2585 6120 2645 6180
rect 2585 6010 2645 6070
rect 2985 6120 3045 6180
rect 2985 6010 3045 6070
rect 3385 6120 3445 6180
rect 3385 6010 3445 6070
rect 3785 6120 3845 6180
rect 3785 6010 3845 6070
rect 4185 6120 4245 6180
rect 4185 6010 4245 6070
rect 4585 6120 4645 6180
rect 4585 6010 4645 6070
rect 4985 6120 5045 6180
rect 4985 6010 5045 6070
rect 5385 6120 5445 6180
rect 5385 6010 5445 6070
rect 5785 6120 5845 6180
rect 5785 6010 5845 6070
rect 6185 6120 6245 6180
rect 6185 6010 6245 6070
rect 6585 6120 6645 6180
rect 6585 6010 6645 6070
rect 6985 6120 7045 6180
rect 6985 6010 7045 6070
rect 7385 6120 7445 6180
rect 7385 6010 7445 6070
rect 7785 6120 7845 6180
rect 7785 6010 7845 6070
rect 8185 6120 8245 6180
rect 8185 6010 8245 6070
rect 8585 6120 8645 6180
rect 8585 6010 8645 6070
rect 8985 6120 9045 6180
rect 8985 6010 9045 6070
rect 9385 6120 9445 6180
rect 9385 6010 9445 6070
rect 9785 6120 9845 6180
rect 9785 6010 9845 6070
rect 10185 6120 10245 6180
rect 10185 6010 10245 6070
rect 10585 6120 10645 6180
rect 10585 6010 10645 6070
rect 10985 6120 11045 6180
rect 10985 6010 11045 6070
rect 11385 6120 11445 6180
rect 11385 6010 11445 6070
rect 11785 6120 11845 6180
rect 11785 6010 11845 6070
rect 12185 6120 12245 6180
rect 12185 6010 12245 6070
rect 12585 6120 12645 6180
rect 12585 6010 12645 6070
rect 12985 6120 13045 6180
rect 12985 6010 13045 6070
rect -215 5750 -155 5810
rect -215 5640 -155 5700
rect 185 5750 245 5810
rect 185 5640 245 5700
rect 585 5750 645 5810
rect 585 5640 645 5700
rect 985 5750 1045 5810
rect 985 5640 1045 5700
rect 1385 5750 1445 5810
rect 1385 5640 1445 5700
rect 1785 5750 1845 5810
rect 1785 5640 1845 5700
rect 2185 5750 2245 5810
rect 2185 5640 2245 5700
rect 2585 5750 2645 5810
rect 2585 5640 2645 5700
rect 2985 5750 3045 5810
rect 2985 5640 3045 5700
rect 3385 5750 3445 5810
rect 3385 5640 3445 5700
rect 3785 5750 3845 5810
rect 3785 5640 3845 5700
rect 4185 5750 4245 5810
rect 4185 5640 4245 5700
rect 4585 5750 4645 5810
rect 4585 5640 4645 5700
rect 4985 5750 5045 5810
rect 4985 5640 5045 5700
rect 5385 5750 5445 5810
rect 5385 5640 5445 5700
rect 5785 5750 5845 5810
rect 5785 5640 5845 5700
rect 6185 5750 6245 5810
rect 6185 5640 6245 5700
rect 6585 5750 6645 5810
rect 6585 5640 6645 5700
rect 6985 5750 7045 5810
rect 6985 5640 7045 5700
rect 7385 5750 7445 5810
rect 7385 5640 7445 5700
rect 7785 5750 7845 5810
rect 7785 5640 7845 5700
rect 8185 5750 8245 5810
rect 8185 5640 8245 5700
rect 8585 5750 8645 5810
rect 8585 5640 8645 5700
rect 8985 5750 9045 5810
rect 8985 5640 9045 5700
rect 9385 5750 9445 5810
rect 9385 5640 9445 5700
rect 9785 5750 9845 5810
rect 9785 5640 9845 5700
rect 10185 5750 10245 5810
rect 10185 5640 10245 5700
rect 10585 5750 10645 5810
rect 10585 5640 10645 5700
rect 10985 5750 11045 5810
rect 10985 5640 11045 5700
rect 11385 5750 11445 5810
rect 11385 5640 11445 5700
rect 11785 5750 11845 5810
rect 11785 5640 11845 5700
rect 12185 5750 12245 5810
rect 12185 5640 12245 5700
rect 12585 5750 12645 5810
rect 12585 5640 12645 5700
rect 12985 5750 13045 5810
rect 12985 5640 13045 5700
rect -215 5380 -155 5440
rect -215 5270 -155 5330
rect 185 5380 245 5440
rect 185 5270 245 5330
rect 585 5380 645 5440
rect 585 5270 645 5330
rect 985 5380 1045 5440
rect 985 5270 1045 5330
rect 1385 5380 1445 5440
rect 1385 5270 1445 5330
rect 1785 5380 1845 5440
rect 1785 5270 1845 5330
rect 2185 5380 2245 5440
rect 2185 5270 2245 5330
rect 2585 5380 2645 5440
rect 2585 5270 2645 5330
rect 2985 5380 3045 5440
rect 2985 5270 3045 5330
rect 3385 5380 3445 5440
rect 3385 5270 3445 5330
rect 3785 5380 3845 5440
rect 3785 5270 3845 5330
rect 4185 5380 4245 5440
rect 4185 5270 4245 5330
rect 4585 5380 4645 5440
rect 4585 5270 4645 5330
rect 4985 5380 5045 5440
rect 4985 5270 5045 5330
rect 5385 5380 5445 5440
rect 5385 5270 5445 5330
rect 5785 5380 5845 5440
rect 5785 5270 5845 5330
rect 6185 5380 6245 5440
rect 6185 5270 6245 5330
rect 6585 5380 6645 5440
rect 6585 5270 6645 5330
rect 6985 5380 7045 5440
rect 6985 5270 7045 5330
rect 7385 5380 7445 5440
rect 7385 5270 7445 5330
rect 7785 5380 7845 5440
rect 7785 5270 7845 5330
rect 8185 5380 8245 5440
rect 8185 5270 8245 5330
rect 8585 5380 8645 5440
rect 8585 5270 8645 5330
rect 8985 5380 9045 5440
rect 8985 5270 9045 5330
rect 9385 5380 9445 5440
rect 9385 5270 9445 5330
rect 9785 5380 9845 5440
rect 9785 5270 9845 5330
rect 10185 5380 10245 5440
rect 10185 5270 10245 5330
rect 10585 5380 10645 5440
rect 10585 5270 10645 5330
rect 10985 5380 11045 5440
rect 10985 5270 11045 5330
rect 11385 5380 11445 5440
rect 11385 5270 11445 5330
rect 11785 5380 11845 5440
rect 11785 5270 11845 5330
rect 12185 5380 12245 5440
rect 12185 5270 12245 5330
rect 12585 5380 12645 5440
rect 12585 5270 12645 5330
rect 12985 5380 13045 5440
rect 12985 5270 13045 5330
rect -215 5010 -155 5070
rect -215 4900 -155 4960
rect 185 5010 245 5070
rect 185 4900 245 4960
rect 585 5010 645 5070
rect 585 4900 645 4960
rect 985 5010 1045 5070
rect 985 4900 1045 4960
rect 1385 5010 1445 5070
rect 1385 4900 1445 4960
rect 1785 5010 1845 5070
rect 1785 4900 1845 4960
rect 2185 5010 2245 5070
rect 2185 4900 2245 4960
rect 2585 5010 2645 5070
rect 2585 4900 2645 4960
rect 2985 5010 3045 5070
rect 2985 4900 3045 4960
rect 3385 5010 3445 5070
rect 3385 4900 3445 4960
rect 3785 5010 3845 5070
rect 3785 4900 3845 4960
rect 4185 5010 4245 5070
rect 4185 4900 4245 4960
rect 4585 5010 4645 5070
rect 4585 4900 4645 4960
rect 4985 5010 5045 5070
rect 4985 4900 5045 4960
rect 5385 5010 5445 5070
rect 5385 4900 5445 4960
rect 5785 5010 5845 5070
rect 5785 4900 5845 4960
rect 6185 5010 6245 5070
rect 6185 4900 6245 4960
rect 6585 5010 6645 5070
rect 6585 4900 6645 4960
rect 6985 5010 7045 5070
rect 6985 4900 7045 4960
rect 7385 5010 7445 5070
rect 7385 4900 7445 4960
rect 7785 5010 7845 5070
rect 7785 4900 7845 4960
rect 8185 5010 8245 5070
rect 8185 4900 8245 4960
rect 8585 5010 8645 5070
rect 8585 4900 8645 4960
rect 8985 5010 9045 5070
rect 8985 4900 9045 4960
rect 9385 5010 9445 5070
rect 9385 4900 9445 4960
rect 9785 5010 9845 5070
rect 9785 4900 9845 4960
rect 10185 5010 10245 5070
rect 10185 4900 10245 4960
rect 10585 5010 10645 5070
rect 10585 4900 10645 4960
rect 10985 5010 11045 5070
rect 10985 4900 11045 4960
rect 11385 5010 11445 5070
rect 11385 4900 11445 4960
rect 11785 5010 11845 5070
rect 11785 4900 11845 4960
rect 12185 5010 12245 5070
rect 12185 4900 12245 4960
rect 12585 5010 12645 5070
rect 12585 4900 12645 4960
rect 12985 5010 13045 5070
rect 12985 4900 13045 4960
rect -215 4640 -155 4700
rect -215 4530 -155 4590
rect 185 4640 245 4700
rect 185 4530 245 4590
rect 585 4640 645 4700
rect 585 4530 645 4590
rect 985 4640 1045 4700
rect 985 4530 1045 4590
rect 1385 4640 1445 4700
rect 1385 4530 1445 4590
rect 1785 4640 1845 4700
rect 1785 4530 1845 4590
rect 2185 4640 2245 4700
rect 2185 4530 2245 4590
rect 2585 4640 2645 4700
rect 2585 4530 2645 4590
rect 2985 4640 3045 4700
rect 2985 4530 3045 4590
rect 3385 4640 3445 4700
rect 3385 4530 3445 4590
rect 3785 4640 3845 4700
rect 3785 4530 3845 4590
rect 4185 4640 4245 4700
rect 4185 4530 4245 4590
rect 4585 4640 4645 4700
rect 4585 4530 4645 4590
rect 4985 4640 5045 4700
rect 4985 4530 5045 4590
rect 5385 4640 5445 4700
rect 5385 4530 5445 4590
rect 5785 4640 5845 4700
rect 5785 4530 5845 4590
rect 6185 4640 6245 4700
rect 6185 4530 6245 4590
rect 6585 4640 6645 4700
rect 6585 4530 6645 4590
rect 6985 4640 7045 4700
rect 6985 4530 7045 4590
rect 7385 4640 7445 4700
rect 7385 4530 7445 4590
rect 7785 4640 7845 4700
rect 7785 4530 7845 4590
rect 8185 4640 8245 4700
rect 8185 4530 8245 4590
rect 8585 4640 8645 4700
rect 8585 4530 8645 4590
rect 8985 4640 9045 4700
rect 8985 4530 9045 4590
rect 9385 4640 9445 4700
rect 9385 4530 9445 4590
rect 9785 4640 9845 4700
rect 9785 4530 9845 4590
rect 10185 4640 10245 4700
rect 10185 4530 10245 4590
rect 10585 4640 10645 4700
rect 10585 4530 10645 4590
rect 10985 4640 11045 4700
rect 10985 4530 11045 4590
rect 11385 4640 11445 4700
rect 11385 4530 11445 4590
rect 11785 4640 11845 4700
rect 11785 4530 11845 4590
rect 12185 4640 12245 4700
rect 12185 4530 12245 4590
rect 12585 4640 12645 4700
rect 12585 4530 12645 4590
rect 12985 4640 13045 4700
rect 12985 4530 13045 4590
rect -215 4270 -155 4330
rect -215 4160 -155 4220
rect 185 4270 245 4330
rect 185 4160 245 4220
rect 585 4270 645 4330
rect 585 4160 645 4220
rect 985 4270 1045 4330
rect 985 4160 1045 4220
rect 1385 4270 1445 4330
rect 1385 4160 1445 4220
rect 1785 4270 1845 4330
rect 1785 4160 1845 4220
rect 2185 4270 2245 4330
rect 2185 4160 2245 4220
rect 2585 4270 2645 4330
rect 2585 4160 2645 4220
rect 2985 4270 3045 4330
rect 2985 4160 3045 4220
rect 3385 4270 3445 4330
rect 3385 4160 3445 4220
rect 3785 4270 3845 4330
rect 3785 4160 3845 4220
rect 4185 4270 4245 4330
rect 4185 4160 4245 4220
rect 4585 4270 4645 4330
rect 4585 4160 4645 4220
rect 4985 4270 5045 4330
rect 4985 4160 5045 4220
rect 5385 4270 5445 4330
rect 5385 4160 5445 4220
rect 5785 4270 5845 4330
rect 5785 4160 5845 4220
rect 6185 4270 6245 4330
rect 6185 4160 6245 4220
rect 6585 4270 6645 4330
rect 6585 4160 6645 4220
rect 6985 4270 7045 4330
rect 6985 4160 7045 4220
rect 7385 4270 7445 4330
rect 7385 4160 7445 4220
rect 7785 4270 7845 4330
rect 7785 4160 7845 4220
rect 8185 4270 8245 4330
rect 8185 4160 8245 4220
rect 8585 4270 8645 4330
rect 8585 4160 8645 4220
rect 8985 4270 9045 4330
rect 8985 4160 9045 4220
rect 9385 4270 9445 4330
rect 9385 4160 9445 4220
rect 9785 4270 9845 4330
rect 9785 4160 9845 4220
rect 10185 4270 10245 4330
rect 10185 4160 10245 4220
rect 10585 4270 10645 4330
rect 10585 4160 10645 4220
rect 10985 4270 11045 4330
rect 10985 4160 11045 4220
rect 11385 4270 11445 4330
rect 11385 4160 11445 4220
rect 11785 4270 11845 4330
rect 11785 4160 11845 4220
rect 12185 4270 12245 4330
rect 12185 4160 12245 4220
rect 12585 4270 12645 4330
rect 12585 4160 12645 4220
rect 12985 4270 13045 4330
rect 12985 4160 13045 4220
rect -215 3900 -155 3960
rect -215 3790 -155 3850
rect 185 3900 245 3960
rect 185 3790 245 3850
rect 585 3900 645 3960
rect 585 3790 645 3850
rect 985 3900 1045 3960
rect 985 3790 1045 3850
rect 1385 3900 1445 3960
rect 1385 3790 1445 3850
rect 1785 3900 1845 3960
rect 1785 3790 1845 3850
rect 2185 3900 2245 3960
rect 2185 3790 2245 3850
rect 2585 3900 2645 3960
rect 2585 3790 2645 3850
rect 2985 3900 3045 3960
rect 2985 3790 3045 3850
rect 3385 3900 3445 3960
rect 3385 3790 3445 3850
rect 3785 3900 3845 3960
rect 3785 3790 3845 3850
rect 4185 3900 4245 3960
rect 4185 3790 4245 3850
rect 4585 3900 4645 3960
rect 4585 3790 4645 3850
rect 4985 3900 5045 3960
rect 4985 3790 5045 3850
rect 5385 3900 5445 3960
rect 5385 3790 5445 3850
rect 5785 3900 5845 3960
rect 5785 3790 5845 3850
rect 6185 3900 6245 3960
rect 6185 3790 6245 3850
rect 6585 3900 6645 3960
rect 6585 3790 6645 3850
rect 6985 3900 7045 3960
rect 6985 3790 7045 3850
rect 7385 3900 7445 3960
rect 7385 3790 7445 3850
rect 7785 3900 7845 3960
rect 7785 3790 7845 3850
rect 8185 3900 8245 3960
rect 8185 3790 8245 3850
rect 8585 3900 8645 3960
rect 8585 3790 8645 3850
rect 8985 3900 9045 3960
rect 8985 3790 9045 3850
rect 9385 3900 9445 3960
rect 9385 3790 9445 3850
rect 9785 3900 9845 3960
rect 9785 3790 9845 3850
rect 10185 3900 10245 3960
rect 10185 3790 10245 3850
rect 10585 3900 10645 3960
rect 10585 3790 10645 3850
rect 10985 3900 11045 3960
rect 10985 3790 11045 3850
rect 11385 3900 11445 3960
rect 11385 3790 11445 3850
rect 11785 3900 11845 3960
rect 11785 3790 11845 3850
rect 12185 3900 12245 3960
rect 12185 3790 12245 3850
rect 12585 3900 12645 3960
rect 12585 3790 12645 3850
rect 12985 3900 13045 3960
rect 12985 3790 13045 3850
rect -215 3530 -155 3590
rect -215 3420 -155 3480
rect 185 3530 245 3590
rect 185 3420 245 3480
rect 585 3530 645 3590
rect 585 3420 645 3480
rect 985 3530 1045 3590
rect 985 3420 1045 3480
rect 1385 3530 1445 3590
rect 1385 3420 1445 3480
rect 1785 3530 1845 3590
rect 1785 3420 1845 3480
rect 2185 3530 2245 3590
rect 2185 3420 2245 3480
rect 2585 3530 2645 3590
rect 2585 3420 2645 3480
rect 2985 3530 3045 3590
rect 2985 3420 3045 3480
rect 3385 3530 3445 3590
rect 3385 3420 3445 3480
rect 3785 3530 3845 3590
rect 3785 3420 3845 3480
rect 4185 3530 4245 3590
rect 4185 3420 4245 3480
rect 4585 3530 4645 3590
rect 4585 3420 4645 3480
rect 4985 3530 5045 3590
rect 4985 3420 5045 3480
rect 5385 3530 5445 3590
rect 5385 3420 5445 3480
rect 5785 3530 5845 3590
rect 5785 3420 5845 3480
rect 6185 3530 6245 3590
rect 6185 3420 6245 3480
rect 6585 3530 6645 3590
rect 6585 3420 6645 3480
rect 6985 3530 7045 3590
rect 6985 3420 7045 3480
rect 7385 3530 7445 3590
rect 7385 3420 7445 3480
rect 7785 3530 7845 3590
rect 7785 3420 7845 3480
rect 8185 3530 8245 3590
rect 8185 3420 8245 3480
rect 8585 3530 8645 3590
rect 8585 3420 8645 3480
rect 8985 3530 9045 3590
rect 8985 3420 9045 3480
rect 9385 3530 9445 3590
rect 9385 3420 9445 3480
rect 9785 3530 9845 3590
rect 9785 3420 9845 3480
rect 10185 3530 10245 3590
rect 10185 3420 10245 3480
rect 10585 3530 10645 3590
rect 10585 3420 10645 3480
rect 10985 3530 11045 3590
rect 10985 3420 11045 3480
rect 11385 3530 11445 3590
rect 11385 3420 11445 3480
rect 11785 3530 11845 3590
rect 11785 3420 11845 3480
rect 12185 3530 12245 3590
rect 12185 3420 12245 3480
rect 12585 3530 12645 3590
rect 12585 3420 12645 3480
rect 12985 3530 13045 3590
rect 12985 3420 13045 3480
rect -215 3160 -155 3220
rect -215 3050 -155 3110
rect 185 3160 245 3220
rect 185 3050 245 3110
rect 585 3160 645 3220
rect 585 3050 645 3110
rect 985 3160 1045 3220
rect 985 3050 1045 3110
rect 1385 3160 1445 3220
rect 1385 3050 1445 3110
rect 1785 3160 1845 3220
rect 1785 3050 1845 3110
rect 2185 3160 2245 3220
rect 2185 3050 2245 3110
rect 2585 3160 2645 3220
rect 2585 3050 2645 3110
rect 2985 3160 3045 3220
rect 2985 3050 3045 3110
rect 3385 3160 3445 3220
rect 3385 3050 3445 3110
rect 3785 3160 3845 3220
rect 3785 3050 3845 3110
rect 4185 3160 4245 3220
rect 4185 3050 4245 3110
rect 4585 3160 4645 3220
rect 4585 3050 4645 3110
rect 4985 3160 5045 3220
rect 4985 3050 5045 3110
rect 5385 3160 5445 3220
rect 5385 3050 5445 3110
rect 5785 3160 5845 3220
rect 5785 3050 5845 3110
rect 6185 3160 6245 3220
rect 6185 3050 6245 3110
rect 6585 3160 6645 3220
rect 6585 3050 6645 3110
rect 6985 3160 7045 3220
rect 6985 3050 7045 3110
rect 7385 3160 7445 3220
rect 7385 3050 7445 3110
rect 7785 3160 7845 3220
rect 7785 3050 7845 3110
rect 8185 3160 8245 3220
rect 8185 3050 8245 3110
rect 8585 3160 8645 3220
rect 8585 3050 8645 3110
rect 8985 3160 9045 3220
rect 8985 3050 9045 3110
rect 9385 3160 9445 3220
rect 9385 3050 9445 3110
rect 9785 3160 9845 3220
rect 9785 3050 9845 3110
rect 10185 3160 10245 3220
rect 10185 3050 10245 3110
rect 10585 3160 10645 3220
rect 10585 3050 10645 3110
rect 10985 3160 11045 3220
rect 10985 3050 11045 3110
rect 11385 3160 11445 3220
rect 11385 3050 11445 3110
rect 11785 3160 11845 3220
rect 11785 3050 11845 3110
rect 12185 3160 12245 3220
rect 12185 3050 12245 3110
rect 12585 3160 12645 3220
rect 12585 3050 12645 3110
rect 12985 3160 13045 3220
rect 12985 3050 13045 3110
rect -215 2790 -155 2850
rect -215 2680 -155 2740
rect 185 2790 245 2850
rect 185 2680 245 2740
rect 585 2790 645 2850
rect 585 2680 645 2740
rect 985 2790 1045 2850
rect 985 2680 1045 2740
rect 1385 2790 1445 2850
rect 1385 2680 1445 2740
rect 1785 2790 1845 2850
rect 1785 2680 1845 2740
rect 2185 2790 2245 2850
rect 2185 2680 2245 2740
rect 2585 2790 2645 2850
rect 2585 2680 2645 2740
rect 2985 2790 3045 2850
rect 2985 2680 3045 2740
rect 3385 2790 3445 2850
rect 3385 2680 3445 2740
rect 3785 2790 3845 2850
rect 3785 2680 3845 2740
rect 4185 2790 4245 2850
rect 4185 2680 4245 2740
rect 4585 2790 4645 2850
rect 4585 2680 4645 2740
rect 4985 2790 5045 2850
rect 4985 2680 5045 2740
rect 5385 2790 5445 2850
rect 5385 2680 5445 2740
rect 5785 2790 5845 2850
rect 5785 2680 5845 2740
rect 6185 2790 6245 2850
rect 6185 2680 6245 2740
rect 6585 2790 6645 2850
rect 6585 2680 6645 2740
rect 6985 2790 7045 2850
rect 6985 2680 7045 2740
rect 7385 2790 7445 2850
rect 7385 2680 7445 2740
rect 7785 2790 7845 2850
rect 7785 2680 7845 2740
rect 8185 2790 8245 2850
rect 8185 2680 8245 2740
rect 8585 2790 8645 2850
rect 8585 2680 8645 2740
rect 8985 2790 9045 2850
rect 8985 2680 9045 2740
rect 9385 2790 9445 2850
rect 9385 2680 9445 2740
rect 9785 2790 9845 2850
rect 9785 2680 9845 2740
rect 10185 2790 10245 2850
rect 10185 2680 10245 2740
rect 10585 2790 10645 2850
rect 10585 2680 10645 2740
rect 10985 2790 11045 2850
rect 10985 2680 11045 2740
rect 11385 2790 11445 2850
rect 11385 2680 11445 2740
rect 11785 2790 11845 2850
rect 11785 2680 11845 2740
rect 12185 2790 12245 2850
rect 12185 2680 12245 2740
rect 12585 2790 12645 2850
rect 12585 2680 12645 2740
rect 12985 2790 13045 2850
rect 12985 2680 13045 2740
rect -215 2420 -155 2480
rect -215 2310 -155 2370
rect 185 2420 245 2480
rect 185 2310 245 2370
rect 585 2420 645 2480
rect 585 2310 645 2370
rect 985 2420 1045 2480
rect 985 2310 1045 2370
rect 1385 2420 1445 2480
rect 1385 2310 1445 2370
rect 1785 2420 1845 2480
rect 1785 2310 1845 2370
rect 2185 2420 2245 2480
rect 2185 2310 2245 2370
rect 2585 2420 2645 2480
rect 2585 2310 2645 2370
rect 2985 2420 3045 2480
rect 2985 2310 3045 2370
rect 3385 2420 3445 2480
rect 3385 2310 3445 2370
rect 3785 2420 3845 2480
rect 3785 2310 3845 2370
rect 4185 2420 4245 2480
rect 4185 2310 4245 2370
rect 4585 2420 4645 2480
rect 4585 2310 4645 2370
rect 4985 2420 5045 2480
rect 4985 2310 5045 2370
rect 5385 2420 5445 2480
rect 5385 2310 5445 2370
rect 5785 2420 5845 2480
rect 5785 2310 5845 2370
rect 6185 2420 6245 2480
rect 6185 2310 6245 2370
rect 6585 2420 6645 2480
rect 6585 2310 6645 2370
rect 6985 2420 7045 2480
rect 6985 2310 7045 2370
rect 7385 2420 7445 2480
rect 7385 2310 7445 2370
rect 7785 2420 7845 2480
rect 7785 2310 7845 2370
rect 8185 2420 8245 2480
rect 8185 2310 8245 2370
rect 8585 2420 8645 2480
rect 8585 2310 8645 2370
rect 8985 2420 9045 2480
rect 8985 2310 9045 2370
rect 9385 2420 9445 2480
rect 9385 2310 9445 2370
rect 9785 2420 9845 2480
rect 9785 2310 9845 2370
rect 10185 2420 10245 2480
rect 10185 2310 10245 2370
rect 10585 2420 10645 2480
rect 10585 2310 10645 2370
rect 10985 2420 11045 2480
rect 10985 2310 11045 2370
rect 11385 2420 11445 2480
rect 11385 2310 11445 2370
rect 11785 2420 11845 2480
rect 11785 2310 11845 2370
rect 12185 2420 12245 2480
rect 12185 2310 12245 2370
rect 12585 2420 12645 2480
rect 12585 2310 12645 2370
rect 12985 2420 13045 2480
rect 12985 2310 13045 2370
rect -215 2050 -155 2110
rect -215 1940 -155 2000
rect 185 2050 245 2110
rect 185 1940 245 2000
rect 585 2050 645 2110
rect 585 1940 645 2000
rect 985 2050 1045 2110
rect 985 1940 1045 2000
rect 1385 2050 1445 2110
rect 1385 1940 1445 2000
rect 1785 2050 1845 2110
rect 1785 1940 1845 2000
rect 2185 2050 2245 2110
rect 2185 1940 2245 2000
rect 2585 2050 2645 2110
rect 2585 1940 2645 2000
rect 2985 2050 3045 2110
rect 2985 1940 3045 2000
rect 3385 2050 3445 2110
rect 3385 1940 3445 2000
rect 3785 2050 3845 2110
rect 3785 1940 3845 2000
rect 4185 2050 4245 2110
rect 4185 1940 4245 2000
rect 4585 2050 4645 2110
rect 4585 1940 4645 2000
rect 4985 2050 5045 2110
rect 4985 1940 5045 2000
rect 5385 2050 5445 2110
rect 5385 1940 5445 2000
rect 5785 2050 5845 2110
rect 5785 1940 5845 2000
rect 6185 2050 6245 2110
rect 6185 1940 6245 2000
rect 6585 2050 6645 2110
rect 6585 1940 6645 2000
rect 6985 2050 7045 2110
rect 6985 1940 7045 2000
rect 7385 2050 7445 2110
rect 7385 1940 7445 2000
rect 7785 2050 7845 2110
rect 7785 1940 7845 2000
rect 8185 2050 8245 2110
rect 8185 1940 8245 2000
rect 8585 2050 8645 2110
rect 8585 1940 8645 2000
rect 8985 2050 9045 2110
rect 8985 1940 9045 2000
rect 9385 2050 9445 2110
rect 9385 1940 9445 2000
rect 9785 2050 9845 2110
rect 9785 1940 9845 2000
rect 10185 2050 10245 2110
rect 10185 1940 10245 2000
rect 10585 2050 10645 2110
rect 10585 1940 10645 2000
rect 10985 2050 11045 2110
rect 10985 1940 11045 2000
rect 11385 2050 11445 2110
rect 11385 1940 11445 2000
rect 11785 2050 11845 2110
rect 11785 1940 11845 2000
rect 12185 2050 12245 2110
rect 12185 1940 12245 2000
rect 12585 2050 12645 2110
rect 12585 1940 12645 2000
rect 12985 2050 13045 2110
rect 12985 1940 13045 2000
rect -215 1680 -155 1740
rect -215 1570 -155 1630
rect 185 1680 245 1740
rect 185 1570 245 1630
rect 585 1680 645 1740
rect 585 1570 645 1630
rect 985 1680 1045 1740
rect 985 1570 1045 1630
rect 1385 1680 1445 1740
rect 1385 1570 1445 1630
rect 1785 1680 1845 1740
rect 1785 1570 1845 1630
rect 2185 1680 2245 1740
rect 2185 1570 2245 1630
rect 2585 1680 2645 1740
rect 2585 1570 2645 1630
rect 2985 1680 3045 1740
rect 2985 1570 3045 1630
rect 3385 1680 3445 1740
rect 3385 1570 3445 1630
rect 3785 1680 3845 1740
rect 3785 1570 3845 1630
rect 4185 1680 4245 1740
rect 4185 1570 4245 1630
rect 4585 1680 4645 1740
rect 4585 1570 4645 1630
rect 4985 1680 5045 1740
rect 4985 1570 5045 1630
rect 5385 1680 5445 1740
rect 5385 1570 5445 1630
rect 5785 1680 5845 1740
rect 5785 1570 5845 1630
rect 6185 1680 6245 1740
rect 6185 1570 6245 1630
rect 6585 1680 6645 1740
rect 6585 1570 6645 1630
rect 6985 1680 7045 1740
rect 6985 1570 7045 1630
rect 7385 1680 7445 1740
rect 7385 1570 7445 1630
rect 7785 1680 7845 1740
rect 7785 1570 7845 1630
rect 8185 1680 8245 1740
rect 8185 1570 8245 1630
rect 8585 1680 8645 1740
rect 8585 1570 8645 1630
rect 8985 1680 9045 1740
rect 8985 1570 9045 1630
rect 9385 1680 9445 1740
rect 9385 1570 9445 1630
rect 9785 1680 9845 1740
rect 9785 1570 9845 1630
rect 10185 1680 10245 1740
rect 10185 1570 10245 1630
rect 10585 1680 10645 1740
rect 10585 1570 10645 1630
rect 10985 1680 11045 1740
rect 10985 1570 11045 1630
rect 11385 1680 11445 1740
rect 11385 1570 11445 1630
rect 11785 1680 11845 1740
rect 11785 1570 11845 1630
rect 12185 1680 12245 1740
rect 12185 1570 12245 1630
rect 12585 1680 12645 1740
rect 12585 1570 12645 1630
rect 12985 1680 13045 1740
rect 12985 1570 13045 1630
rect -215 1310 -155 1370
rect -215 1200 -155 1260
rect 185 1310 245 1370
rect 185 1200 245 1260
rect 585 1310 645 1370
rect 585 1200 645 1260
rect 985 1310 1045 1370
rect 985 1200 1045 1260
rect 1385 1310 1445 1370
rect 1385 1200 1445 1260
rect 1785 1310 1845 1370
rect 1785 1200 1845 1260
rect 2185 1310 2245 1370
rect 2185 1200 2245 1260
rect 2585 1310 2645 1370
rect 2585 1200 2645 1260
rect 2985 1310 3045 1370
rect 2985 1200 3045 1260
rect 3385 1310 3445 1370
rect 3385 1200 3445 1260
rect 3785 1310 3845 1370
rect 3785 1200 3845 1260
rect 4185 1310 4245 1370
rect 4185 1200 4245 1260
rect 4585 1310 4645 1370
rect 4585 1200 4645 1260
rect 4985 1310 5045 1370
rect 4985 1200 5045 1260
rect 5385 1310 5445 1370
rect 5385 1200 5445 1260
rect 5785 1310 5845 1370
rect 5785 1200 5845 1260
rect 6185 1310 6245 1370
rect 6185 1200 6245 1260
rect 6585 1310 6645 1370
rect 6585 1200 6645 1260
rect 6985 1310 7045 1370
rect 6985 1200 7045 1260
rect 7385 1310 7445 1370
rect 7385 1200 7445 1260
rect 7785 1310 7845 1370
rect 7785 1200 7845 1260
rect 8185 1310 8245 1370
rect 8185 1200 8245 1260
rect 8585 1310 8645 1370
rect 8585 1200 8645 1260
rect 8985 1310 9045 1370
rect 8985 1200 9045 1260
rect 9385 1310 9445 1370
rect 9385 1200 9445 1260
rect 9785 1310 9845 1370
rect 9785 1200 9845 1260
rect 10185 1310 10245 1370
rect 10185 1200 10245 1260
rect 10585 1310 10645 1370
rect 10585 1200 10645 1260
rect 10985 1310 11045 1370
rect 10985 1200 11045 1260
rect 11385 1310 11445 1370
rect 11385 1200 11445 1260
rect 11785 1310 11845 1370
rect 11785 1200 11845 1260
rect 12185 1310 12245 1370
rect 12185 1200 12245 1260
rect 12585 1310 12645 1370
rect 12585 1200 12645 1260
rect 12985 1310 13045 1370
rect 12985 1200 13045 1260
rect -215 940 -155 1000
rect -215 830 -155 890
rect 185 940 245 1000
rect 185 830 245 890
rect 585 940 645 1000
rect 585 830 645 890
rect 985 940 1045 1000
rect 985 830 1045 890
rect 1385 940 1445 1000
rect 1385 830 1445 890
rect 1785 940 1845 1000
rect 1785 830 1845 890
rect 2185 940 2245 1000
rect 2185 830 2245 890
rect 2585 940 2645 1000
rect 2585 830 2645 890
rect 2985 940 3045 1000
rect 2985 830 3045 890
rect 3385 940 3445 1000
rect 3385 830 3445 890
rect 3785 940 3845 1000
rect 3785 830 3845 890
rect 4185 940 4245 1000
rect 4185 830 4245 890
rect 4585 940 4645 1000
rect 4585 830 4645 890
rect 4985 940 5045 1000
rect 4985 830 5045 890
rect 5385 940 5445 1000
rect 5385 830 5445 890
rect 5785 940 5845 1000
rect 5785 830 5845 890
rect 6185 940 6245 1000
rect 6185 830 6245 890
rect 6585 940 6645 1000
rect 6585 830 6645 890
rect 6985 940 7045 1000
rect 6985 830 7045 890
rect 7385 940 7445 1000
rect 7385 830 7445 890
rect 7785 940 7845 1000
rect 7785 830 7845 890
rect 8185 940 8245 1000
rect 8185 830 8245 890
rect 8585 940 8645 1000
rect 8585 830 8645 890
rect 8985 940 9045 1000
rect 8985 830 9045 890
rect 9385 940 9445 1000
rect 9385 830 9445 890
rect 9785 940 9845 1000
rect 9785 830 9845 890
rect 10185 940 10245 1000
rect 10185 830 10245 890
rect 10585 940 10645 1000
rect 10585 830 10645 890
rect 10985 940 11045 1000
rect 10985 830 11045 890
rect 11385 940 11445 1000
rect 11385 830 11445 890
rect 11785 940 11845 1000
rect 11785 830 11845 890
rect 12185 940 12245 1000
rect 12185 830 12245 890
rect 12585 940 12645 1000
rect 12585 830 12645 890
rect 12985 940 13045 1000
rect 12985 830 13045 890
rect -215 570 -155 630
rect -215 460 -155 520
rect 185 570 245 630
rect 185 460 245 520
rect 585 570 645 630
rect 585 460 645 520
rect 985 570 1045 630
rect 985 460 1045 520
rect 1385 570 1445 630
rect 1385 460 1445 520
rect 1785 570 1845 630
rect 1785 460 1845 520
rect 2185 570 2245 630
rect 2185 460 2245 520
rect 2585 570 2645 630
rect 2585 460 2645 520
rect 2985 570 3045 630
rect 2985 460 3045 520
rect 3385 570 3445 630
rect 3385 460 3445 520
rect 3785 570 3845 630
rect 3785 460 3845 520
rect 4185 570 4245 630
rect 4185 460 4245 520
rect 4585 570 4645 630
rect 4585 460 4645 520
rect 4985 570 5045 630
rect 4985 460 5045 520
rect 5385 570 5445 630
rect 5385 460 5445 520
rect 5785 570 5845 630
rect 5785 460 5845 520
rect 6185 570 6245 630
rect 6185 460 6245 520
rect 6585 570 6645 630
rect 6585 460 6645 520
rect 6985 570 7045 630
rect 6985 460 7045 520
rect 7385 570 7445 630
rect 7385 460 7445 520
rect 7785 570 7845 630
rect 7785 460 7845 520
rect 8185 570 8245 630
rect 8185 460 8245 520
rect 8585 570 8645 630
rect 8585 460 8645 520
rect 8985 570 9045 630
rect 8985 460 9045 520
rect 9385 570 9445 630
rect 9385 460 9445 520
rect 9785 570 9845 630
rect 9785 460 9845 520
rect 10185 570 10245 630
rect 10185 460 10245 520
rect 10585 570 10645 630
rect 10585 460 10645 520
rect 10985 570 11045 630
rect 10985 460 11045 520
rect 11385 570 11445 630
rect 11385 460 11445 520
rect 11785 570 11845 630
rect 11785 460 11845 520
rect 12185 570 12245 630
rect 12185 460 12245 520
rect 12585 570 12645 630
rect 12585 460 12645 520
rect 12985 570 13045 630
rect 12985 460 13045 520
rect -215 200 -155 260
rect -215 90 -155 150
rect 185 200 245 260
rect 185 90 245 150
rect 585 200 645 260
rect 585 90 645 150
rect 985 200 1045 260
rect 985 90 1045 150
rect 1385 200 1445 260
rect 1385 90 1445 150
rect 1785 200 1845 260
rect 1785 90 1845 150
rect 2185 200 2245 260
rect 2185 90 2245 150
rect 2585 200 2645 260
rect 2585 90 2645 150
rect 2985 200 3045 260
rect 2985 90 3045 150
rect 3385 200 3445 260
rect 3385 90 3445 150
rect 3785 200 3845 260
rect 3785 90 3845 150
rect 4185 200 4245 260
rect 4185 90 4245 150
rect 4585 200 4645 260
rect 4585 90 4645 150
rect 4985 200 5045 260
rect 4985 90 5045 150
rect 5385 200 5445 260
rect 5385 90 5445 150
rect 5785 200 5845 260
rect 5785 90 5845 150
rect 6185 200 6245 260
rect 6185 90 6245 150
rect 6585 200 6645 260
rect 6585 90 6645 150
rect 6985 200 7045 260
rect 6985 90 7045 150
rect 7385 200 7445 260
rect 7385 90 7445 150
rect 7785 200 7845 260
rect 7785 90 7845 150
rect 8185 200 8245 260
rect 8185 90 8245 150
rect 8585 200 8645 260
rect 8585 90 8645 150
rect 8985 200 9045 260
rect 8985 90 9045 150
rect 9385 200 9445 260
rect 9385 90 9445 150
rect 9785 200 9845 260
rect 9785 90 9845 150
rect 10185 200 10245 260
rect 10185 90 10245 150
rect 10585 200 10645 260
rect 10585 90 10645 150
rect 10985 200 11045 260
rect 10985 90 11045 150
rect 11385 200 11445 260
rect 11385 90 11445 150
rect 11785 200 11845 260
rect 11785 90 11845 150
rect 12185 200 12245 260
rect 12185 90 12245 150
rect 12585 200 12645 260
rect 12585 90 12645 150
rect 12985 200 13045 260
rect 12985 90 13045 150
rect -215 -170 -155 -110
rect -215 -280 -155 -220
rect 185 -170 245 -110
rect 185 -280 245 -220
rect 585 -170 645 -110
rect 585 -280 645 -220
rect 985 -170 1045 -110
rect 985 -280 1045 -220
rect 1385 -170 1445 -110
rect 1385 -280 1445 -220
rect 1785 -170 1845 -110
rect 1785 -280 1845 -220
rect 2185 -170 2245 -110
rect 2185 -280 2245 -220
rect 2585 -170 2645 -110
rect 2585 -280 2645 -220
rect 2985 -170 3045 -110
rect 2985 -280 3045 -220
rect 3385 -170 3445 -110
rect 3385 -280 3445 -220
rect 3785 -170 3845 -110
rect 3785 -280 3845 -220
rect 4185 -170 4245 -110
rect 4185 -280 4245 -220
rect 4585 -170 4645 -110
rect 4585 -280 4645 -220
rect 4985 -170 5045 -110
rect 4985 -280 5045 -220
rect 5385 -170 5445 -110
rect 5385 -280 5445 -220
rect 5785 -170 5845 -110
rect 5785 -280 5845 -220
rect 6185 -170 6245 -110
rect 6185 -280 6245 -220
rect 6585 -170 6645 -110
rect 6585 -280 6645 -220
rect 6985 -170 7045 -110
rect 6985 -280 7045 -220
rect 7385 -170 7445 -110
rect 7385 -280 7445 -220
rect 7785 -170 7845 -110
rect 7785 -280 7845 -220
rect 8185 -170 8245 -110
rect 8185 -280 8245 -220
rect 8585 -170 8645 -110
rect 8585 -280 8645 -220
rect 8985 -170 9045 -110
rect 8985 -280 9045 -220
rect 9385 -170 9445 -110
rect 9385 -280 9445 -220
rect 9785 -170 9845 -110
rect 9785 -280 9845 -220
rect 10185 -170 10245 -110
rect 10185 -280 10245 -220
rect 10585 -170 10645 -110
rect 10585 -280 10645 -220
rect 10985 -170 11045 -110
rect 10985 -280 11045 -220
rect 11385 -170 11445 -110
rect 11385 -280 11445 -220
rect 11785 -170 11845 -110
rect 11785 -280 11845 -220
rect 12185 -170 12245 -110
rect 12185 -280 12245 -220
rect 12585 -170 12645 -110
rect 12585 -280 12645 -220
rect 12985 -170 13045 -110
rect 12985 -280 13045 -220
<< metal3 >>
rect -275 24180 -95 24185
rect -275 24120 -265 24180
rect -205 24120 -165 24180
rect -105 24120 -95 24180
rect -275 24115 -95 24120
rect -215 23945 -155 24115
rect 12895 24055 12905 24135
rect 12985 24055 13035 24135
rect 13115 24055 13125 24135
rect 185 23945 245 24040
rect 585 23945 645 24040
rect 985 23945 1045 24040
rect 1385 23945 1445 24040
rect 1785 23945 1845 24040
rect 2185 23945 2245 24040
rect 2585 23945 2645 24040
rect 2985 23945 3045 24040
rect 3385 23945 3445 24040
rect 3785 23945 3845 24040
rect 4185 23945 4245 24040
rect 4585 23945 4645 24040
rect 4985 23945 5045 24040
rect 5385 23945 5445 24040
rect 5785 23945 5845 24040
rect 6185 23945 6245 24040
rect 6585 23945 6645 24040
rect 6985 23945 7045 24040
rect 7385 23945 7445 24040
rect 7785 23945 7845 24040
rect 8185 23945 8245 24040
rect 8585 23945 8645 24040
rect 8985 23945 9045 24040
rect 9385 23945 9445 24040
rect 9785 23945 9845 24040
rect 10185 23945 10245 24040
rect 10585 23945 10645 24040
rect 10985 23945 11045 24040
rect 11385 23945 11445 24040
rect 11785 23945 11845 24040
rect 12185 23945 12245 24040
rect 12585 23945 12645 24040
rect 12985 23945 13045 24055
rect -225 23940 -145 23945
rect -225 23880 -215 23940
rect -155 23880 -145 23940
rect -225 23830 -145 23880
rect 170 23875 180 23945
rect 250 23875 260 23945
rect 570 23875 580 23945
rect 650 23875 660 23945
rect 970 23875 980 23945
rect 1050 23875 1060 23945
rect 1370 23875 1380 23945
rect 1450 23875 1460 23945
rect 1770 23875 1780 23945
rect 1850 23875 1860 23945
rect 2170 23875 2180 23945
rect 2250 23875 2260 23945
rect 2570 23875 2580 23945
rect 2650 23875 2660 23945
rect 2970 23875 2980 23945
rect 3050 23875 3060 23945
rect 3370 23875 3380 23945
rect 3450 23875 3460 23945
rect 3770 23875 3780 23945
rect 3850 23875 3860 23945
rect 4170 23875 4180 23945
rect 4250 23875 4260 23945
rect 4570 23875 4580 23945
rect 4650 23875 4660 23945
rect 4970 23875 4980 23945
rect 5050 23875 5060 23945
rect 5370 23875 5380 23945
rect 5450 23875 5460 23945
rect 5770 23875 5780 23945
rect 5850 23875 5860 23945
rect 6170 23875 6180 23945
rect 6250 23875 6260 23945
rect 6570 23875 6580 23945
rect 6650 23875 6660 23945
rect 6970 23875 6980 23945
rect 7050 23875 7060 23945
rect 7370 23875 7380 23945
rect 7450 23875 7460 23945
rect 7770 23875 7780 23945
rect 7850 23875 7860 23945
rect 8170 23875 8180 23945
rect 8250 23875 8260 23945
rect 8570 23875 8580 23945
rect 8650 23875 8660 23945
rect 8970 23875 8980 23945
rect 9050 23875 9060 23945
rect 9370 23875 9380 23945
rect 9450 23875 9460 23945
rect 9770 23875 9780 23945
rect 9850 23875 9860 23945
rect 10170 23875 10180 23945
rect 10250 23875 10260 23945
rect 10570 23875 10580 23945
rect 10650 23875 10660 23945
rect 10970 23875 10980 23945
rect 11050 23875 11060 23945
rect 11370 23875 11380 23945
rect 11450 23875 11460 23945
rect 11770 23875 11780 23945
rect 11850 23875 11860 23945
rect 12170 23875 12180 23945
rect 12250 23875 12260 23945
rect 12570 23875 12580 23945
rect 12650 23875 12660 23945
rect 12975 23940 13055 23945
rect 12975 23880 12985 23940
rect 13045 23880 13055 23940
rect -225 23770 -215 23830
rect -155 23770 -145 23830
rect -225 23765 -145 23770
rect 175 23830 255 23875
rect 175 23770 185 23830
rect 245 23770 255 23830
rect 175 23765 255 23770
rect 575 23830 655 23875
rect 575 23770 585 23830
rect 645 23770 655 23830
rect 575 23765 655 23770
rect 975 23830 1055 23875
rect 975 23770 985 23830
rect 1045 23770 1055 23830
rect 975 23765 1055 23770
rect 1375 23830 1455 23875
rect 1375 23770 1385 23830
rect 1445 23770 1455 23830
rect 1375 23765 1455 23770
rect 1775 23830 1855 23875
rect 1775 23770 1785 23830
rect 1845 23770 1855 23830
rect 1775 23765 1855 23770
rect 2175 23830 2255 23875
rect 2175 23770 2185 23830
rect 2245 23770 2255 23830
rect 2175 23765 2255 23770
rect 2575 23830 2655 23875
rect 2575 23770 2585 23830
rect 2645 23770 2655 23830
rect 2575 23765 2655 23770
rect 2975 23830 3055 23875
rect 2975 23770 2985 23830
rect 3045 23770 3055 23830
rect 2975 23765 3055 23770
rect 3375 23830 3455 23875
rect 3375 23770 3385 23830
rect 3445 23770 3455 23830
rect 3375 23765 3455 23770
rect 3775 23830 3855 23875
rect 3775 23770 3785 23830
rect 3845 23770 3855 23830
rect 3775 23765 3855 23770
rect 4175 23830 4255 23875
rect 4175 23770 4185 23830
rect 4245 23770 4255 23830
rect 4175 23765 4255 23770
rect 4575 23830 4655 23875
rect 4575 23770 4585 23830
rect 4645 23770 4655 23830
rect 4575 23765 4655 23770
rect 4975 23830 5055 23875
rect 4975 23770 4985 23830
rect 5045 23770 5055 23830
rect 4975 23765 5055 23770
rect 5375 23830 5455 23875
rect 5375 23770 5385 23830
rect 5445 23770 5455 23830
rect 5375 23765 5455 23770
rect 5775 23830 5855 23875
rect 5775 23770 5785 23830
rect 5845 23770 5855 23830
rect 5775 23765 5855 23770
rect 6175 23830 6255 23875
rect 6175 23770 6185 23830
rect 6245 23770 6255 23830
rect 6175 23765 6255 23770
rect 6575 23830 6655 23875
rect 6575 23770 6585 23830
rect 6645 23770 6655 23830
rect 6575 23765 6655 23770
rect 6975 23830 7055 23875
rect 6975 23770 6985 23830
rect 7045 23770 7055 23830
rect 6975 23765 7055 23770
rect 7375 23830 7455 23875
rect 7375 23770 7385 23830
rect 7445 23770 7455 23830
rect 7375 23765 7455 23770
rect 7775 23830 7855 23875
rect 7775 23770 7785 23830
rect 7845 23770 7855 23830
rect 7775 23765 7855 23770
rect 8175 23830 8255 23875
rect 8175 23770 8185 23830
rect 8245 23770 8255 23830
rect 8175 23765 8255 23770
rect 8575 23830 8655 23875
rect 8575 23770 8585 23830
rect 8645 23770 8655 23830
rect 8575 23765 8655 23770
rect 8975 23830 9055 23875
rect 8975 23770 8985 23830
rect 9045 23770 9055 23830
rect 8975 23765 9055 23770
rect 9375 23830 9455 23875
rect 9375 23770 9385 23830
rect 9445 23770 9455 23830
rect 9375 23765 9455 23770
rect 9775 23830 9855 23875
rect 9775 23770 9785 23830
rect 9845 23770 9855 23830
rect 9775 23765 9855 23770
rect 10175 23830 10255 23875
rect 10175 23770 10185 23830
rect 10245 23770 10255 23830
rect 10175 23765 10255 23770
rect 10575 23830 10655 23875
rect 10575 23770 10585 23830
rect 10645 23770 10655 23830
rect 10575 23765 10655 23770
rect 10975 23830 11055 23875
rect 10975 23770 10985 23830
rect 11045 23770 11055 23830
rect 10975 23765 11055 23770
rect 11375 23830 11455 23875
rect 11375 23770 11385 23830
rect 11445 23770 11455 23830
rect 11375 23765 11455 23770
rect 11775 23830 11855 23875
rect 11775 23770 11785 23830
rect 11845 23770 11855 23830
rect 11775 23765 11855 23770
rect 12175 23830 12255 23875
rect 12175 23770 12185 23830
rect 12245 23770 12255 23830
rect 12175 23765 12255 23770
rect 12575 23830 12655 23875
rect 12575 23770 12585 23830
rect 12645 23770 12655 23830
rect 12575 23765 12655 23770
rect 12975 23830 13055 23880
rect 12975 23770 12985 23830
rect 13045 23770 13055 23830
rect 12975 23765 13055 23770
rect -215 23575 -155 23765
rect 185 23575 245 23765
rect 585 23575 645 23765
rect 985 23575 1045 23765
rect 1385 23575 1445 23765
rect 1785 23575 1845 23765
rect 2185 23575 2245 23765
rect 2585 23575 2645 23765
rect 2985 23575 3045 23765
rect 3385 23575 3445 23765
rect 3785 23575 3845 23765
rect 4185 23575 4245 23765
rect 4585 23575 4645 23765
rect 4985 23575 5045 23765
rect 5385 23575 5445 23765
rect 5785 23575 5845 23765
rect 6185 23575 6245 23765
rect 6585 23575 6645 23765
rect 6985 23575 7045 23765
rect 7385 23575 7445 23765
rect 7785 23575 7845 23765
rect 8185 23575 8245 23765
rect 8585 23575 8645 23765
rect 8985 23575 9045 23765
rect 9385 23575 9445 23765
rect 9785 23575 9845 23765
rect 10185 23575 10245 23765
rect 10585 23575 10645 23765
rect 10985 23575 11045 23765
rect 11385 23575 11445 23765
rect 11785 23575 11845 23765
rect 12185 23575 12245 23765
rect 12585 23575 12645 23765
rect 12985 23575 13045 23765
rect -225 23570 -145 23575
rect -225 23510 -215 23570
rect -155 23510 -145 23570
rect -225 23460 -145 23510
rect -225 23400 -215 23460
rect -155 23400 -145 23460
rect -225 23395 -145 23400
rect 175 23570 255 23575
rect 175 23510 185 23570
rect 245 23510 255 23570
rect 175 23460 255 23510
rect 175 23400 185 23460
rect 245 23400 255 23460
rect 175 23395 255 23400
rect 575 23570 655 23575
rect 575 23510 585 23570
rect 645 23510 655 23570
rect 575 23460 655 23510
rect 575 23400 585 23460
rect 645 23400 655 23460
rect 575 23395 655 23400
rect 975 23570 1055 23575
rect 975 23510 985 23570
rect 1045 23510 1055 23570
rect 975 23460 1055 23510
rect 975 23400 985 23460
rect 1045 23400 1055 23460
rect 975 23395 1055 23400
rect 1375 23570 1455 23575
rect 1375 23510 1385 23570
rect 1445 23510 1455 23570
rect 1375 23460 1455 23510
rect 1375 23400 1385 23460
rect 1445 23400 1455 23460
rect 1375 23395 1455 23400
rect 1775 23570 1855 23575
rect 1775 23510 1785 23570
rect 1845 23510 1855 23570
rect 1775 23460 1855 23510
rect 1775 23400 1785 23460
rect 1845 23400 1855 23460
rect 1775 23395 1855 23400
rect 2175 23570 2255 23575
rect 2175 23510 2185 23570
rect 2245 23510 2255 23570
rect 2175 23460 2255 23510
rect 2175 23400 2185 23460
rect 2245 23400 2255 23460
rect 2175 23395 2255 23400
rect 2575 23570 2655 23575
rect 2575 23510 2585 23570
rect 2645 23510 2655 23570
rect 2575 23460 2655 23510
rect 2575 23400 2585 23460
rect 2645 23400 2655 23460
rect 2575 23395 2655 23400
rect 2975 23570 3055 23575
rect 2975 23510 2985 23570
rect 3045 23510 3055 23570
rect 2975 23460 3055 23510
rect 2975 23400 2985 23460
rect 3045 23400 3055 23460
rect 2975 23395 3055 23400
rect 3375 23570 3455 23575
rect 3375 23510 3385 23570
rect 3445 23510 3455 23570
rect 3375 23460 3455 23510
rect 3375 23400 3385 23460
rect 3445 23400 3455 23460
rect 3375 23395 3455 23400
rect 3775 23570 3855 23575
rect 3775 23510 3785 23570
rect 3845 23510 3855 23570
rect 3775 23460 3855 23510
rect 3775 23400 3785 23460
rect 3845 23400 3855 23460
rect 3775 23395 3855 23400
rect 4175 23570 4255 23575
rect 4175 23510 4185 23570
rect 4245 23510 4255 23570
rect 4175 23460 4255 23510
rect 4175 23400 4185 23460
rect 4245 23400 4255 23460
rect 4175 23395 4255 23400
rect 4575 23570 4655 23575
rect 4575 23510 4585 23570
rect 4645 23510 4655 23570
rect 4575 23460 4655 23510
rect 4575 23400 4585 23460
rect 4645 23400 4655 23460
rect 4575 23395 4655 23400
rect 4975 23570 5055 23575
rect 4975 23510 4985 23570
rect 5045 23510 5055 23570
rect 4975 23460 5055 23510
rect 4975 23400 4985 23460
rect 5045 23400 5055 23460
rect 4975 23395 5055 23400
rect 5375 23570 5455 23575
rect 5375 23510 5385 23570
rect 5445 23510 5455 23570
rect 5375 23460 5455 23510
rect 5375 23400 5385 23460
rect 5445 23400 5455 23460
rect 5375 23395 5455 23400
rect 5775 23570 5855 23575
rect 5775 23510 5785 23570
rect 5845 23510 5855 23570
rect 5775 23460 5855 23510
rect 5775 23400 5785 23460
rect 5845 23400 5855 23460
rect 5775 23395 5855 23400
rect 6175 23570 6255 23575
rect 6175 23510 6185 23570
rect 6245 23510 6255 23570
rect 6175 23460 6255 23510
rect 6175 23400 6185 23460
rect 6245 23400 6255 23460
rect 6175 23395 6255 23400
rect 6575 23570 6655 23575
rect 6575 23510 6585 23570
rect 6645 23510 6655 23570
rect 6575 23460 6655 23510
rect 6575 23400 6585 23460
rect 6645 23400 6655 23460
rect 6575 23395 6655 23400
rect 6975 23570 7055 23575
rect 6975 23510 6985 23570
rect 7045 23510 7055 23570
rect 6975 23460 7055 23510
rect 6975 23400 6985 23460
rect 7045 23400 7055 23460
rect 6975 23395 7055 23400
rect 7375 23570 7455 23575
rect 7375 23510 7385 23570
rect 7445 23510 7455 23570
rect 7375 23460 7455 23510
rect 7375 23400 7385 23460
rect 7445 23400 7455 23460
rect 7375 23395 7455 23400
rect 7775 23570 7855 23575
rect 7775 23510 7785 23570
rect 7845 23510 7855 23570
rect 7775 23460 7855 23510
rect 7775 23400 7785 23460
rect 7845 23400 7855 23460
rect 7775 23395 7855 23400
rect 8175 23570 8255 23575
rect 8175 23510 8185 23570
rect 8245 23510 8255 23570
rect 8175 23460 8255 23510
rect 8175 23400 8185 23460
rect 8245 23400 8255 23460
rect 8175 23395 8255 23400
rect 8575 23570 8655 23575
rect 8575 23510 8585 23570
rect 8645 23510 8655 23570
rect 8575 23460 8655 23510
rect 8575 23400 8585 23460
rect 8645 23400 8655 23460
rect 8575 23395 8655 23400
rect 8975 23570 9055 23575
rect 8975 23510 8985 23570
rect 9045 23510 9055 23570
rect 8975 23460 9055 23510
rect 8975 23400 8985 23460
rect 9045 23400 9055 23460
rect 8975 23395 9055 23400
rect 9375 23570 9455 23575
rect 9375 23510 9385 23570
rect 9445 23510 9455 23570
rect 9375 23460 9455 23510
rect 9375 23400 9385 23460
rect 9445 23400 9455 23460
rect 9375 23395 9455 23400
rect 9775 23570 9855 23575
rect 9775 23510 9785 23570
rect 9845 23510 9855 23570
rect 9775 23460 9855 23510
rect 9775 23400 9785 23460
rect 9845 23400 9855 23460
rect 9775 23395 9855 23400
rect 10175 23570 10255 23575
rect 10175 23510 10185 23570
rect 10245 23510 10255 23570
rect 10175 23460 10255 23510
rect 10175 23400 10185 23460
rect 10245 23400 10255 23460
rect 10175 23395 10255 23400
rect 10575 23570 10655 23575
rect 10575 23510 10585 23570
rect 10645 23510 10655 23570
rect 10575 23460 10655 23510
rect 10575 23400 10585 23460
rect 10645 23400 10655 23460
rect 10575 23395 10655 23400
rect 10975 23570 11055 23575
rect 10975 23510 10985 23570
rect 11045 23510 11055 23570
rect 10975 23460 11055 23510
rect 10975 23400 10985 23460
rect 11045 23400 11055 23460
rect 10975 23395 11055 23400
rect 11375 23570 11455 23575
rect 11375 23510 11385 23570
rect 11445 23510 11455 23570
rect 11375 23460 11455 23510
rect 11375 23400 11385 23460
rect 11445 23400 11455 23460
rect 11375 23395 11455 23400
rect 11775 23570 11855 23575
rect 11775 23510 11785 23570
rect 11845 23510 11855 23570
rect 11775 23460 11855 23510
rect 11775 23400 11785 23460
rect 11845 23400 11855 23460
rect 11775 23395 11855 23400
rect 12175 23570 12255 23575
rect 12175 23510 12185 23570
rect 12245 23510 12255 23570
rect 12175 23460 12255 23510
rect 12175 23400 12185 23460
rect 12245 23400 12255 23460
rect 12175 23395 12255 23400
rect 12575 23570 12655 23575
rect 12575 23510 12585 23570
rect 12645 23510 12655 23570
rect 12575 23460 12655 23510
rect 12575 23400 12585 23460
rect 12645 23400 12655 23460
rect 12575 23395 12655 23400
rect 12975 23570 13055 23575
rect 12975 23510 12985 23570
rect 13045 23510 13055 23570
rect 12975 23460 13055 23510
rect 12975 23400 12985 23460
rect 13045 23400 13055 23460
rect 12975 23395 13055 23400
rect -215 23205 -155 23395
rect 185 23205 245 23395
rect 585 23205 645 23395
rect 985 23205 1045 23395
rect 1385 23205 1445 23395
rect 1785 23205 1845 23395
rect 2185 23205 2245 23395
rect 2585 23205 2645 23395
rect 2985 23205 3045 23395
rect 3385 23205 3445 23395
rect 3785 23205 3845 23395
rect 4185 23205 4245 23395
rect 4585 23205 4645 23395
rect 4985 23205 5045 23395
rect 5385 23205 5445 23395
rect 5785 23205 5845 23395
rect 6185 23205 6245 23395
rect 6585 23205 6645 23395
rect 6985 23205 7045 23395
rect 7385 23205 7445 23395
rect 7785 23205 7845 23395
rect 8185 23205 8245 23395
rect 8585 23205 8645 23395
rect 8985 23205 9045 23395
rect 9385 23205 9445 23395
rect 9785 23205 9845 23395
rect 10185 23205 10245 23395
rect 10585 23205 10645 23395
rect 10985 23205 11045 23395
rect 11385 23205 11445 23395
rect 11785 23205 11845 23395
rect 12185 23205 12245 23395
rect 12585 23205 12645 23395
rect 12985 23205 13045 23395
rect -225 23200 -145 23205
rect -225 23140 -215 23200
rect -155 23140 -145 23200
rect -225 23090 -145 23140
rect -225 23030 -215 23090
rect -155 23030 -145 23090
rect -225 23025 -145 23030
rect 175 23200 255 23205
rect 175 23140 185 23200
rect 245 23140 255 23200
rect 175 23090 255 23140
rect 175 23030 185 23090
rect 245 23030 255 23090
rect 175 23025 255 23030
rect 575 23200 655 23205
rect 575 23140 585 23200
rect 645 23140 655 23200
rect 575 23090 655 23140
rect 575 23030 585 23090
rect 645 23030 655 23090
rect 575 23025 655 23030
rect 975 23200 1055 23205
rect 975 23140 985 23200
rect 1045 23140 1055 23200
rect 975 23090 1055 23140
rect 975 23030 985 23090
rect 1045 23030 1055 23090
rect 975 23025 1055 23030
rect 1375 23200 1455 23205
rect 1375 23140 1385 23200
rect 1445 23140 1455 23200
rect 1375 23090 1455 23140
rect 1375 23030 1385 23090
rect 1445 23030 1455 23090
rect 1375 23025 1455 23030
rect 1775 23200 1855 23205
rect 1775 23140 1785 23200
rect 1845 23140 1855 23200
rect 1775 23090 1855 23140
rect 1775 23030 1785 23090
rect 1845 23030 1855 23090
rect 1775 23025 1855 23030
rect 2175 23200 2255 23205
rect 2175 23140 2185 23200
rect 2245 23140 2255 23200
rect 2175 23090 2255 23140
rect 2175 23030 2185 23090
rect 2245 23030 2255 23090
rect 2175 23025 2255 23030
rect 2575 23200 2655 23205
rect 2575 23140 2585 23200
rect 2645 23140 2655 23200
rect 2575 23090 2655 23140
rect 2575 23030 2585 23090
rect 2645 23030 2655 23090
rect 2575 23025 2655 23030
rect 2975 23200 3055 23205
rect 2975 23140 2985 23200
rect 3045 23140 3055 23200
rect 2975 23090 3055 23140
rect 2975 23030 2985 23090
rect 3045 23030 3055 23090
rect 2975 23025 3055 23030
rect 3375 23200 3455 23205
rect 3375 23140 3385 23200
rect 3445 23140 3455 23200
rect 3375 23090 3455 23140
rect 3375 23030 3385 23090
rect 3445 23030 3455 23090
rect 3375 23025 3455 23030
rect 3775 23200 3855 23205
rect 3775 23140 3785 23200
rect 3845 23140 3855 23200
rect 3775 23090 3855 23140
rect 3775 23030 3785 23090
rect 3845 23030 3855 23090
rect 3775 23025 3855 23030
rect 4175 23200 4255 23205
rect 4175 23140 4185 23200
rect 4245 23140 4255 23200
rect 4175 23090 4255 23140
rect 4175 23030 4185 23090
rect 4245 23030 4255 23090
rect 4175 23025 4255 23030
rect 4575 23200 4655 23205
rect 4575 23140 4585 23200
rect 4645 23140 4655 23200
rect 4575 23090 4655 23140
rect 4575 23030 4585 23090
rect 4645 23030 4655 23090
rect 4575 23025 4655 23030
rect 4975 23200 5055 23205
rect 4975 23140 4985 23200
rect 5045 23140 5055 23200
rect 4975 23090 5055 23140
rect 4975 23030 4985 23090
rect 5045 23030 5055 23090
rect 4975 23025 5055 23030
rect 5375 23200 5455 23205
rect 5375 23140 5385 23200
rect 5445 23140 5455 23200
rect 5375 23090 5455 23140
rect 5375 23030 5385 23090
rect 5445 23030 5455 23090
rect 5375 23025 5455 23030
rect 5775 23200 5855 23205
rect 5775 23140 5785 23200
rect 5845 23140 5855 23200
rect 5775 23090 5855 23140
rect 5775 23030 5785 23090
rect 5845 23030 5855 23090
rect 5775 23025 5855 23030
rect 6175 23200 6255 23205
rect 6175 23140 6185 23200
rect 6245 23140 6255 23200
rect 6175 23090 6255 23140
rect 6175 23030 6185 23090
rect 6245 23030 6255 23090
rect 6175 23025 6255 23030
rect 6575 23200 6655 23205
rect 6575 23140 6585 23200
rect 6645 23140 6655 23200
rect 6575 23090 6655 23140
rect 6575 23030 6585 23090
rect 6645 23030 6655 23090
rect 6575 23025 6655 23030
rect 6975 23200 7055 23205
rect 6975 23140 6985 23200
rect 7045 23140 7055 23200
rect 6975 23090 7055 23140
rect 6975 23030 6985 23090
rect 7045 23030 7055 23090
rect 6975 23025 7055 23030
rect 7375 23200 7455 23205
rect 7375 23140 7385 23200
rect 7445 23140 7455 23200
rect 7375 23090 7455 23140
rect 7375 23030 7385 23090
rect 7445 23030 7455 23090
rect 7375 23025 7455 23030
rect 7775 23200 7855 23205
rect 7775 23140 7785 23200
rect 7845 23140 7855 23200
rect 7775 23090 7855 23140
rect 7775 23030 7785 23090
rect 7845 23030 7855 23090
rect 7775 23025 7855 23030
rect 8175 23200 8255 23205
rect 8175 23140 8185 23200
rect 8245 23140 8255 23200
rect 8175 23090 8255 23140
rect 8175 23030 8185 23090
rect 8245 23030 8255 23090
rect 8175 23025 8255 23030
rect 8575 23200 8655 23205
rect 8575 23140 8585 23200
rect 8645 23140 8655 23200
rect 8575 23090 8655 23140
rect 8575 23030 8585 23090
rect 8645 23030 8655 23090
rect 8575 23025 8655 23030
rect 8975 23200 9055 23205
rect 8975 23140 8985 23200
rect 9045 23140 9055 23200
rect 8975 23090 9055 23140
rect 8975 23030 8985 23090
rect 9045 23030 9055 23090
rect 8975 23025 9055 23030
rect 9375 23200 9455 23205
rect 9375 23140 9385 23200
rect 9445 23140 9455 23200
rect 9375 23090 9455 23140
rect 9375 23030 9385 23090
rect 9445 23030 9455 23090
rect 9375 23025 9455 23030
rect 9775 23200 9855 23205
rect 9775 23140 9785 23200
rect 9845 23140 9855 23200
rect 9775 23090 9855 23140
rect 9775 23030 9785 23090
rect 9845 23030 9855 23090
rect 9775 23025 9855 23030
rect 10175 23200 10255 23205
rect 10175 23140 10185 23200
rect 10245 23140 10255 23200
rect 10175 23090 10255 23140
rect 10175 23030 10185 23090
rect 10245 23030 10255 23090
rect 10175 23025 10255 23030
rect 10575 23200 10655 23205
rect 10575 23140 10585 23200
rect 10645 23140 10655 23200
rect 10575 23090 10655 23140
rect 10575 23030 10585 23090
rect 10645 23030 10655 23090
rect 10575 23025 10655 23030
rect 10975 23200 11055 23205
rect 10975 23140 10985 23200
rect 11045 23140 11055 23200
rect 10975 23090 11055 23140
rect 10975 23030 10985 23090
rect 11045 23030 11055 23090
rect 10975 23025 11055 23030
rect 11375 23200 11455 23205
rect 11375 23140 11385 23200
rect 11445 23140 11455 23200
rect 11375 23090 11455 23140
rect 11375 23030 11385 23090
rect 11445 23030 11455 23090
rect 11375 23025 11455 23030
rect 11775 23200 11855 23205
rect 11775 23140 11785 23200
rect 11845 23140 11855 23200
rect 11775 23090 11855 23140
rect 11775 23030 11785 23090
rect 11845 23030 11855 23090
rect 11775 23025 11855 23030
rect 12175 23200 12255 23205
rect 12175 23140 12185 23200
rect 12245 23140 12255 23200
rect 12175 23090 12255 23140
rect 12175 23030 12185 23090
rect 12245 23030 12255 23090
rect 12175 23025 12255 23030
rect 12575 23200 12655 23205
rect 12575 23140 12585 23200
rect 12645 23140 12655 23200
rect 12575 23090 12655 23140
rect 12575 23030 12585 23090
rect 12645 23030 12655 23090
rect 12575 23025 12655 23030
rect 12975 23200 13055 23205
rect 12975 23140 12985 23200
rect 13045 23140 13055 23200
rect 12975 23090 13055 23140
rect 12975 23030 12985 23090
rect 13045 23030 13055 23090
rect 12975 23025 13055 23030
rect -215 22835 -155 23025
rect 185 22835 245 23025
rect 585 22835 645 23025
rect 985 22835 1045 23025
rect 1385 22835 1445 23025
rect 1785 22835 1845 23025
rect 2185 22835 2245 23025
rect 2585 22835 2645 23025
rect 2985 22835 3045 23025
rect 3385 22835 3445 23025
rect 3785 22835 3845 23025
rect 4185 22835 4245 23025
rect 4585 22835 4645 23025
rect 4985 22835 5045 23025
rect 5385 22835 5445 23025
rect 5785 22835 5845 23025
rect 6185 22835 6245 23025
rect 6585 22835 6645 23025
rect 6985 22835 7045 23025
rect 7385 22835 7445 23025
rect 7785 22835 7845 23025
rect 8185 22835 8245 23025
rect 8585 22835 8645 23025
rect 8985 22835 9045 23025
rect 9385 22835 9445 23025
rect 9785 22835 9845 23025
rect 10185 22835 10245 23025
rect 10585 22835 10645 23025
rect 10985 22835 11045 23025
rect 11385 22835 11445 23025
rect 11785 22835 11845 23025
rect 12185 22835 12245 23025
rect 12585 22835 12645 23025
rect 12985 22835 13045 23025
rect -225 22830 -145 22835
rect -225 22770 -215 22830
rect -155 22770 -145 22830
rect -225 22720 -145 22770
rect -225 22660 -215 22720
rect -155 22660 -145 22720
rect -225 22655 -145 22660
rect 175 22830 255 22835
rect 175 22770 185 22830
rect 245 22770 255 22830
rect 175 22720 255 22770
rect 175 22660 185 22720
rect 245 22660 255 22720
rect 175 22655 255 22660
rect 575 22830 655 22835
rect 575 22770 585 22830
rect 645 22770 655 22830
rect 575 22720 655 22770
rect 575 22660 585 22720
rect 645 22660 655 22720
rect 575 22655 655 22660
rect 975 22830 1055 22835
rect 975 22770 985 22830
rect 1045 22770 1055 22830
rect 975 22720 1055 22770
rect 975 22660 985 22720
rect 1045 22660 1055 22720
rect 975 22655 1055 22660
rect 1375 22830 1455 22835
rect 1375 22770 1385 22830
rect 1445 22770 1455 22830
rect 1375 22720 1455 22770
rect 1375 22660 1385 22720
rect 1445 22660 1455 22720
rect 1375 22655 1455 22660
rect 1775 22830 1855 22835
rect 1775 22770 1785 22830
rect 1845 22770 1855 22830
rect 1775 22720 1855 22770
rect 1775 22660 1785 22720
rect 1845 22660 1855 22720
rect 1775 22655 1855 22660
rect 2175 22830 2255 22835
rect 2175 22770 2185 22830
rect 2245 22770 2255 22830
rect 2175 22720 2255 22770
rect 2175 22660 2185 22720
rect 2245 22660 2255 22720
rect 2175 22655 2255 22660
rect 2575 22830 2655 22835
rect 2575 22770 2585 22830
rect 2645 22770 2655 22830
rect 2575 22720 2655 22770
rect 2575 22660 2585 22720
rect 2645 22660 2655 22720
rect 2575 22655 2655 22660
rect 2975 22830 3055 22835
rect 2975 22770 2985 22830
rect 3045 22770 3055 22830
rect 2975 22720 3055 22770
rect 2975 22660 2985 22720
rect 3045 22660 3055 22720
rect 2975 22655 3055 22660
rect 3375 22830 3455 22835
rect 3375 22770 3385 22830
rect 3445 22770 3455 22830
rect 3375 22720 3455 22770
rect 3375 22660 3385 22720
rect 3445 22660 3455 22720
rect 3375 22655 3455 22660
rect 3775 22830 3855 22835
rect 3775 22770 3785 22830
rect 3845 22770 3855 22830
rect 3775 22720 3855 22770
rect 3775 22660 3785 22720
rect 3845 22660 3855 22720
rect 3775 22655 3855 22660
rect 4175 22830 4255 22835
rect 4175 22770 4185 22830
rect 4245 22770 4255 22830
rect 4175 22720 4255 22770
rect 4175 22660 4185 22720
rect 4245 22660 4255 22720
rect 4175 22655 4255 22660
rect 4575 22830 4655 22835
rect 4575 22770 4585 22830
rect 4645 22770 4655 22830
rect 4575 22720 4655 22770
rect 4575 22660 4585 22720
rect 4645 22660 4655 22720
rect 4575 22655 4655 22660
rect 4975 22830 5055 22835
rect 4975 22770 4985 22830
rect 5045 22770 5055 22830
rect 4975 22720 5055 22770
rect 4975 22660 4985 22720
rect 5045 22660 5055 22720
rect 4975 22655 5055 22660
rect 5375 22830 5455 22835
rect 5375 22770 5385 22830
rect 5445 22770 5455 22830
rect 5375 22720 5455 22770
rect 5375 22660 5385 22720
rect 5445 22660 5455 22720
rect 5375 22655 5455 22660
rect 5775 22830 5855 22835
rect 5775 22770 5785 22830
rect 5845 22770 5855 22830
rect 5775 22720 5855 22770
rect 5775 22660 5785 22720
rect 5845 22660 5855 22720
rect 5775 22655 5855 22660
rect 6175 22830 6255 22835
rect 6175 22770 6185 22830
rect 6245 22770 6255 22830
rect 6175 22720 6255 22770
rect 6175 22660 6185 22720
rect 6245 22660 6255 22720
rect 6175 22655 6255 22660
rect 6575 22830 6655 22835
rect 6575 22770 6585 22830
rect 6645 22770 6655 22830
rect 6575 22720 6655 22770
rect 6575 22660 6585 22720
rect 6645 22660 6655 22720
rect 6575 22655 6655 22660
rect 6975 22830 7055 22835
rect 6975 22770 6985 22830
rect 7045 22770 7055 22830
rect 6975 22720 7055 22770
rect 6975 22660 6985 22720
rect 7045 22660 7055 22720
rect 6975 22655 7055 22660
rect 7375 22830 7455 22835
rect 7375 22770 7385 22830
rect 7445 22770 7455 22830
rect 7375 22720 7455 22770
rect 7375 22660 7385 22720
rect 7445 22660 7455 22720
rect 7375 22655 7455 22660
rect 7775 22830 7855 22835
rect 7775 22770 7785 22830
rect 7845 22770 7855 22830
rect 7775 22720 7855 22770
rect 7775 22660 7785 22720
rect 7845 22660 7855 22720
rect 7775 22655 7855 22660
rect 8175 22830 8255 22835
rect 8175 22770 8185 22830
rect 8245 22770 8255 22830
rect 8175 22720 8255 22770
rect 8175 22660 8185 22720
rect 8245 22660 8255 22720
rect 8175 22655 8255 22660
rect 8575 22830 8655 22835
rect 8575 22770 8585 22830
rect 8645 22770 8655 22830
rect 8575 22720 8655 22770
rect 8575 22660 8585 22720
rect 8645 22660 8655 22720
rect 8575 22655 8655 22660
rect 8975 22830 9055 22835
rect 8975 22770 8985 22830
rect 9045 22770 9055 22830
rect 8975 22720 9055 22770
rect 8975 22660 8985 22720
rect 9045 22660 9055 22720
rect 8975 22655 9055 22660
rect 9375 22830 9455 22835
rect 9375 22770 9385 22830
rect 9445 22770 9455 22830
rect 9375 22720 9455 22770
rect 9375 22660 9385 22720
rect 9445 22660 9455 22720
rect 9375 22655 9455 22660
rect 9775 22830 9855 22835
rect 9775 22770 9785 22830
rect 9845 22770 9855 22830
rect 9775 22720 9855 22770
rect 9775 22660 9785 22720
rect 9845 22660 9855 22720
rect 9775 22655 9855 22660
rect 10175 22830 10255 22835
rect 10175 22770 10185 22830
rect 10245 22770 10255 22830
rect 10175 22720 10255 22770
rect 10175 22660 10185 22720
rect 10245 22660 10255 22720
rect 10175 22655 10255 22660
rect 10575 22830 10655 22835
rect 10575 22770 10585 22830
rect 10645 22770 10655 22830
rect 10575 22720 10655 22770
rect 10575 22660 10585 22720
rect 10645 22660 10655 22720
rect 10575 22655 10655 22660
rect 10975 22830 11055 22835
rect 10975 22770 10985 22830
rect 11045 22770 11055 22830
rect 10975 22720 11055 22770
rect 10975 22660 10985 22720
rect 11045 22660 11055 22720
rect 10975 22655 11055 22660
rect 11375 22830 11455 22835
rect 11375 22770 11385 22830
rect 11445 22770 11455 22830
rect 11375 22720 11455 22770
rect 11375 22660 11385 22720
rect 11445 22660 11455 22720
rect 11375 22655 11455 22660
rect 11775 22830 11855 22835
rect 11775 22770 11785 22830
rect 11845 22770 11855 22830
rect 11775 22720 11855 22770
rect 11775 22660 11785 22720
rect 11845 22660 11855 22720
rect 11775 22655 11855 22660
rect 12175 22830 12255 22835
rect 12175 22770 12185 22830
rect 12245 22770 12255 22830
rect 12175 22720 12255 22770
rect 12175 22660 12185 22720
rect 12245 22660 12255 22720
rect 12175 22655 12255 22660
rect 12575 22830 12655 22835
rect 12575 22770 12585 22830
rect 12645 22770 12655 22830
rect 12575 22720 12655 22770
rect 12575 22660 12585 22720
rect 12645 22660 12655 22720
rect 12575 22655 12655 22660
rect 12975 22830 13055 22835
rect 12975 22770 12985 22830
rect 13045 22770 13055 22830
rect 12975 22720 13055 22770
rect 12975 22660 12985 22720
rect 13045 22660 13055 22720
rect 12975 22655 13055 22660
rect -215 22465 -155 22655
rect 185 22465 245 22655
rect 585 22465 645 22655
rect 985 22465 1045 22655
rect 1385 22465 1445 22655
rect 1785 22465 1845 22655
rect 2185 22465 2245 22655
rect 2585 22465 2645 22655
rect 2985 22465 3045 22655
rect 3385 22465 3445 22655
rect 3785 22465 3845 22655
rect 4185 22465 4245 22655
rect 4585 22465 4645 22655
rect 4985 22465 5045 22655
rect 5385 22465 5445 22655
rect 5785 22465 5845 22655
rect 6185 22465 6245 22655
rect 6585 22465 6645 22655
rect 6985 22465 7045 22655
rect 7385 22465 7445 22655
rect 7785 22465 7845 22655
rect 8185 22465 8245 22655
rect 8585 22465 8645 22655
rect 8985 22465 9045 22655
rect 9385 22465 9445 22655
rect 9785 22465 9845 22655
rect 10185 22465 10245 22655
rect 10585 22465 10645 22655
rect 10985 22465 11045 22655
rect 11385 22465 11445 22655
rect 11785 22465 11845 22655
rect 12185 22465 12245 22655
rect 12585 22465 12645 22655
rect 12985 22465 13045 22655
rect -225 22460 -145 22465
rect -225 22400 -215 22460
rect -155 22400 -145 22460
rect -225 22350 -145 22400
rect -225 22290 -215 22350
rect -155 22290 -145 22350
rect -225 22285 -145 22290
rect 175 22460 255 22465
rect 175 22400 185 22460
rect 245 22400 255 22460
rect 175 22350 255 22400
rect 175 22290 185 22350
rect 245 22290 255 22350
rect 175 22285 255 22290
rect 575 22460 655 22465
rect 575 22400 585 22460
rect 645 22400 655 22460
rect 575 22350 655 22400
rect 575 22290 585 22350
rect 645 22290 655 22350
rect 575 22285 655 22290
rect 975 22460 1055 22465
rect 975 22400 985 22460
rect 1045 22400 1055 22460
rect 975 22350 1055 22400
rect 975 22290 985 22350
rect 1045 22290 1055 22350
rect 975 22285 1055 22290
rect 1375 22460 1455 22465
rect 1375 22400 1385 22460
rect 1445 22400 1455 22460
rect 1375 22350 1455 22400
rect 1375 22290 1385 22350
rect 1445 22290 1455 22350
rect 1375 22285 1455 22290
rect 1775 22460 1855 22465
rect 1775 22400 1785 22460
rect 1845 22400 1855 22460
rect 1775 22350 1855 22400
rect 1775 22290 1785 22350
rect 1845 22290 1855 22350
rect 1775 22285 1855 22290
rect 2175 22460 2255 22465
rect 2175 22400 2185 22460
rect 2245 22400 2255 22460
rect 2175 22350 2255 22400
rect 2175 22290 2185 22350
rect 2245 22290 2255 22350
rect 2175 22285 2255 22290
rect 2575 22460 2655 22465
rect 2575 22400 2585 22460
rect 2645 22400 2655 22460
rect 2575 22350 2655 22400
rect 2575 22290 2585 22350
rect 2645 22290 2655 22350
rect 2575 22285 2655 22290
rect 2975 22460 3055 22465
rect 2975 22400 2985 22460
rect 3045 22400 3055 22460
rect 2975 22350 3055 22400
rect 2975 22290 2985 22350
rect 3045 22290 3055 22350
rect 2975 22285 3055 22290
rect 3375 22460 3455 22465
rect 3375 22400 3385 22460
rect 3445 22400 3455 22460
rect 3375 22350 3455 22400
rect 3375 22290 3385 22350
rect 3445 22290 3455 22350
rect 3375 22285 3455 22290
rect 3775 22460 3855 22465
rect 3775 22400 3785 22460
rect 3845 22400 3855 22460
rect 3775 22350 3855 22400
rect 3775 22290 3785 22350
rect 3845 22290 3855 22350
rect 3775 22285 3855 22290
rect 4175 22460 4255 22465
rect 4175 22400 4185 22460
rect 4245 22400 4255 22460
rect 4175 22350 4255 22400
rect 4175 22290 4185 22350
rect 4245 22290 4255 22350
rect 4175 22285 4255 22290
rect 4575 22460 4655 22465
rect 4575 22400 4585 22460
rect 4645 22400 4655 22460
rect 4575 22350 4655 22400
rect 4575 22290 4585 22350
rect 4645 22290 4655 22350
rect 4575 22285 4655 22290
rect 4975 22460 5055 22465
rect 4975 22400 4985 22460
rect 5045 22400 5055 22460
rect 4975 22350 5055 22400
rect 4975 22290 4985 22350
rect 5045 22290 5055 22350
rect 4975 22285 5055 22290
rect 5375 22460 5455 22465
rect 5375 22400 5385 22460
rect 5445 22400 5455 22460
rect 5375 22350 5455 22400
rect 5375 22290 5385 22350
rect 5445 22290 5455 22350
rect 5375 22285 5455 22290
rect 5775 22460 5855 22465
rect 5775 22400 5785 22460
rect 5845 22400 5855 22460
rect 5775 22350 5855 22400
rect 5775 22290 5785 22350
rect 5845 22290 5855 22350
rect 5775 22285 5855 22290
rect 6175 22460 6255 22465
rect 6175 22400 6185 22460
rect 6245 22400 6255 22460
rect 6175 22350 6255 22400
rect 6175 22290 6185 22350
rect 6245 22290 6255 22350
rect 6175 22285 6255 22290
rect 6575 22460 6655 22465
rect 6575 22400 6585 22460
rect 6645 22400 6655 22460
rect 6575 22350 6655 22400
rect 6575 22290 6585 22350
rect 6645 22290 6655 22350
rect 6575 22285 6655 22290
rect 6975 22460 7055 22465
rect 6975 22400 6985 22460
rect 7045 22400 7055 22460
rect 6975 22350 7055 22400
rect 6975 22290 6985 22350
rect 7045 22290 7055 22350
rect 6975 22285 7055 22290
rect 7375 22460 7455 22465
rect 7375 22400 7385 22460
rect 7445 22400 7455 22460
rect 7375 22350 7455 22400
rect 7375 22290 7385 22350
rect 7445 22290 7455 22350
rect 7375 22285 7455 22290
rect 7775 22460 7855 22465
rect 7775 22400 7785 22460
rect 7845 22400 7855 22460
rect 7775 22350 7855 22400
rect 7775 22290 7785 22350
rect 7845 22290 7855 22350
rect 7775 22285 7855 22290
rect 8175 22460 8255 22465
rect 8175 22400 8185 22460
rect 8245 22400 8255 22460
rect 8175 22350 8255 22400
rect 8175 22290 8185 22350
rect 8245 22290 8255 22350
rect 8175 22285 8255 22290
rect 8575 22460 8655 22465
rect 8575 22400 8585 22460
rect 8645 22400 8655 22460
rect 8575 22350 8655 22400
rect 8575 22290 8585 22350
rect 8645 22290 8655 22350
rect 8575 22285 8655 22290
rect 8975 22460 9055 22465
rect 8975 22400 8985 22460
rect 9045 22400 9055 22460
rect 8975 22350 9055 22400
rect 8975 22290 8985 22350
rect 9045 22290 9055 22350
rect 8975 22285 9055 22290
rect 9375 22460 9455 22465
rect 9375 22400 9385 22460
rect 9445 22400 9455 22460
rect 9375 22350 9455 22400
rect 9375 22290 9385 22350
rect 9445 22290 9455 22350
rect 9375 22285 9455 22290
rect 9775 22460 9855 22465
rect 9775 22400 9785 22460
rect 9845 22400 9855 22460
rect 9775 22350 9855 22400
rect 9775 22290 9785 22350
rect 9845 22290 9855 22350
rect 9775 22285 9855 22290
rect 10175 22460 10255 22465
rect 10175 22400 10185 22460
rect 10245 22400 10255 22460
rect 10175 22350 10255 22400
rect 10175 22290 10185 22350
rect 10245 22290 10255 22350
rect 10175 22285 10255 22290
rect 10575 22460 10655 22465
rect 10575 22400 10585 22460
rect 10645 22400 10655 22460
rect 10575 22350 10655 22400
rect 10575 22290 10585 22350
rect 10645 22290 10655 22350
rect 10575 22285 10655 22290
rect 10975 22460 11055 22465
rect 10975 22400 10985 22460
rect 11045 22400 11055 22460
rect 10975 22350 11055 22400
rect 10975 22290 10985 22350
rect 11045 22290 11055 22350
rect 10975 22285 11055 22290
rect 11375 22460 11455 22465
rect 11375 22400 11385 22460
rect 11445 22400 11455 22460
rect 11375 22350 11455 22400
rect 11375 22290 11385 22350
rect 11445 22290 11455 22350
rect 11375 22285 11455 22290
rect 11775 22460 11855 22465
rect 11775 22400 11785 22460
rect 11845 22400 11855 22460
rect 11775 22350 11855 22400
rect 11775 22290 11785 22350
rect 11845 22290 11855 22350
rect 11775 22285 11855 22290
rect 12175 22460 12255 22465
rect 12175 22400 12185 22460
rect 12245 22400 12255 22460
rect 12175 22350 12255 22400
rect 12175 22290 12185 22350
rect 12245 22290 12255 22350
rect 12175 22285 12255 22290
rect 12575 22460 12655 22465
rect 12575 22400 12585 22460
rect 12645 22400 12655 22460
rect 12575 22350 12655 22400
rect 12575 22290 12585 22350
rect 12645 22290 12655 22350
rect 12575 22285 12655 22290
rect 12975 22460 13055 22465
rect 12975 22400 12985 22460
rect 13045 22400 13055 22460
rect 12975 22350 13055 22400
rect 12975 22290 12985 22350
rect 13045 22290 13055 22350
rect 12975 22285 13055 22290
rect -215 22095 -155 22285
rect 185 22095 245 22285
rect 585 22095 645 22285
rect 985 22095 1045 22285
rect 1385 22095 1445 22285
rect 1785 22095 1845 22285
rect 2185 22095 2245 22285
rect 2585 22095 2645 22285
rect 2985 22095 3045 22285
rect 3385 22095 3445 22285
rect 3785 22095 3845 22285
rect 4185 22095 4245 22285
rect 4585 22095 4645 22285
rect 4985 22095 5045 22285
rect 5385 22095 5445 22285
rect 5785 22095 5845 22285
rect 6185 22095 6245 22285
rect 6585 22095 6645 22285
rect 6985 22095 7045 22285
rect 7385 22095 7445 22285
rect 7785 22095 7845 22285
rect 8185 22095 8245 22285
rect 8585 22095 8645 22285
rect 8985 22095 9045 22285
rect 9385 22095 9445 22285
rect 9785 22095 9845 22285
rect 10185 22095 10245 22285
rect 10585 22095 10645 22285
rect 10985 22095 11045 22285
rect 11385 22095 11445 22285
rect 11785 22095 11845 22285
rect 12185 22095 12245 22285
rect 12585 22095 12645 22285
rect 12985 22095 13045 22285
rect -225 22090 -145 22095
rect -225 22030 -215 22090
rect -155 22030 -145 22090
rect -225 21980 -145 22030
rect -225 21920 -215 21980
rect -155 21920 -145 21980
rect -225 21915 -145 21920
rect 175 22090 255 22095
rect 175 22030 185 22090
rect 245 22030 255 22090
rect 175 21980 255 22030
rect 175 21920 185 21980
rect 245 21920 255 21980
rect 175 21915 255 21920
rect 575 22090 655 22095
rect 575 22030 585 22090
rect 645 22030 655 22090
rect 575 21980 655 22030
rect 575 21920 585 21980
rect 645 21920 655 21980
rect 575 21915 655 21920
rect 975 22090 1055 22095
rect 975 22030 985 22090
rect 1045 22030 1055 22090
rect 975 21980 1055 22030
rect 975 21920 985 21980
rect 1045 21920 1055 21980
rect 975 21915 1055 21920
rect 1375 22090 1455 22095
rect 1375 22030 1385 22090
rect 1445 22030 1455 22090
rect 1375 21980 1455 22030
rect 1375 21920 1385 21980
rect 1445 21920 1455 21980
rect 1375 21915 1455 21920
rect 1775 22090 1855 22095
rect 1775 22030 1785 22090
rect 1845 22030 1855 22090
rect 1775 21980 1855 22030
rect 1775 21920 1785 21980
rect 1845 21920 1855 21980
rect 1775 21915 1855 21920
rect 2175 22090 2255 22095
rect 2175 22030 2185 22090
rect 2245 22030 2255 22090
rect 2175 21980 2255 22030
rect 2175 21920 2185 21980
rect 2245 21920 2255 21980
rect 2175 21915 2255 21920
rect 2575 22090 2655 22095
rect 2575 22030 2585 22090
rect 2645 22030 2655 22090
rect 2575 21980 2655 22030
rect 2575 21920 2585 21980
rect 2645 21920 2655 21980
rect 2575 21915 2655 21920
rect 2975 22090 3055 22095
rect 2975 22030 2985 22090
rect 3045 22030 3055 22090
rect 2975 21980 3055 22030
rect 2975 21920 2985 21980
rect 3045 21920 3055 21980
rect 2975 21915 3055 21920
rect 3375 22090 3455 22095
rect 3375 22030 3385 22090
rect 3445 22030 3455 22090
rect 3375 21980 3455 22030
rect 3375 21920 3385 21980
rect 3445 21920 3455 21980
rect 3375 21915 3455 21920
rect 3775 22090 3855 22095
rect 3775 22030 3785 22090
rect 3845 22030 3855 22090
rect 3775 21980 3855 22030
rect 3775 21920 3785 21980
rect 3845 21920 3855 21980
rect 3775 21915 3855 21920
rect 4175 22090 4255 22095
rect 4175 22030 4185 22090
rect 4245 22030 4255 22090
rect 4175 21980 4255 22030
rect 4175 21920 4185 21980
rect 4245 21920 4255 21980
rect 4175 21915 4255 21920
rect 4575 22090 4655 22095
rect 4575 22030 4585 22090
rect 4645 22030 4655 22090
rect 4575 21980 4655 22030
rect 4575 21920 4585 21980
rect 4645 21920 4655 21980
rect 4575 21915 4655 21920
rect 4975 22090 5055 22095
rect 4975 22030 4985 22090
rect 5045 22030 5055 22090
rect 4975 21980 5055 22030
rect 4975 21920 4985 21980
rect 5045 21920 5055 21980
rect 4975 21915 5055 21920
rect 5375 22090 5455 22095
rect 5375 22030 5385 22090
rect 5445 22030 5455 22090
rect 5375 21980 5455 22030
rect 5375 21920 5385 21980
rect 5445 21920 5455 21980
rect 5375 21915 5455 21920
rect 5775 22090 5855 22095
rect 5775 22030 5785 22090
rect 5845 22030 5855 22090
rect 5775 21980 5855 22030
rect 5775 21920 5785 21980
rect 5845 21920 5855 21980
rect 5775 21915 5855 21920
rect 6175 22090 6255 22095
rect 6175 22030 6185 22090
rect 6245 22030 6255 22090
rect 6175 21980 6255 22030
rect 6175 21920 6185 21980
rect 6245 21920 6255 21980
rect 6175 21915 6255 21920
rect 6575 22090 6655 22095
rect 6575 22030 6585 22090
rect 6645 22030 6655 22090
rect 6575 21980 6655 22030
rect 6575 21920 6585 21980
rect 6645 21920 6655 21980
rect 6575 21915 6655 21920
rect 6975 22090 7055 22095
rect 6975 22030 6985 22090
rect 7045 22030 7055 22090
rect 6975 21980 7055 22030
rect 6975 21920 6985 21980
rect 7045 21920 7055 21980
rect 6975 21915 7055 21920
rect 7375 22090 7455 22095
rect 7375 22030 7385 22090
rect 7445 22030 7455 22090
rect 7375 21980 7455 22030
rect 7375 21920 7385 21980
rect 7445 21920 7455 21980
rect 7375 21915 7455 21920
rect 7775 22090 7855 22095
rect 7775 22030 7785 22090
rect 7845 22030 7855 22090
rect 7775 21980 7855 22030
rect 7775 21920 7785 21980
rect 7845 21920 7855 21980
rect 7775 21915 7855 21920
rect 8175 22090 8255 22095
rect 8175 22030 8185 22090
rect 8245 22030 8255 22090
rect 8175 21980 8255 22030
rect 8175 21920 8185 21980
rect 8245 21920 8255 21980
rect 8175 21915 8255 21920
rect 8575 22090 8655 22095
rect 8575 22030 8585 22090
rect 8645 22030 8655 22090
rect 8575 21980 8655 22030
rect 8575 21920 8585 21980
rect 8645 21920 8655 21980
rect 8575 21915 8655 21920
rect 8975 22090 9055 22095
rect 8975 22030 8985 22090
rect 9045 22030 9055 22090
rect 8975 21980 9055 22030
rect 8975 21920 8985 21980
rect 9045 21920 9055 21980
rect 8975 21915 9055 21920
rect 9375 22090 9455 22095
rect 9375 22030 9385 22090
rect 9445 22030 9455 22090
rect 9375 21980 9455 22030
rect 9375 21920 9385 21980
rect 9445 21920 9455 21980
rect 9375 21915 9455 21920
rect 9775 22090 9855 22095
rect 9775 22030 9785 22090
rect 9845 22030 9855 22090
rect 9775 21980 9855 22030
rect 9775 21920 9785 21980
rect 9845 21920 9855 21980
rect 9775 21915 9855 21920
rect 10175 22090 10255 22095
rect 10175 22030 10185 22090
rect 10245 22030 10255 22090
rect 10175 21980 10255 22030
rect 10175 21920 10185 21980
rect 10245 21920 10255 21980
rect 10175 21915 10255 21920
rect 10575 22090 10655 22095
rect 10575 22030 10585 22090
rect 10645 22030 10655 22090
rect 10575 21980 10655 22030
rect 10575 21920 10585 21980
rect 10645 21920 10655 21980
rect 10575 21915 10655 21920
rect 10975 22090 11055 22095
rect 10975 22030 10985 22090
rect 11045 22030 11055 22090
rect 10975 21980 11055 22030
rect 10975 21920 10985 21980
rect 11045 21920 11055 21980
rect 10975 21915 11055 21920
rect 11375 22090 11455 22095
rect 11375 22030 11385 22090
rect 11445 22030 11455 22090
rect 11375 21980 11455 22030
rect 11375 21920 11385 21980
rect 11445 21920 11455 21980
rect 11375 21915 11455 21920
rect 11775 22090 11855 22095
rect 11775 22030 11785 22090
rect 11845 22030 11855 22090
rect 11775 21980 11855 22030
rect 11775 21920 11785 21980
rect 11845 21920 11855 21980
rect 11775 21915 11855 21920
rect 12175 22090 12255 22095
rect 12175 22030 12185 22090
rect 12245 22030 12255 22090
rect 12175 21980 12255 22030
rect 12175 21920 12185 21980
rect 12245 21920 12255 21980
rect 12175 21915 12255 21920
rect 12575 22090 12655 22095
rect 12575 22030 12585 22090
rect 12645 22030 12655 22090
rect 12575 21980 12655 22030
rect 12575 21920 12585 21980
rect 12645 21920 12655 21980
rect 12575 21915 12655 21920
rect 12975 22090 13055 22095
rect 12975 22030 12985 22090
rect 13045 22030 13055 22090
rect 12975 21980 13055 22030
rect 12975 21920 12985 21980
rect 13045 21920 13055 21980
rect 12975 21915 13055 21920
rect -215 21725 -155 21915
rect 185 21725 245 21915
rect 585 21725 645 21915
rect 985 21725 1045 21915
rect 1385 21725 1445 21915
rect 1785 21725 1845 21915
rect 2185 21725 2245 21915
rect 2585 21725 2645 21915
rect 2985 21725 3045 21915
rect 3385 21725 3445 21915
rect 3785 21725 3845 21915
rect 4185 21725 4245 21915
rect 4585 21725 4645 21915
rect 4985 21725 5045 21915
rect 5385 21725 5445 21915
rect 5785 21725 5845 21915
rect 6185 21725 6245 21915
rect 6585 21725 6645 21915
rect 6985 21725 7045 21915
rect 7385 21725 7445 21915
rect 7785 21725 7845 21915
rect 8185 21725 8245 21915
rect 8585 21725 8645 21915
rect 8985 21725 9045 21915
rect 9385 21725 9445 21915
rect 9785 21725 9845 21915
rect 10185 21725 10245 21915
rect 10585 21725 10645 21915
rect 10985 21725 11045 21915
rect 11385 21725 11445 21915
rect 11785 21725 11845 21915
rect 12185 21725 12245 21915
rect 12585 21725 12645 21915
rect 12985 21725 13045 21915
rect -225 21720 -145 21725
rect -225 21660 -215 21720
rect -155 21660 -145 21720
rect -225 21610 -145 21660
rect -225 21550 -215 21610
rect -155 21550 -145 21610
rect -225 21545 -145 21550
rect 175 21720 255 21725
rect 175 21660 185 21720
rect 245 21660 255 21720
rect 175 21610 255 21660
rect 175 21550 185 21610
rect 245 21550 255 21610
rect 175 21545 255 21550
rect 575 21720 655 21725
rect 575 21660 585 21720
rect 645 21660 655 21720
rect 575 21610 655 21660
rect 575 21550 585 21610
rect 645 21550 655 21610
rect 575 21545 655 21550
rect 975 21720 1055 21725
rect 975 21660 985 21720
rect 1045 21660 1055 21720
rect 975 21610 1055 21660
rect 975 21550 985 21610
rect 1045 21550 1055 21610
rect 975 21545 1055 21550
rect 1375 21720 1455 21725
rect 1375 21660 1385 21720
rect 1445 21660 1455 21720
rect 1375 21610 1455 21660
rect 1375 21550 1385 21610
rect 1445 21550 1455 21610
rect 1375 21545 1455 21550
rect 1775 21720 1855 21725
rect 1775 21660 1785 21720
rect 1845 21660 1855 21720
rect 1775 21610 1855 21660
rect 1775 21550 1785 21610
rect 1845 21550 1855 21610
rect 1775 21545 1855 21550
rect 2175 21720 2255 21725
rect 2175 21660 2185 21720
rect 2245 21660 2255 21720
rect 2175 21610 2255 21660
rect 2175 21550 2185 21610
rect 2245 21550 2255 21610
rect 2175 21545 2255 21550
rect 2575 21720 2655 21725
rect 2575 21660 2585 21720
rect 2645 21660 2655 21720
rect 2575 21610 2655 21660
rect 2575 21550 2585 21610
rect 2645 21550 2655 21610
rect 2575 21545 2655 21550
rect 2975 21720 3055 21725
rect 2975 21660 2985 21720
rect 3045 21660 3055 21720
rect 2975 21610 3055 21660
rect 2975 21550 2985 21610
rect 3045 21550 3055 21610
rect 2975 21545 3055 21550
rect 3375 21720 3455 21725
rect 3375 21660 3385 21720
rect 3445 21660 3455 21720
rect 3375 21610 3455 21660
rect 3375 21550 3385 21610
rect 3445 21550 3455 21610
rect 3375 21545 3455 21550
rect 3775 21720 3855 21725
rect 3775 21660 3785 21720
rect 3845 21660 3855 21720
rect 3775 21610 3855 21660
rect 3775 21550 3785 21610
rect 3845 21550 3855 21610
rect 3775 21545 3855 21550
rect 4175 21720 4255 21725
rect 4175 21660 4185 21720
rect 4245 21660 4255 21720
rect 4175 21610 4255 21660
rect 4175 21550 4185 21610
rect 4245 21550 4255 21610
rect 4175 21545 4255 21550
rect 4575 21720 4655 21725
rect 4575 21660 4585 21720
rect 4645 21660 4655 21720
rect 4575 21610 4655 21660
rect 4575 21550 4585 21610
rect 4645 21550 4655 21610
rect 4575 21545 4655 21550
rect 4975 21720 5055 21725
rect 4975 21660 4985 21720
rect 5045 21660 5055 21720
rect 4975 21610 5055 21660
rect 4975 21550 4985 21610
rect 5045 21550 5055 21610
rect 4975 21545 5055 21550
rect 5375 21720 5455 21725
rect 5375 21660 5385 21720
rect 5445 21660 5455 21720
rect 5375 21610 5455 21660
rect 5375 21550 5385 21610
rect 5445 21550 5455 21610
rect 5375 21545 5455 21550
rect 5775 21720 5855 21725
rect 5775 21660 5785 21720
rect 5845 21660 5855 21720
rect 5775 21610 5855 21660
rect 5775 21550 5785 21610
rect 5845 21550 5855 21610
rect 5775 21545 5855 21550
rect 6175 21720 6255 21725
rect 6175 21660 6185 21720
rect 6245 21660 6255 21720
rect 6175 21610 6255 21660
rect 6175 21550 6185 21610
rect 6245 21550 6255 21610
rect 6175 21545 6255 21550
rect 6575 21720 6655 21725
rect 6575 21660 6585 21720
rect 6645 21660 6655 21720
rect 6575 21610 6655 21660
rect 6575 21550 6585 21610
rect 6645 21550 6655 21610
rect 6575 21545 6655 21550
rect 6975 21720 7055 21725
rect 6975 21660 6985 21720
rect 7045 21660 7055 21720
rect 6975 21610 7055 21660
rect 6975 21550 6985 21610
rect 7045 21550 7055 21610
rect 6975 21545 7055 21550
rect 7375 21720 7455 21725
rect 7375 21660 7385 21720
rect 7445 21660 7455 21720
rect 7375 21610 7455 21660
rect 7375 21550 7385 21610
rect 7445 21550 7455 21610
rect 7375 21545 7455 21550
rect 7775 21720 7855 21725
rect 7775 21660 7785 21720
rect 7845 21660 7855 21720
rect 7775 21610 7855 21660
rect 7775 21550 7785 21610
rect 7845 21550 7855 21610
rect 7775 21545 7855 21550
rect 8175 21720 8255 21725
rect 8175 21660 8185 21720
rect 8245 21660 8255 21720
rect 8175 21610 8255 21660
rect 8175 21550 8185 21610
rect 8245 21550 8255 21610
rect 8175 21545 8255 21550
rect 8575 21720 8655 21725
rect 8575 21660 8585 21720
rect 8645 21660 8655 21720
rect 8575 21610 8655 21660
rect 8575 21550 8585 21610
rect 8645 21550 8655 21610
rect 8575 21545 8655 21550
rect 8975 21720 9055 21725
rect 8975 21660 8985 21720
rect 9045 21660 9055 21720
rect 8975 21610 9055 21660
rect 8975 21550 8985 21610
rect 9045 21550 9055 21610
rect 8975 21545 9055 21550
rect 9375 21720 9455 21725
rect 9375 21660 9385 21720
rect 9445 21660 9455 21720
rect 9375 21610 9455 21660
rect 9375 21550 9385 21610
rect 9445 21550 9455 21610
rect 9375 21545 9455 21550
rect 9775 21720 9855 21725
rect 9775 21660 9785 21720
rect 9845 21660 9855 21720
rect 9775 21610 9855 21660
rect 9775 21550 9785 21610
rect 9845 21550 9855 21610
rect 9775 21545 9855 21550
rect 10175 21720 10255 21725
rect 10175 21660 10185 21720
rect 10245 21660 10255 21720
rect 10175 21610 10255 21660
rect 10175 21550 10185 21610
rect 10245 21550 10255 21610
rect 10175 21545 10255 21550
rect 10575 21720 10655 21725
rect 10575 21660 10585 21720
rect 10645 21660 10655 21720
rect 10575 21610 10655 21660
rect 10575 21550 10585 21610
rect 10645 21550 10655 21610
rect 10575 21545 10655 21550
rect 10975 21720 11055 21725
rect 10975 21660 10985 21720
rect 11045 21660 11055 21720
rect 10975 21610 11055 21660
rect 10975 21550 10985 21610
rect 11045 21550 11055 21610
rect 10975 21545 11055 21550
rect 11375 21720 11455 21725
rect 11375 21660 11385 21720
rect 11445 21660 11455 21720
rect 11375 21610 11455 21660
rect 11375 21550 11385 21610
rect 11445 21550 11455 21610
rect 11375 21545 11455 21550
rect 11775 21720 11855 21725
rect 11775 21660 11785 21720
rect 11845 21660 11855 21720
rect 11775 21610 11855 21660
rect 11775 21550 11785 21610
rect 11845 21550 11855 21610
rect 11775 21545 11855 21550
rect 12175 21720 12255 21725
rect 12175 21660 12185 21720
rect 12245 21660 12255 21720
rect 12175 21610 12255 21660
rect 12175 21550 12185 21610
rect 12245 21550 12255 21610
rect 12175 21545 12255 21550
rect 12575 21720 12655 21725
rect 12575 21660 12585 21720
rect 12645 21660 12655 21720
rect 12575 21610 12655 21660
rect 12575 21550 12585 21610
rect 12645 21550 12655 21610
rect 12575 21545 12655 21550
rect 12975 21720 13055 21725
rect 12975 21660 12985 21720
rect 13045 21660 13055 21720
rect 12975 21610 13055 21660
rect 12975 21550 12985 21610
rect 13045 21550 13055 21610
rect 12975 21545 13055 21550
rect -215 21355 -155 21545
rect 185 21355 245 21545
rect 585 21355 645 21545
rect 985 21355 1045 21545
rect 1385 21355 1445 21545
rect 1785 21355 1845 21545
rect 2185 21355 2245 21545
rect 2585 21355 2645 21545
rect 2985 21355 3045 21545
rect 3385 21355 3445 21545
rect 3785 21355 3845 21545
rect 4185 21355 4245 21545
rect 4585 21355 4645 21545
rect 4985 21355 5045 21545
rect 5385 21355 5445 21545
rect 5785 21355 5845 21545
rect 6185 21355 6245 21545
rect 6585 21355 6645 21545
rect 6985 21355 7045 21545
rect 7385 21355 7445 21545
rect 7785 21355 7845 21545
rect 8185 21355 8245 21545
rect 8585 21355 8645 21545
rect 8985 21355 9045 21545
rect 9385 21355 9445 21545
rect 9785 21355 9845 21545
rect 10185 21355 10245 21545
rect 10585 21355 10645 21545
rect 10985 21355 11045 21545
rect 11385 21355 11445 21545
rect 11785 21355 11845 21545
rect 12185 21355 12245 21545
rect 12585 21355 12645 21545
rect 12985 21355 13045 21545
rect -225 21350 -145 21355
rect -225 21290 -215 21350
rect -155 21290 -145 21350
rect -225 21240 -145 21290
rect -225 21180 -215 21240
rect -155 21180 -145 21240
rect -225 21175 -145 21180
rect 175 21350 255 21355
rect 175 21290 185 21350
rect 245 21290 255 21350
rect 175 21240 255 21290
rect 175 21180 185 21240
rect 245 21180 255 21240
rect 175 21175 255 21180
rect 575 21350 655 21355
rect 575 21290 585 21350
rect 645 21290 655 21350
rect 575 21240 655 21290
rect 575 21180 585 21240
rect 645 21180 655 21240
rect 575 21175 655 21180
rect 975 21350 1055 21355
rect 975 21290 985 21350
rect 1045 21290 1055 21350
rect 975 21240 1055 21290
rect 975 21180 985 21240
rect 1045 21180 1055 21240
rect 975 21175 1055 21180
rect 1375 21350 1455 21355
rect 1375 21290 1385 21350
rect 1445 21290 1455 21350
rect 1375 21240 1455 21290
rect 1375 21180 1385 21240
rect 1445 21180 1455 21240
rect 1375 21175 1455 21180
rect 1775 21350 1855 21355
rect 1775 21290 1785 21350
rect 1845 21290 1855 21350
rect 1775 21240 1855 21290
rect 1775 21180 1785 21240
rect 1845 21180 1855 21240
rect 1775 21175 1855 21180
rect 2175 21350 2255 21355
rect 2175 21290 2185 21350
rect 2245 21290 2255 21350
rect 2175 21240 2255 21290
rect 2175 21180 2185 21240
rect 2245 21180 2255 21240
rect 2175 21175 2255 21180
rect 2575 21350 2655 21355
rect 2575 21290 2585 21350
rect 2645 21290 2655 21350
rect 2575 21240 2655 21290
rect 2575 21180 2585 21240
rect 2645 21180 2655 21240
rect 2575 21175 2655 21180
rect 2975 21350 3055 21355
rect 2975 21290 2985 21350
rect 3045 21290 3055 21350
rect 2975 21240 3055 21290
rect 2975 21180 2985 21240
rect 3045 21180 3055 21240
rect 2975 21175 3055 21180
rect 3375 21350 3455 21355
rect 3375 21290 3385 21350
rect 3445 21290 3455 21350
rect 3375 21240 3455 21290
rect 3375 21180 3385 21240
rect 3445 21180 3455 21240
rect 3375 21175 3455 21180
rect 3775 21350 3855 21355
rect 3775 21290 3785 21350
rect 3845 21290 3855 21350
rect 3775 21240 3855 21290
rect 3775 21180 3785 21240
rect 3845 21180 3855 21240
rect 3775 21175 3855 21180
rect 4175 21350 4255 21355
rect 4175 21290 4185 21350
rect 4245 21290 4255 21350
rect 4175 21240 4255 21290
rect 4175 21180 4185 21240
rect 4245 21180 4255 21240
rect 4175 21175 4255 21180
rect 4575 21350 4655 21355
rect 4575 21290 4585 21350
rect 4645 21290 4655 21350
rect 4575 21240 4655 21290
rect 4575 21180 4585 21240
rect 4645 21180 4655 21240
rect 4575 21175 4655 21180
rect 4975 21350 5055 21355
rect 4975 21290 4985 21350
rect 5045 21290 5055 21350
rect 4975 21240 5055 21290
rect 4975 21180 4985 21240
rect 5045 21180 5055 21240
rect 4975 21175 5055 21180
rect 5375 21350 5455 21355
rect 5375 21290 5385 21350
rect 5445 21290 5455 21350
rect 5375 21240 5455 21290
rect 5375 21180 5385 21240
rect 5445 21180 5455 21240
rect 5375 21175 5455 21180
rect 5775 21350 5855 21355
rect 5775 21290 5785 21350
rect 5845 21290 5855 21350
rect 5775 21240 5855 21290
rect 5775 21180 5785 21240
rect 5845 21180 5855 21240
rect 5775 21175 5855 21180
rect 6175 21350 6255 21355
rect 6175 21290 6185 21350
rect 6245 21290 6255 21350
rect 6175 21240 6255 21290
rect 6175 21180 6185 21240
rect 6245 21180 6255 21240
rect 6175 21175 6255 21180
rect 6575 21350 6655 21355
rect 6575 21290 6585 21350
rect 6645 21290 6655 21350
rect 6575 21240 6655 21290
rect 6575 21180 6585 21240
rect 6645 21180 6655 21240
rect 6575 21175 6655 21180
rect 6975 21350 7055 21355
rect 6975 21290 6985 21350
rect 7045 21290 7055 21350
rect 6975 21240 7055 21290
rect 6975 21180 6985 21240
rect 7045 21180 7055 21240
rect 6975 21175 7055 21180
rect 7375 21350 7455 21355
rect 7375 21290 7385 21350
rect 7445 21290 7455 21350
rect 7375 21240 7455 21290
rect 7375 21180 7385 21240
rect 7445 21180 7455 21240
rect 7375 21175 7455 21180
rect 7775 21350 7855 21355
rect 7775 21290 7785 21350
rect 7845 21290 7855 21350
rect 7775 21240 7855 21290
rect 7775 21180 7785 21240
rect 7845 21180 7855 21240
rect 7775 21175 7855 21180
rect 8175 21350 8255 21355
rect 8175 21290 8185 21350
rect 8245 21290 8255 21350
rect 8175 21240 8255 21290
rect 8175 21180 8185 21240
rect 8245 21180 8255 21240
rect 8175 21175 8255 21180
rect 8575 21350 8655 21355
rect 8575 21290 8585 21350
rect 8645 21290 8655 21350
rect 8575 21240 8655 21290
rect 8575 21180 8585 21240
rect 8645 21180 8655 21240
rect 8575 21175 8655 21180
rect 8975 21350 9055 21355
rect 8975 21290 8985 21350
rect 9045 21290 9055 21350
rect 8975 21240 9055 21290
rect 8975 21180 8985 21240
rect 9045 21180 9055 21240
rect 8975 21175 9055 21180
rect 9375 21350 9455 21355
rect 9375 21290 9385 21350
rect 9445 21290 9455 21350
rect 9375 21240 9455 21290
rect 9375 21180 9385 21240
rect 9445 21180 9455 21240
rect 9375 21175 9455 21180
rect 9775 21350 9855 21355
rect 9775 21290 9785 21350
rect 9845 21290 9855 21350
rect 9775 21240 9855 21290
rect 9775 21180 9785 21240
rect 9845 21180 9855 21240
rect 9775 21175 9855 21180
rect 10175 21350 10255 21355
rect 10175 21290 10185 21350
rect 10245 21290 10255 21350
rect 10175 21240 10255 21290
rect 10175 21180 10185 21240
rect 10245 21180 10255 21240
rect 10175 21175 10255 21180
rect 10575 21350 10655 21355
rect 10575 21290 10585 21350
rect 10645 21290 10655 21350
rect 10575 21240 10655 21290
rect 10575 21180 10585 21240
rect 10645 21180 10655 21240
rect 10575 21175 10655 21180
rect 10975 21350 11055 21355
rect 10975 21290 10985 21350
rect 11045 21290 11055 21350
rect 10975 21240 11055 21290
rect 10975 21180 10985 21240
rect 11045 21180 11055 21240
rect 10975 21175 11055 21180
rect 11375 21350 11455 21355
rect 11375 21290 11385 21350
rect 11445 21290 11455 21350
rect 11375 21240 11455 21290
rect 11375 21180 11385 21240
rect 11445 21180 11455 21240
rect 11375 21175 11455 21180
rect 11775 21350 11855 21355
rect 11775 21290 11785 21350
rect 11845 21290 11855 21350
rect 11775 21240 11855 21290
rect 11775 21180 11785 21240
rect 11845 21180 11855 21240
rect 11775 21175 11855 21180
rect 12175 21350 12255 21355
rect 12175 21290 12185 21350
rect 12245 21290 12255 21350
rect 12175 21240 12255 21290
rect 12175 21180 12185 21240
rect 12245 21180 12255 21240
rect 12175 21175 12255 21180
rect 12575 21350 12655 21355
rect 12575 21290 12585 21350
rect 12645 21290 12655 21350
rect 12575 21240 12655 21290
rect 12575 21180 12585 21240
rect 12645 21180 12655 21240
rect 12575 21175 12655 21180
rect 12975 21350 13055 21355
rect 12975 21290 12985 21350
rect 13045 21290 13055 21350
rect 12975 21240 13055 21290
rect 12975 21180 12985 21240
rect 13045 21180 13055 21240
rect 12975 21175 13055 21180
rect -215 20985 -155 21175
rect 185 20985 245 21175
rect 585 20985 645 21175
rect 985 20985 1045 21175
rect 1385 20985 1445 21175
rect 1785 20985 1845 21175
rect 2185 20985 2245 21175
rect 2585 20985 2645 21175
rect 2985 20985 3045 21175
rect 3385 20985 3445 21175
rect 3785 20985 3845 21175
rect 4185 20985 4245 21175
rect 4585 20985 4645 21175
rect 4985 20985 5045 21175
rect 5385 20985 5445 21175
rect 5785 20985 5845 21175
rect 6185 20985 6245 21175
rect 6585 20985 6645 21175
rect 6985 20985 7045 21175
rect 7385 20985 7445 21175
rect 7785 20985 7845 21175
rect 8185 20985 8245 21175
rect 8585 20985 8645 21175
rect 8985 20985 9045 21175
rect 9385 20985 9445 21175
rect 9785 20985 9845 21175
rect 10185 20985 10245 21175
rect 10585 20985 10645 21175
rect 10985 20985 11045 21175
rect 11385 20985 11445 21175
rect 11785 20985 11845 21175
rect 12185 20985 12245 21175
rect 12585 20985 12645 21175
rect 12985 20985 13045 21175
rect -225 20980 -145 20985
rect -225 20920 -215 20980
rect -155 20920 -145 20980
rect -225 20870 -145 20920
rect -225 20810 -215 20870
rect -155 20810 -145 20870
rect -225 20805 -145 20810
rect 175 20980 255 20985
rect 175 20920 185 20980
rect 245 20920 255 20980
rect 175 20870 255 20920
rect 175 20810 185 20870
rect 245 20810 255 20870
rect 175 20805 255 20810
rect 575 20980 655 20985
rect 575 20920 585 20980
rect 645 20920 655 20980
rect 575 20870 655 20920
rect 575 20810 585 20870
rect 645 20810 655 20870
rect 575 20805 655 20810
rect 975 20980 1055 20985
rect 975 20920 985 20980
rect 1045 20920 1055 20980
rect 975 20870 1055 20920
rect 975 20810 985 20870
rect 1045 20810 1055 20870
rect 975 20805 1055 20810
rect 1375 20980 1455 20985
rect 1375 20920 1385 20980
rect 1445 20920 1455 20980
rect 1375 20870 1455 20920
rect 1375 20810 1385 20870
rect 1445 20810 1455 20870
rect 1375 20805 1455 20810
rect 1775 20980 1855 20985
rect 1775 20920 1785 20980
rect 1845 20920 1855 20980
rect 1775 20870 1855 20920
rect 1775 20810 1785 20870
rect 1845 20810 1855 20870
rect 1775 20805 1855 20810
rect 2175 20980 2255 20985
rect 2175 20920 2185 20980
rect 2245 20920 2255 20980
rect 2175 20870 2255 20920
rect 2175 20810 2185 20870
rect 2245 20810 2255 20870
rect 2175 20805 2255 20810
rect 2575 20980 2655 20985
rect 2575 20920 2585 20980
rect 2645 20920 2655 20980
rect 2575 20870 2655 20920
rect 2575 20810 2585 20870
rect 2645 20810 2655 20870
rect 2575 20805 2655 20810
rect 2975 20980 3055 20985
rect 2975 20920 2985 20980
rect 3045 20920 3055 20980
rect 2975 20870 3055 20920
rect 2975 20810 2985 20870
rect 3045 20810 3055 20870
rect 2975 20805 3055 20810
rect 3375 20980 3455 20985
rect 3375 20920 3385 20980
rect 3445 20920 3455 20980
rect 3375 20870 3455 20920
rect 3375 20810 3385 20870
rect 3445 20810 3455 20870
rect 3375 20805 3455 20810
rect 3775 20980 3855 20985
rect 3775 20920 3785 20980
rect 3845 20920 3855 20980
rect 3775 20870 3855 20920
rect 3775 20810 3785 20870
rect 3845 20810 3855 20870
rect 3775 20805 3855 20810
rect 4175 20980 4255 20985
rect 4175 20920 4185 20980
rect 4245 20920 4255 20980
rect 4175 20870 4255 20920
rect 4175 20810 4185 20870
rect 4245 20810 4255 20870
rect 4175 20805 4255 20810
rect 4575 20980 4655 20985
rect 4575 20920 4585 20980
rect 4645 20920 4655 20980
rect 4575 20870 4655 20920
rect 4575 20810 4585 20870
rect 4645 20810 4655 20870
rect 4575 20805 4655 20810
rect 4975 20980 5055 20985
rect 4975 20920 4985 20980
rect 5045 20920 5055 20980
rect 4975 20870 5055 20920
rect 4975 20810 4985 20870
rect 5045 20810 5055 20870
rect 4975 20805 5055 20810
rect 5375 20980 5455 20985
rect 5375 20920 5385 20980
rect 5445 20920 5455 20980
rect 5375 20870 5455 20920
rect 5375 20810 5385 20870
rect 5445 20810 5455 20870
rect 5375 20805 5455 20810
rect 5775 20980 5855 20985
rect 5775 20920 5785 20980
rect 5845 20920 5855 20980
rect 5775 20870 5855 20920
rect 5775 20810 5785 20870
rect 5845 20810 5855 20870
rect 5775 20805 5855 20810
rect 6175 20980 6255 20985
rect 6175 20920 6185 20980
rect 6245 20920 6255 20980
rect 6175 20870 6255 20920
rect 6175 20810 6185 20870
rect 6245 20810 6255 20870
rect 6175 20805 6255 20810
rect 6575 20980 6655 20985
rect 6575 20920 6585 20980
rect 6645 20920 6655 20980
rect 6575 20870 6655 20920
rect 6575 20810 6585 20870
rect 6645 20810 6655 20870
rect 6575 20805 6655 20810
rect 6975 20980 7055 20985
rect 6975 20920 6985 20980
rect 7045 20920 7055 20980
rect 6975 20870 7055 20920
rect 6975 20810 6985 20870
rect 7045 20810 7055 20870
rect 6975 20805 7055 20810
rect 7375 20980 7455 20985
rect 7375 20920 7385 20980
rect 7445 20920 7455 20980
rect 7375 20870 7455 20920
rect 7375 20810 7385 20870
rect 7445 20810 7455 20870
rect 7375 20805 7455 20810
rect 7775 20980 7855 20985
rect 7775 20920 7785 20980
rect 7845 20920 7855 20980
rect 7775 20870 7855 20920
rect 7775 20810 7785 20870
rect 7845 20810 7855 20870
rect 7775 20805 7855 20810
rect 8175 20980 8255 20985
rect 8175 20920 8185 20980
rect 8245 20920 8255 20980
rect 8175 20870 8255 20920
rect 8175 20810 8185 20870
rect 8245 20810 8255 20870
rect 8175 20805 8255 20810
rect 8575 20980 8655 20985
rect 8575 20920 8585 20980
rect 8645 20920 8655 20980
rect 8575 20870 8655 20920
rect 8575 20810 8585 20870
rect 8645 20810 8655 20870
rect 8575 20805 8655 20810
rect 8975 20980 9055 20985
rect 8975 20920 8985 20980
rect 9045 20920 9055 20980
rect 8975 20870 9055 20920
rect 8975 20810 8985 20870
rect 9045 20810 9055 20870
rect 8975 20805 9055 20810
rect 9375 20980 9455 20985
rect 9375 20920 9385 20980
rect 9445 20920 9455 20980
rect 9375 20870 9455 20920
rect 9375 20810 9385 20870
rect 9445 20810 9455 20870
rect 9375 20805 9455 20810
rect 9775 20980 9855 20985
rect 9775 20920 9785 20980
rect 9845 20920 9855 20980
rect 9775 20870 9855 20920
rect 9775 20810 9785 20870
rect 9845 20810 9855 20870
rect 9775 20805 9855 20810
rect 10175 20980 10255 20985
rect 10175 20920 10185 20980
rect 10245 20920 10255 20980
rect 10175 20870 10255 20920
rect 10175 20810 10185 20870
rect 10245 20810 10255 20870
rect 10175 20805 10255 20810
rect 10575 20980 10655 20985
rect 10575 20920 10585 20980
rect 10645 20920 10655 20980
rect 10575 20870 10655 20920
rect 10575 20810 10585 20870
rect 10645 20810 10655 20870
rect 10575 20805 10655 20810
rect 10975 20980 11055 20985
rect 10975 20920 10985 20980
rect 11045 20920 11055 20980
rect 10975 20870 11055 20920
rect 10975 20810 10985 20870
rect 11045 20810 11055 20870
rect 10975 20805 11055 20810
rect 11375 20980 11455 20985
rect 11375 20920 11385 20980
rect 11445 20920 11455 20980
rect 11375 20870 11455 20920
rect 11375 20810 11385 20870
rect 11445 20810 11455 20870
rect 11375 20805 11455 20810
rect 11775 20980 11855 20985
rect 11775 20920 11785 20980
rect 11845 20920 11855 20980
rect 11775 20870 11855 20920
rect 11775 20810 11785 20870
rect 11845 20810 11855 20870
rect 11775 20805 11855 20810
rect 12175 20980 12255 20985
rect 12175 20920 12185 20980
rect 12245 20920 12255 20980
rect 12175 20870 12255 20920
rect 12175 20810 12185 20870
rect 12245 20810 12255 20870
rect 12175 20805 12255 20810
rect 12575 20980 12655 20985
rect 12575 20920 12585 20980
rect 12645 20920 12655 20980
rect 12575 20870 12655 20920
rect 12575 20810 12585 20870
rect 12645 20810 12655 20870
rect 12575 20805 12655 20810
rect 12975 20980 13055 20985
rect 12975 20920 12985 20980
rect 13045 20920 13055 20980
rect 12975 20870 13055 20920
rect 12975 20810 12985 20870
rect 13045 20810 13055 20870
rect 12975 20805 13055 20810
rect -215 20615 -155 20805
rect 185 20615 245 20805
rect 585 20615 645 20805
rect 985 20615 1045 20805
rect 1385 20615 1445 20805
rect 1785 20615 1845 20805
rect 2185 20615 2245 20805
rect 2585 20615 2645 20805
rect 2985 20615 3045 20805
rect 3385 20615 3445 20805
rect 3785 20615 3845 20805
rect 4185 20615 4245 20805
rect 4585 20615 4645 20805
rect 4985 20615 5045 20805
rect 5385 20615 5445 20805
rect 5785 20615 5845 20805
rect 6185 20615 6245 20805
rect 6585 20615 6645 20805
rect 6985 20615 7045 20805
rect 7385 20615 7445 20805
rect 7785 20615 7845 20805
rect 8185 20615 8245 20805
rect 8585 20615 8645 20805
rect 8985 20615 9045 20805
rect 9385 20615 9445 20805
rect 9785 20615 9845 20805
rect 10185 20615 10245 20805
rect 10585 20615 10645 20805
rect 10985 20615 11045 20805
rect 11385 20615 11445 20805
rect 11785 20615 11845 20805
rect 12185 20615 12245 20805
rect 12585 20615 12645 20805
rect 12985 20615 13045 20805
rect -225 20610 -145 20615
rect -225 20550 -215 20610
rect -155 20550 -145 20610
rect -225 20500 -145 20550
rect -225 20440 -215 20500
rect -155 20440 -145 20500
rect -225 20435 -145 20440
rect 175 20610 255 20615
rect 175 20550 185 20610
rect 245 20550 255 20610
rect 175 20500 255 20550
rect 175 20440 185 20500
rect 245 20440 255 20500
rect 175 20435 255 20440
rect 575 20610 655 20615
rect 575 20550 585 20610
rect 645 20550 655 20610
rect 575 20500 655 20550
rect 575 20440 585 20500
rect 645 20440 655 20500
rect 575 20435 655 20440
rect 975 20610 1055 20615
rect 975 20550 985 20610
rect 1045 20550 1055 20610
rect 975 20500 1055 20550
rect 975 20440 985 20500
rect 1045 20440 1055 20500
rect 975 20435 1055 20440
rect 1375 20610 1455 20615
rect 1375 20550 1385 20610
rect 1445 20550 1455 20610
rect 1375 20500 1455 20550
rect 1375 20440 1385 20500
rect 1445 20440 1455 20500
rect 1375 20435 1455 20440
rect 1775 20610 1855 20615
rect 1775 20550 1785 20610
rect 1845 20550 1855 20610
rect 1775 20500 1855 20550
rect 1775 20440 1785 20500
rect 1845 20440 1855 20500
rect 1775 20435 1855 20440
rect 2175 20610 2255 20615
rect 2175 20550 2185 20610
rect 2245 20550 2255 20610
rect 2175 20500 2255 20550
rect 2175 20440 2185 20500
rect 2245 20440 2255 20500
rect 2175 20435 2255 20440
rect 2575 20610 2655 20615
rect 2575 20550 2585 20610
rect 2645 20550 2655 20610
rect 2575 20500 2655 20550
rect 2575 20440 2585 20500
rect 2645 20440 2655 20500
rect 2575 20435 2655 20440
rect 2975 20610 3055 20615
rect 2975 20550 2985 20610
rect 3045 20550 3055 20610
rect 2975 20500 3055 20550
rect 2975 20440 2985 20500
rect 3045 20440 3055 20500
rect 2975 20435 3055 20440
rect 3375 20610 3455 20615
rect 3375 20550 3385 20610
rect 3445 20550 3455 20610
rect 3375 20500 3455 20550
rect 3375 20440 3385 20500
rect 3445 20440 3455 20500
rect 3375 20435 3455 20440
rect 3775 20610 3855 20615
rect 3775 20550 3785 20610
rect 3845 20550 3855 20610
rect 3775 20500 3855 20550
rect 3775 20440 3785 20500
rect 3845 20440 3855 20500
rect 3775 20435 3855 20440
rect 4175 20610 4255 20615
rect 4175 20550 4185 20610
rect 4245 20550 4255 20610
rect 4175 20500 4255 20550
rect 4175 20440 4185 20500
rect 4245 20440 4255 20500
rect 4175 20435 4255 20440
rect 4575 20610 4655 20615
rect 4575 20550 4585 20610
rect 4645 20550 4655 20610
rect 4575 20500 4655 20550
rect 4575 20440 4585 20500
rect 4645 20440 4655 20500
rect 4575 20435 4655 20440
rect 4975 20610 5055 20615
rect 4975 20550 4985 20610
rect 5045 20550 5055 20610
rect 4975 20500 5055 20550
rect 4975 20440 4985 20500
rect 5045 20440 5055 20500
rect 4975 20435 5055 20440
rect 5375 20610 5455 20615
rect 5375 20550 5385 20610
rect 5445 20550 5455 20610
rect 5375 20500 5455 20550
rect 5375 20440 5385 20500
rect 5445 20440 5455 20500
rect 5375 20435 5455 20440
rect 5775 20610 5855 20615
rect 5775 20550 5785 20610
rect 5845 20550 5855 20610
rect 5775 20500 5855 20550
rect 5775 20440 5785 20500
rect 5845 20440 5855 20500
rect 5775 20435 5855 20440
rect 6175 20610 6255 20615
rect 6175 20550 6185 20610
rect 6245 20550 6255 20610
rect 6175 20500 6255 20550
rect 6175 20440 6185 20500
rect 6245 20440 6255 20500
rect 6175 20435 6255 20440
rect 6575 20610 6655 20615
rect 6575 20550 6585 20610
rect 6645 20550 6655 20610
rect 6575 20500 6655 20550
rect 6575 20440 6585 20500
rect 6645 20440 6655 20500
rect 6575 20435 6655 20440
rect 6975 20610 7055 20615
rect 6975 20550 6985 20610
rect 7045 20550 7055 20610
rect 6975 20500 7055 20550
rect 6975 20440 6985 20500
rect 7045 20440 7055 20500
rect 6975 20435 7055 20440
rect 7375 20610 7455 20615
rect 7375 20550 7385 20610
rect 7445 20550 7455 20610
rect 7375 20500 7455 20550
rect 7375 20440 7385 20500
rect 7445 20440 7455 20500
rect 7375 20435 7455 20440
rect 7775 20610 7855 20615
rect 7775 20550 7785 20610
rect 7845 20550 7855 20610
rect 7775 20500 7855 20550
rect 7775 20440 7785 20500
rect 7845 20440 7855 20500
rect 7775 20435 7855 20440
rect 8175 20610 8255 20615
rect 8175 20550 8185 20610
rect 8245 20550 8255 20610
rect 8175 20500 8255 20550
rect 8175 20440 8185 20500
rect 8245 20440 8255 20500
rect 8175 20435 8255 20440
rect 8575 20610 8655 20615
rect 8575 20550 8585 20610
rect 8645 20550 8655 20610
rect 8575 20500 8655 20550
rect 8575 20440 8585 20500
rect 8645 20440 8655 20500
rect 8575 20435 8655 20440
rect 8975 20610 9055 20615
rect 8975 20550 8985 20610
rect 9045 20550 9055 20610
rect 8975 20500 9055 20550
rect 8975 20440 8985 20500
rect 9045 20440 9055 20500
rect 8975 20435 9055 20440
rect 9375 20610 9455 20615
rect 9375 20550 9385 20610
rect 9445 20550 9455 20610
rect 9375 20500 9455 20550
rect 9375 20440 9385 20500
rect 9445 20440 9455 20500
rect 9375 20435 9455 20440
rect 9775 20610 9855 20615
rect 9775 20550 9785 20610
rect 9845 20550 9855 20610
rect 9775 20500 9855 20550
rect 9775 20440 9785 20500
rect 9845 20440 9855 20500
rect 9775 20435 9855 20440
rect 10175 20610 10255 20615
rect 10175 20550 10185 20610
rect 10245 20550 10255 20610
rect 10175 20500 10255 20550
rect 10175 20440 10185 20500
rect 10245 20440 10255 20500
rect 10175 20435 10255 20440
rect 10575 20610 10655 20615
rect 10575 20550 10585 20610
rect 10645 20550 10655 20610
rect 10575 20500 10655 20550
rect 10575 20440 10585 20500
rect 10645 20440 10655 20500
rect 10575 20435 10655 20440
rect 10975 20610 11055 20615
rect 10975 20550 10985 20610
rect 11045 20550 11055 20610
rect 10975 20500 11055 20550
rect 10975 20440 10985 20500
rect 11045 20440 11055 20500
rect 10975 20435 11055 20440
rect 11375 20610 11455 20615
rect 11375 20550 11385 20610
rect 11445 20550 11455 20610
rect 11375 20500 11455 20550
rect 11375 20440 11385 20500
rect 11445 20440 11455 20500
rect 11375 20435 11455 20440
rect 11775 20610 11855 20615
rect 11775 20550 11785 20610
rect 11845 20550 11855 20610
rect 11775 20500 11855 20550
rect 11775 20440 11785 20500
rect 11845 20440 11855 20500
rect 11775 20435 11855 20440
rect 12175 20610 12255 20615
rect 12175 20550 12185 20610
rect 12245 20550 12255 20610
rect 12175 20500 12255 20550
rect 12175 20440 12185 20500
rect 12245 20440 12255 20500
rect 12175 20435 12255 20440
rect 12575 20610 12655 20615
rect 12575 20550 12585 20610
rect 12645 20550 12655 20610
rect 12575 20500 12655 20550
rect 12575 20440 12585 20500
rect 12645 20440 12655 20500
rect 12575 20435 12655 20440
rect 12975 20610 13055 20615
rect 12975 20550 12985 20610
rect 13045 20550 13055 20610
rect 12975 20500 13055 20550
rect 12975 20440 12985 20500
rect 13045 20440 13055 20500
rect 12975 20435 13055 20440
rect -215 20245 -155 20435
rect 185 20245 245 20435
rect 585 20245 645 20435
rect 985 20245 1045 20435
rect 1385 20245 1445 20435
rect 1785 20245 1845 20435
rect 2185 20245 2245 20435
rect 2585 20245 2645 20435
rect 2985 20245 3045 20435
rect 3385 20245 3445 20435
rect 3785 20245 3845 20435
rect 4185 20245 4245 20435
rect 4585 20245 4645 20435
rect 4985 20245 5045 20435
rect 5385 20245 5445 20435
rect 5785 20245 5845 20435
rect 6185 20245 6245 20435
rect 6585 20245 6645 20435
rect 6985 20245 7045 20435
rect 7385 20245 7445 20435
rect 7785 20245 7845 20435
rect 8185 20245 8245 20435
rect 8585 20245 8645 20435
rect 8985 20245 9045 20435
rect 9385 20245 9445 20435
rect 9785 20245 9845 20435
rect 10185 20245 10245 20435
rect 10585 20245 10645 20435
rect 10985 20245 11045 20435
rect 11385 20245 11445 20435
rect 11785 20245 11845 20435
rect 12185 20245 12245 20435
rect 12585 20245 12645 20435
rect 12985 20245 13045 20435
rect -225 20240 -145 20245
rect -225 20180 -215 20240
rect -155 20180 -145 20240
rect -225 20130 -145 20180
rect -225 20070 -215 20130
rect -155 20070 -145 20130
rect -225 20065 -145 20070
rect 175 20240 255 20245
rect 175 20180 185 20240
rect 245 20180 255 20240
rect 175 20130 255 20180
rect 175 20070 185 20130
rect 245 20070 255 20130
rect 175 20065 255 20070
rect 575 20240 655 20245
rect 575 20180 585 20240
rect 645 20180 655 20240
rect 575 20130 655 20180
rect 575 20070 585 20130
rect 645 20070 655 20130
rect 575 20065 655 20070
rect 975 20240 1055 20245
rect 975 20180 985 20240
rect 1045 20180 1055 20240
rect 975 20130 1055 20180
rect 975 20070 985 20130
rect 1045 20070 1055 20130
rect 975 20065 1055 20070
rect 1375 20240 1455 20245
rect 1375 20180 1385 20240
rect 1445 20180 1455 20240
rect 1375 20130 1455 20180
rect 1375 20070 1385 20130
rect 1445 20070 1455 20130
rect 1375 20065 1455 20070
rect 1775 20240 1855 20245
rect 1775 20180 1785 20240
rect 1845 20180 1855 20240
rect 1775 20130 1855 20180
rect 1775 20070 1785 20130
rect 1845 20070 1855 20130
rect 1775 20065 1855 20070
rect 2175 20240 2255 20245
rect 2175 20180 2185 20240
rect 2245 20180 2255 20240
rect 2175 20130 2255 20180
rect 2175 20070 2185 20130
rect 2245 20070 2255 20130
rect 2175 20065 2255 20070
rect 2575 20240 2655 20245
rect 2575 20180 2585 20240
rect 2645 20180 2655 20240
rect 2575 20130 2655 20180
rect 2575 20070 2585 20130
rect 2645 20070 2655 20130
rect 2575 20065 2655 20070
rect 2975 20240 3055 20245
rect 2975 20180 2985 20240
rect 3045 20180 3055 20240
rect 2975 20130 3055 20180
rect 2975 20070 2985 20130
rect 3045 20070 3055 20130
rect 2975 20065 3055 20070
rect 3375 20240 3455 20245
rect 3375 20180 3385 20240
rect 3445 20180 3455 20240
rect 3375 20130 3455 20180
rect 3375 20070 3385 20130
rect 3445 20070 3455 20130
rect 3375 20065 3455 20070
rect 3775 20240 3855 20245
rect 3775 20180 3785 20240
rect 3845 20180 3855 20240
rect 3775 20130 3855 20180
rect 3775 20070 3785 20130
rect 3845 20070 3855 20130
rect 3775 20065 3855 20070
rect 4175 20240 4255 20245
rect 4175 20180 4185 20240
rect 4245 20180 4255 20240
rect 4175 20130 4255 20180
rect 4175 20070 4185 20130
rect 4245 20070 4255 20130
rect 4175 20065 4255 20070
rect 4575 20240 4655 20245
rect 4575 20180 4585 20240
rect 4645 20180 4655 20240
rect 4575 20130 4655 20180
rect 4575 20070 4585 20130
rect 4645 20070 4655 20130
rect 4575 20065 4655 20070
rect 4975 20240 5055 20245
rect 4975 20180 4985 20240
rect 5045 20180 5055 20240
rect 4975 20130 5055 20180
rect 4975 20070 4985 20130
rect 5045 20070 5055 20130
rect 4975 20065 5055 20070
rect 5375 20240 5455 20245
rect 5375 20180 5385 20240
rect 5445 20180 5455 20240
rect 5375 20130 5455 20180
rect 5375 20070 5385 20130
rect 5445 20070 5455 20130
rect 5375 20065 5455 20070
rect 5775 20240 5855 20245
rect 5775 20180 5785 20240
rect 5845 20180 5855 20240
rect 5775 20130 5855 20180
rect 5775 20070 5785 20130
rect 5845 20070 5855 20130
rect 5775 20065 5855 20070
rect 6175 20240 6255 20245
rect 6175 20180 6185 20240
rect 6245 20180 6255 20240
rect 6175 20130 6255 20180
rect 6175 20070 6185 20130
rect 6245 20070 6255 20130
rect 6175 20065 6255 20070
rect 6575 20240 6655 20245
rect 6575 20180 6585 20240
rect 6645 20180 6655 20240
rect 6575 20130 6655 20180
rect 6575 20070 6585 20130
rect 6645 20070 6655 20130
rect 6575 20065 6655 20070
rect 6975 20240 7055 20245
rect 6975 20180 6985 20240
rect 7045 20180 7055 20240
rect 6975 20130 7055 20180
rect 6975 20070 6985 20130
rect 7045 20070 7055 20130
rect 6975 20065 7055 20070
rect 7375 20240 7455 20245
rect 7375 20180 7385 20240
rect 7445 20180 7455 20240
rect 7375 20130 7455 20180
rect 7375 20070 7385 20130
rect 7445 20070 7455 20130
rect 7375 20065 7455 20070
rect 7775 20240 7855 20245
rect 7775 20180 7785 20240
rect 7845 20180 7855 20240
rect 7775 20130 7855 20180
rect 7775 20070 7785 20130
rect 7845 20070 7855 20130
rect 7775 20065 7855 20070
rect 8175 20240 8255 20245
rect 8175 20180 8185 20240
rect 8245 20180 8255 20240
rect 8175 20130 8255 20180
rect 8175 20070 8185 20130
rect 8245 20070 8255 20130
rect 8175 20065 8255 20070
rect 8575 20240 8655 20245
rect 8575 20180 8585 20240
rect 8645 20180 8655 20240
rect 8575 20130 8655 20180
rect 8575 20070 8585 20130
rect 8645 20070 8655 20130
rect 8575 20065 8655 20070
rect 8975 20240 9055 20245
rect 8975 20180 8985 20240
rect 9045 20180 9055 20240
rect 8975 20130 9055 20180
rect 8975 20070 8985 20130
rect 9045 20070 9055 20130
rect 8975 20065 9055 20070
rect 9375 20240 9455 20245
rect 9375 20180 9385 20240
rect 9445 20180 9455 20240
rect 9375 20130 9455 20180
rect 9375 20070 9385 20130
rect 9445 20070 9455 20130
rect 9375 20065 9455 20070
rect 9775 20240 9855 20245
rect 9775 20180 9785 20240
rect 9845 20180 9855 20240
rect 9775 20130 9855 20180
rect 9775 20070 9785 20130
rect 9845 20070 9855 20130
rect 9775 20065 9855 20070
rect 10175 20240 10255 20245
rect 10175 20180 10185 20240
rect 10245 20180 10255 20240
rect 10175 20130 10255 20180
rect 10175 20070 10185 20130
rect 10245 20070 10255 20130
rect 10175 20065 10255 20070
rect 10575 20240 10655 20245
rect 10575 20180 10585 20240
rect 10645 20180 10655 20240
rect 10575 20130 10655 20180
rect 10575 20070 10585 20130
rect 10645 20070 10655 20130
rect 10575 20065 10655 20070
rect 10975 20240 11055 20245
rect 10975 20180 10985 20240
rect 11045 20180 11055 20240
rect 10975 20130 11055 20180
rect 10975 20070 10985 20130
rect 11045 20070 11055 20130
rect 10975 20065 11055 20070
rect 11375 20240 11455 20245
rect 11375 20180 11385 20240
rect 11445 20180 11455 20240
rect 11375 20130 11455 20180
rect 11375 20070 11385 20130
rect 11445 20070 11455 20130
rect 11375 20065 11455 20070
rect 11775 20240 11855 20245
rect 11775 20180 11785 20240
rect 11845 20180 11855 20240
rect 11775 20130 11855 20180
rect 11775 20070 11785 20130
rect 11845 20070 11855 20130
rect 11775 20065 11855 20070
rect 12175 20240 12255 20245
rect 12175 20180 12185 20240
rect 12245 20180 12255 20240
rect 12175 20130 12255 20180
rect 12175 20070 12185 20130
rect 12245 20070 12255 20130
rect 12175 20065 12255 20070
rect 12575 20240 12655 20245
rect 12575 20180 12585 20240
rect 12645 20180 12655 20240
rect 12575 20130 12655 20180
rect 12575 20070 12585 20130
rect 12645 20070 12655 20130
rect 12575 20065 12655 20070
rect 12975 20240 13055 20245
rect 12975 20180 12985 20240
rect 13045 20180 13055 20240
rect 12975 20130 13055 20180
rect 12975 20070 12985 20130
rect 13045 20070 13055 20130
rect 12975 20065 13055 20070
rect -215 19875 -155 20065
rect 185 19875 245 20065
rect 585 19875 645 20065
rect 985 19875 1045 20065
rect 1385 19875 1445 20065
rect 1785 19875 1845 20065
rect 2185 19875 2245 20065
rect 2585 19875 2645 20065
rect 2985 19875 3045 20065
rect 3385 19875 3445 20065
rect 3785 19875 3845 20065
rect 4185 19875 4245 20065
rect 4585 19875 4645 20065
rect 4985 19875 5045 20065
rect 5385 19875 5445 20065
rect 5785 19875 5845 20065
rect 6185 19875 6245 20065
rect 6585 19875 6645 20065
rect 6985 19875 7045 20065
rect 7385 19875 7445 20065
rect 7785 19875 7845 20065
rect 8185 19875 8245 20065
rect 8585 19875 8645 20065
rect 8985 19875 9045 20065
rect 9385 19875 9445 20065
rect 9785 19875 9845 20065
rect 10185 19875 10245 20065
rect 10585 19875 10645 20065
rect 10985 19875 11045 20065
rect 11385 19875 11445 20065
rect 11785 19875 11845 20065
rect 12185 19875 12245 20065
rect 12585 19875 12645 20065
rect 12985 19875 13045 20065
rect -225 19870 -145 19875
rect -225 19810 -215 19870
rect -155 19810 -145 19870
rect -225 19760 -145 19810
rect -225 19700 -215 19760
rect -155 19700 -145 19760
rect -225 19695 -145 19700
rect 175 19870 255 19875
rect 175 19810 185 19870
rect 245 19810 255 19870
rect 175 19760 255 19810
rect 175 19700 185 19760
rect 245 19700 255 19760
rect 175 19695 255 19700
rect 575 19870 655 19875
rect 575 19810 585 19870
rect 645 19810 655 19870
rect 575 19760 655 19810
rect 575 19700 585 19760
rect 645 19700 655 19760
rect 575 19695 655 19700
rect 975 19870 1055 19875
rect 975 19810 985 19870
rect 1045 19810 1055 19870
rect 975 19760 1055 19810
rect 975 19700 985 19760
rect 1045 19700 1055 19760
rect 975 19695 1055 19700
rect 1375 19870 1455 19875
rect 1375 19810 1385 19870
rect 1445 19810 1455 19870
rect 1375 19760 1455 19810
rect 1375 19700 1385 19760
rect 1445 19700 1455 19760
rect 1375 19695 1455 19700
rect 1775 19870 1855 19875
rect 1775 19810 1785 19870
rect 1845 19810 1855 19870
rect 1775 19760 1855 19810
rect 1775 19700 1785 19760
rect 1845 19700 1855 19760
rect 1775 19695 1855 19700
rect 2175 19870 2255 19875
rect 2175 19810 2185 19870
rect 2245 19810 2255 19870
rect 2175 19760 2255 19810
rect 2175 19700 2185 19760
rect 2245 19700 2255 19760
rect 2175 19695 2255 19700
rect 2575 19870 2655 19875
rect 2575 19810 2585 19870
rect 2645 19810 2655 19870
rect 2575 19760 2655 19810
rect 2575 19700 2585 19760
rect 2645 19700 2655 19760
rect 2575 19695 2655 19700
rect 2975 19870 3055 19875
rect 2975 19810 2985 19870
rect 3045 19810 3055 19870
rect 2975 19760 3055 19810
rect 2975 19700 2985 19760
rect 3045 19700 3055 19760
rect 2975 19695 3055 19700
rect 3375 19870 3455 19875
rect 3375 19810 3385 19870
rect 3445 19810 3455 19870
rect 3375 19760 3455 19810
rect 3375 19700 3385 19760
rect 3445 19700 3455 19760
rect 3375 19695 3455 19700
rect 3775 19870 3855 19875
rect 3775 19810 3785 19870
rect 3845 19810 3855 19870
rect 3775 19760 3855 19810
rect 3775 19700 3785 19760
rect 3845 19700 3855 19760
rect 3775 19695 3855 19700
rect 4175 19870 4255 19875
rect 4175 19810 4185 19870
rect 4245 19810 4255 19870
rect 4175 19760 4255 19810
rect 4175 19700 4185 19760
rect 4245 19700 4255 19760
rect 4175 19695 4255 19700
rect 4575 19870 4655 19875
rect 4575 19810 4585 19870
rect 4645 19810 4655 19870
rect 4575 19760 4655 19810
rect 4575 19700 4585 19760
rect 4645 19700 4655 19760
rect 4575 19695 4655 19700
rect 4975 19870 5055 19875
rect 4975 19810 4985 19870
rect 5045 19810 5055 19870
rect 4975 19760 5055 19810
rect 4975 19700 4985 19760
rect 5045 19700 5055 19760
rect 4975 19695 5055 19700
rect 5375 19870 5455 19875
rect 5375 19810 5385 19870
rect 5445 19810 5455 19870
rect 5375 19760 5455 19810
rect 5375 19700 5385 19760
rect 5445 19700 5455 19760
rect 5375 19695 5455 19700
rect 5775 19870 5855 19875
rect 5775 19810 5785 19870
rect 5845 19810 5855 19870
rect 5775 19760 5855 19810
rect 5775 19700 5785 19760
rect 5845 19700 5855 19760
rect 5775 19695 5855 19700
rect 6175 19870 6255 19875
rect 6175 19810 6185 19870
rect 6245 19810 6255 19870
rect 6175 19760 6255 19810
rect 6175 19700 6185 19760
rect 6245 19700 6255 19760
rect 6175 19695 6255 19700
rect 6575 19870 6655 19875
rect 6575 19810 6585 19870
rect 6645 19810 6655 19870
rect 6575 19760 6655 19810
rect 6575 19700 6585 19760
rect 6645 19700 6655 19760
rect 6575 19695 6655 19700
rect 6975 19870 7055 19875
rect 6975 19810 6985 19870
rect 7045 19810 7055 19870
rect 6975 19760 7055 19810
rect 6975 19700 6985 19760
rect 7045 19700 7055 19760
rect 6975 19695 7055 19700
rect 7375 19870 7455 19875
rect 7375 19810 7385 19870
rect 7445 19810 7455 19870
rect 7375 19760 7455 19810
rect 7375 19700 7385 19760
rect 7445 19700 7455 19760
rect 7375 19695 7455 19700
rect 7775 19870 7855 19875
rect 7775 19810 7785 19870
rect 7845 19810 7855 19870
rect 7775 19760 7855 19810
rect 7775 19700 7785 19760
rect 7845 19700 7855 19760
rect 7775 19695 7855 19700
rect 8175 19870 8255 19875
rect 8175 19810 8185 19870
rect 8245 19810 8255 19870
rect 8175 19760 8255 19810
rect 8175 19700 8185 19760
rect 8245 19700 8255 19760
rect 8175 19695 8255 19700
rect 8575 19870 8655 19875
rect 8575 19810 8585 19870
rect 8645 19810 8655 19870
rect 8575 19760 8655 19810
rect 8575 19700 8585 19760
rect 8645 19700 8655 19760
rect 8575 19695 8655 19700
rect 8975 19870 9055 19875
rect 8975 19810 8985 19870
rect 9045 19810 9055 19870
rect 8975 19760 9055 19810
rect 8975 19700 8985 19760
rect 9045 19700 9055 19760
rect 8975 19695 9055 19700
rect 9375 19870 9455 19875
rect 9375 19810 9385 19870
rect 9445 19810 9455 19870
rect 9375 19760 9455 19810
rect 9375 19700 9385 19760
rect 9445 19700 9455 19760
rect 9375 19695 9455 19700
rect 9775 19870 9855 19875
rect 9775 19810 9785 19870
rect 9845 19810 9855 19870
rect 9775 19760 9855 19810
rect 9775 19700 9785 19760
rect 9845 19700 9855 19760
rect 9775 19695 9855 19700
rect 10175 19870 10255 19875
rect 10175 19810 10185 19870
rect 10245 19810 10255 19870
rect 10175 19760 10255 19810
rect 10175 19700 10185 19760
rect 10245 19700 10255 19760
rect 10175 19695 10255 19700
rect 10575 19870 10655 19875
rect 10575 19810 10585 19870
rect 10645 19810 10655 19870
rect 10575 19760 10655 19810
rect 10575 19700 10585 19760
rect 10645 19700 10655 19760
rect 10575 19695 10655 19700
rect 10975 19870 11055 19875
rect 10975 19810 10985 19870
rect 11045 19810 11055 19870
rect 10975 19760 11055 19810
rect 10975 19700 10985 19760
rect 11045 19700 11055 19760
rect 10975 19695 11055 19700
rect 11375 19870 11455 19875
rect 11375 19810 11385 19870
rect 11445 19810 11455 19870
rect 11375 19760 11455 19810
rect 11375 19700 11385 19760
rect 11445 19700 11455 19760
rect 11375 19695 11455 19700
rect 11775 19870 11855 19875
rect 11775 19810 11785 19870
rect 11845 19810 11855 19870
rect 11775 19760 11855 19810
rect 11775 19700 11785 19760
rect 11845 19700 11855 19760
rect 11775 19695 11855 19700
rect 12175 19870 12255 19875
rect 12175 19810 12185 19870
rect 12245 19810 12255 19870
rect 12175 19760 12255 19810
rect 12175 19700 12185 19760
rect 12245 19700 12255 19760
rect 12175 19695 12255 19700
rect 12575 19870 12655 19875
rect 12575 19810 12585 19870
rect 12645 19810 12655 19870
rect 12575 19760 12655 19810
rect 12575 19700 12585 19760
rect 12645 19700 12655 19760
rect 12575 19695 12655 19700
rect 12975 19870 13055 19875
rect 12975 19810 12985 19870
rect 13045 19810 13055 19870
rect 12975 19760 13055 19810
rect 12975 19700 12985 19760
rect 13045 19700 13055 19760
rect 12975 19695 13055 19700
rect -215 19505 -155 19695
rect 185 19505 245 19695
rect 585 19505 645 19695
rect 985 19505 1045 19695
rect 1385 19505 1445 19695
rect 1785 19505 1845 19695
rect 2185 19505 2245 19695
rect 2585 19505 2645 19695
rect 2985 19505 3045 19695
rect 3385 19505 3445 19695
rect 3785 19505 3845 19695
rect 4185 19505 4245 19695
rect 4585 19505 4645 19695
rect 4985 19505 5045 19695
rect 5385 19505 5445 19695
rect 5785 19505 5845 19695
rect 6185 19505 6245 19695
rect 6585 19505 6645 19695
rect 6985 19505 7045 19695
rect 7385 19505 7445 19695
rect 7785 19505 7845 19695
rect 8185 19505 8245 19695
rect 8585 19505 8645 19695
rect 8985 19505 9045 19695
rect 9385 19505 9445 19695
rect 9785 19505 9845 19695
rect 10185 19505 10245 19695
rect 10585 19505 10645 19695
rect 10985 19505 11045 19695
rect 11385 19505 11445 19695
rect 11785 19505 11845 19695
rect 12185 19505 12245 19695
rect 12585 19505 12645 19695
rect 12985 19505 13045 19695
rect -225 19500 -145 19505
rect -225 19440 -215 19500
rect -155 19440 -145 19500
rect -225 19390 -145 19440
rect -225 19330 -215 19390
rect -155 19330 -145 19390
rect -225 19325 -145 19330
rect 175 19500 255 19505
rect 175 19440 185 19500
rect 245 19440 255 19500
rect 175 19390 255 19440
rect 175 19330 185 19390
rect 245 19330 255 19390
rect 175 19325 255 19330
rect 575 19500 655 19505
rect 575 19440 585 19500
rect 645 19440 655 19500
rect 575 19390 655 19440
rect 575 19330 585 19390
rect 645 19330 655 19390
rect 575 19325 655 19330
rect 975 19500 1055 19505
rect 975 19440 985 19500
rect 1045 19440 1055 19500
rect 975 19390 1055 19440
rect 975 19330 985 19390
rect 1045 19330 1055 19390
rect 975 19325 1055 19330
rect 1375 19500 1455 19505
rect 1375 19440 1385 19500
rect 1445 19440 1455 19500
rect 1375 19390 1455 19440
rect 1375 19330 1385 19390
rect 1445 19330 1455 19390
rect 1375 19325 1455 19330
rect 1775 19500 1855 19505
rect 1775 19440 1785 19500
rect 1845 19440 1855 19500
rect 1775 19390 1855 19440
rect 1775 19330 1785 19390
rect 1845 19330 1855 19390
rect 1775 19325 1855 19330
rect 2175 19500 2255 19505
rect 2175 19440 2185 19500
rect 2245 19440 2255 19500
rect 2175 19390 2255 19440
rect 2175 19330 2185 19390
rect 2245 19330 2255 19390
rect 2175 19325 2255 19330
rect 2575 19500 2655 19505
rect 2575 19440 2585 19500
rect 2645 19440 2655 19500
rect 2575 19390 2655 19440
rect 2575 19330 2585 19390
rect 2645 19330 2655 19390
rect 2575 19325 2655 19330
rect 2975 19500 3055 19505
rect 2975 19440 2985 19500
rect 3045 19440 3055 19500
rect 2975 19390 3055 19440
rect 2975 19330 2985 19390
rect 3045 19330 3055 19390
rect 2975 19325 3055 19330
rect 3375 19500 3455 19505
rect 3375 19440 3385 19500
rect 3445 19440 3455 19500
rect 3375 19390 3455 19440
rect 3375 19330 3385 19390
rect 3445 19330 3455 19390
rect 3375 19325 3455 19330
rect 3775 19500 3855 19505
rect 3775 19440 3785 19500
rect 3845 19440 3855 19500
rect 3775 19390 3855 19440
rect 3775 19330 3785 19390
rect 3845 19330 3855 19390
rect 3775 19325 3855 19330
rect 4175 19500 4255 19505
rect 4175 19440 4185 19500
rect 4245 19440 4255 19500
rect 4175 19390 4255 19440
rect 4175 19330 4185 19390
rect 4245 19330 4255 19390
rect 4175 19325 4255 19330
rect 4575 19500 4655 19505
rect 4575 19440 4585 19500
rect 4645 19440 4655 19500
rect 4575 19390 4655 19440
rect 4575 19330 4585 19390
rect 4645 19330 4655 19390
rect 4575 19325 4655 19330
rect 4975 19500 5055 19505
rect 4975 19440 4985 19500
rect 5045 19440 5055 19500
rect 4975 19390 5055 19440
rect 4975 19330 4985 19390
rect 5045 19330 5055 19390
rect 4975 19325 5055 19330
rect 5375 19500 5455 19505
rect 5375 19440 5385 19500
rect 5445 19440 5455 19500
rect 5375 19390 5455 19440
rect 5375 19330 5385 19390
rect 5445 19330 5455 19390
rect 5375 19325 5455 19330
rect 5775 19500 5855 19505
rect 5775 19440 5785 19500
rect 5845 19440 5855 19500
rect 5775 19390 5855 19440
rect 5775 19330 5785 19390
rect 5845 19330 5855 19390
rect 5775 19325 5855 19330
rect 6175 19500 6255 19505
rect 6175 19440 6185 19500
rect 6245 19440 6255 19500
rect 6175 19390 6255 19440
rect 6175 19330 6185 19390
rect 6245 19330 6255 19390
rect 6175 19325 6255 19330
rect 6575 19500 6655 19505
rect 6575 19440 6585 19500
rect 6645 19440 6655 19500
rect 6575 19390 6655 19440
rect 6575 19330 6585 19390
rect 6645 19330 6655 19390
rect 6575 19325 6655 19330
rect 6975 19500 7055 19505
rect 6975 19440 6985 19500
rect 7045 19440 7055 19500
rect 6975 19390 7055 19440
rect 6975 19330 6985 19390
rect 7045 19330 7055 19390
rect 6975 19325 7055 19330
rect 7375 19500 7455 19505
rect 7375 19440 7385 19500
rect 7445 19440 7455 19500
rect 7375 19390 7455 19440
rect 7375 19330 7385 19390
rect 7445 19330 7455 19390
rect 7375 19325 7455 19330
rect 7775 19500 7855 19505
rect 7775 19440 7785 19500
rect 7845 19440 7855 19500
rect 7775 19390 7855 19440
rect 7775 19330 7785 19390
rect 7845 19330 7855 19390
rect 7775 19325 7855 19330
rect 8175 19500 8255 19505
rect 8175 19440 8185 19500
rect 8245 19440 8255 19500
rect 8175 19390 8255 19440
rect 8175 19330 8185 19390
rect 8245 19330 8255 19390
rect 8175 19325 8255 19330
rect 8575 19500 8655 19505
rect 8575 19440 8585 19500
rect 8645 19440 8655 19500
rect 8575 19390 8655 19440
rect 8575 19330 8585 19390
rect 8645 19330 8655 19390
rect 8575 19325 8655 19330
rect 8975 19500 9055 19505
rect 8975 19440 8985 19500
rect 9045 19440 9055 19500
rect 8975 19390 9055 19440
rect 8975 19330 8985 19390
rect 9045 19330 9055 19390
rect 8975 19325 9055 19330
rect 9375 19500 9455 19505
rect 9375 19440 9385 19500
rect 9445 19440 9455 19500
rect 9375 19390 9455 19440
rect 9375 19330 9385 19390
rect 9445 19330 9455 19390
rect 9375 19325 9455 19330
rect 9775 19500 9855 19505
rect 9775 19440 9785 19500
rect 9845 19440 9855 19500
rect 9775 19390 9855 19440
rect 9775 19330 9785 19390
rect 9845 19330 9855 19390
rect 9775 19325 9855 19330
rect 10175 19500 10255 19505
rect 10175 19440 10185 19500
rect 10245 19440 10255 19500
rect 10175 19390 10255 19440
rect 10175 19330 10185 19390
rect 10245 19330 10255 19390
rect 10175 19325 10255 19330
rect 10575 19500 10655 19505
rect 10575 19440 10585 19500
rect 10645 19440 10655 19500
rect 10575 19390 10655 19440
rect 10575 19330 10585 19390
rect 10645 19330 10655 19390
rect 10575 19325 10655 19330
rect 10975 19500 11055 19505
rect 10975 19440 10985 19500
rect 11045 19440 11055 19500
rect 10975 19390 11055 19440
rect 10975 19330 10985 19390
rect 11045 19330 11055 19390
rect 10975 19325 11055 19330
rect 11375 19500 11455 19505
rect 11375 19440 11385 19500
rect 11445 19440 11455 19500
rect 11375 19390 11455 19440
rect 11375 19330 11385 19390
rect 11445 19330 11455 19390
rect 11375 19325 11455 19330
rect 11775 19500 11855 19505
rect 11775 19440 11785 19500
rect 11845 19440 11855 19500
rect 11775 19390 11855 19440
rect 11775 19330 11785 19390
rect 11845 19330 11855 19390
rect 11775 19325 11855 19330
rect 12175 19500 12255 19505
rect 12175 19440 12185 19500
rect 12245 19440 12255 19500
rect 12175 19390 12255 19440
rect 12175 19330 12185 19390
rect 12245 19330 12255 19390
rect 12175 19325 12255 19330
rect 12575 19500 12655 19505
rect 12575 19440 12585 19500
rect 12645 19440 12655 19500
rect 12575 19390 12655 19440
rect 12575 19330 12585 19390
rect 12645 19330 12655 19390
rect 12575 19325 12655 19330
rect 12975 19500 13055 19505
rect 12975 19440 12985 19500
rect 13045 19440 13055 19500
rect 12975 19390 13055 19440
rect 12975 19330 12985 19390
rect 13045 19330 13055 19390
rect 12975 19325 13055 19330
rect -215 19135 -155 19325
rect 185 19135 245 19325
rect 585 19135 645 19325
rect 985 19135 1045 19325
rect 1385 19135 1445 19325
rect 1785 19135 1845 19325
rect 2185 19135 2245 19325
rect 2585 19135 2645 19325
rect 2985 19135 3045 19325
rect 3385 19135 3445 19325
rect 3785 19135 3845 19325
rect 4185 19135 4245 19325
rect 4585 19135 4645 19325
rect 4985 19135 5045 19325
rect 5385 19135 5445 19325
rect 5785 19135 5845 19325
rect 6185 19135 6245 19325
rect 6585 19135 6645 19325
rect 6985 19135 7045 19325
rect 7385 19135 7445 19325
rect 7785 19135 7845 19325
rect 8185 19135 8245 19325
rect 8585 19135 8645 19325
rect 8985 19135 9045 19325
rect 9385 19135 9445 19325
rect 9785 19135 9845 19325
rect 10185 19135 10245 19325
rect 10585 19135 10645 19325
rect 10985 19135 11045 19325
rect 11385 19135 11445 19325
rect 11785 19135 11845 19325
rect 12185 19135 12245 19325
rect 12585 19135 12645 19325
rect 12985 19135 13045 19325
rect -225 19130 -145 19135
rect -225 19070 -215 19130
rect -155 19070 -145 19130
rect -225 19020 -145 19070
rect -225 18960 -215 19020
rect -155 18960 -145 19020
rect -225 18955 -145 18960
rect 175 19130 255 19135
rect 175 19070 185 19130
rect 245 19070 255 19130
rect 175 19020 255 19070
rect 175 18960 185 19020
rect 245 18960 255 19020
rect 175 18955 255 18960
rect 575 19130 655 19135
rect 575 19070 585 19130
rect 645 19070 655 19130
rect 575 19020 655 19070
rect 575 18960 585 19020
rect 645 18960 655 19020
rect 575 18955 655 18960
rect 975 19130 1055 19135
rect 975 19070 985 19130
rect 1045 19070 1055 19130
rect 975 19020 1055 19070
rect 975 18960 985 19020
rect 1045 18960 1055 19020
rect 975 18955 1055 18960
rect 1375 19130 1455 19135
rect 1375 19070 1385 19130
rect 1445 19070 1455 19130
rect 1375 19020 1455 19070
rect 1375 18960 1385 19020
rect 1445 18960 1455 19020
rect 1375 18955 1455 18960
rect 1775 19130 1855 19135
rect 1775 19070 1785 19130
rect 1845 19070 1855 19130
rect 1775 19020 1855 19070
rect 1775 18960 1785 19020
rect 1845 18960 1855 19020
rect 1775 18955 1855 18960
rect 2175 19130 2255 19135
rect 2175 19070 2185 19130
rect 2245 19070 2255 19130
rect 2175 19020 2255 19070
rect 2175 18960 2185 19020
rect 2245 18960 2255 19020
rect 2175 18955 2255 18960
rect 2575 19130 2655 19135
rect 2575 19070 2585 19130
rect 2645 19070 2655 19130
rect 2575 19020 2655 19070
rect 2575 18960 2585 19020
rect 2645 18960 2655 19020
rect 2575 18955 2655 18960
rect 2975 19130 3055 19135
rect 2975 19070 2985 19130
rect 3045 19070 3055 19130
rect 2975 19020 3055 19070
rect 2975 18960 2985 19020
rect 3045 18960 3055 19020
rect 2975 18955 3055 18960
rect 3375 19130 3455 19135
rect 3375 19070 3385 19130
rect 3445 19070 3455 19130
rect 3375 19020 3455 19070
rect 3375 18960 3385 19020
rect 3445 18960 3455 19020
rect 3375 18955 3455 18960
rect 3775 19130 3855 19135
rect 3775 19070 3785 19130
rect 3845 19070 3855 19130
rect 3775 19020 3855 19070
rect 3775 18960 3785 19020
rect 3845 18960 3855 19020
rect 3775 18955 3855 18960
rect 4175 19130 4255 19135
rect 4175 19070 4185 19130
rect 4245 19070 4255 19130
rect 4175 19020 4255 19070
rect 4175 18960 4185 19020
rect 4245 18960 4255 19020
rect 4175 18955 4255 18960
rect 4575 19130 4655 19135
rect 4575 19070 4585 19130
rect 4645 19070 4655 19130
rect 4575 19020 4655 19070
rect 4575 18960 4585 19020
rect 4645 18960 4655 19020
rect 4575 18955 4655 18960
rect 4975 19130 5055 19135
rect 4975 19070 4985 19130
rect 5045 19070 5055 19130
rect 4975 19020 5055 19070
rect 4975 18960 4985 19020
rect 5045 18960 5055 19020
rect 4975 18955 5055 18960
rect 5375 19130 5455 19135
rect 5375 19070 5385 19130
rect 5445 19070 5455 19130
rect 5375 19020 5455 19070
rect 5375 18960 5385 19020
rect 5445 18960 5455 19020
rect 5375 18955 5455 18960
rect 5775 19130 5855 19135
rect 5775 19070 5785 19130
rect 5845 19070 5855 19130
rect 5775 19020 5855 19070
rect 5775 18960 5785 19020
rect 5845 18960 5855 19020
rect 5775 18955 5855 18960
rect 6175 19130 6255 19135
rect 6175 19070 6185 19130
rect 6245 19070 6255 19130
rect 6175 19020 6255 19070
rect 6175 18960 6185 19020
rect 6245 18960 6255 19020
rect 6175 18955 6255 18960
rect 6575 19130 6655 19135
rect 6575 19070 6585 19130
rect 6645 19070 6655 19130
rect 6575 19020 6655 19070
rect 6575 18960 6585 19020
rect 6645 18960 6655 19020
rect 6575 18955 6655 18960
rect 6975 19130 7055 19135
rect 6975 19070 6985 19130
rect 7045 19070 7055 19130
rect 6975 19020 7055 19070
rect 6975 18960 6985 19020
rect 7045 18960 7055 19020
rect 6975 18955 7055 18960
rect 7375 19130 7455 19135
rect 7375 19070 7385 19130
rect 7445 19070 7455 19130
rect 7375 19020 7455 19070
rect 7375 18960 7385 19020
rect 7445 18960 7455 19020
rect 7375 18955 7455 18960
rect 7775 19130 7855 19135
rect 7775 19070 7785 19130
rect 7845 19070 7855 19130
rect 7775 19020 7855 19070
rect 7775 18960 7785 19020
rect 7845 18960 7855 19020
rect 7775 18955 7855 18960
rect 8175 19130 8255 19135
rect 8175 19070 8185 19130
rect 8245 19070 8255 19130
rect 8175 19020 8255 19070
rect 8175 18960 8185 19020
rect 8245 18960 8255 19020
rect 8175 18955 8255 18960
rect 8575 19130 8655 19135
rect 8575 19070 8585 19130
rect 8645 19070 8655 19130
rect 8575 19020 8655 19070
rect 8575 18960 8585 19020
rect 8645 18960 8655 19020
rect 8575 18955 8655 18960
rect 8975 19130 9055 19135
rect 8975 19070 8985 19130
rect 9045 19070 9055 19130
rect 8975 19020 9055 19070
rect 8975 18960 8985 19020
rect 9045 18960 9055 19020
rect 8975 18955 9055 18960
rect 9375 19130 9455 19135
rect 9375 19070 9385 19130
rect 9445 19070 9455 19130
rect 9375 19020 9455 19070
rect 9375 18960 9385 19020
rect 9445 18960 9455 19020
rect 9375 18955 9455 18960
rect 9775 19130 9855 19135
rect 9775 19070 9785 19130
rect 9845 19070 9855 19130
rect 9775 19020 9855 19070
rect 9775 18960 9785 19020
rect 9845 18960 9855 19020
rect 9775 18955 9855 18960
rect 10175 19130 10255 19135
rect 10175 19070 10185 19130
rect 10245 19070 10255 19130
rect 10175 19020 10255 19070
rect 10175 18960 10185 19020
rect 10245 18960 10255 19020
rect 10175 18955 10255 18960
rect 10575 19130 10655 19135
rect 10575 19070 10585 19130
rect 10645 19070 10655 19130
rect 10575 19020 10655 19070
rect 10575 18960 10585 19020
rect 10645 18960 10655 19020
rect 10575 18955 10655 18960
rect 10975 19130 11055 19135
rect 10975 19070 10985 19130
rect 11045 19070 11055 19130
rect 10975 19020 11055 19070
rect 10975 18960 10985 19020
rect 11045 18960 11055 19020
rect 10975 18955 11055 18960
rect 11375 19130 11455 19135
rect 11375 19070 11385 19130
rect 11445 19070 11455 19130
rect 11375 19020 11455 19070
rect 11375 18960 11385 19020
rect 11445 18960 11455 19020
rect 11375 18955 11455 18960
rect 11775 19130 11855 19135
rect 11775 19070 11785 19130
rect 11845 19070 11855 19130
rect 11775 19020 11855 19070
rect 11775 18960 11785 19020
rect 11845 18960 11855 19020
rect 11775 18955 11855 18960
rect 12175 19130 12255 19135
rect 12175 19070 12185 19130
rect 12245 19070 12255 19130
rect 12175 19020 12255 19070
rect 12175 18960 12185 19020
rect 12245 18960 12255 19020
rect 12175 18955 12255 18960
rect 12575 19130 12655 19135
rect 12575 19070 12585 19130
rect 12645 19070 12655 19130
rect 12575 19020 12655 19070
rect 12575 18960 12585 19020
rect 12645 18960 12655 19020
rect 12575 18955 12655 18960
rect 12975 19130 13055 19135
rect 12975 19070 12985 19130
rect 13045 19070 13055 19130
rect 12975 19020 13055 19070
rect 12975 18960 12985 19020
rect 13045 18960 13055 19020
rect 12975 18955 13055 18960
rect -215 18765 -155 18955
rect 185 18765 245 18955
rect 585 18765 645 18955
rect 985 18765 1045 18955
rect 1385 18765 1445 18955
rect 1785 18765 1845 18955
rect 2185 18765 2245 18955
rect 2585 18765 2645 18955
rect 2985 18765 3045 18955
rect 3385 18765 3445 18955
rect 3785 18765 3845 18955
rect 4185 18765 4245 18955
rect 4585 18765 4645 18955
rect 4985 18765 5045 18955
rect 5385 18765 5445 18955
rect 5785 18765 5845 18955
rect 6185 18765 6245 18955
rect 6585 18765 6645 18955
rect 6985 18765 7045 18955
rect 7385 18765 7445 18955
rect 7785 18765 7845 18955
rect 8185 18765 8245 18955
rect 8585 18765 8645 18955
rect 8985 18765 9045 18955
rect 9385 18765 9445 18955
rect 9785 18765 9845 18955
rect 10185 18765 10245 18955
rect 10585 18765 10645 18955
rect 10985 18765 11045 18955
rect 11385 18765 11445 18955
rect 11785 18765 11845 18955
rect 12185 18765 12245 18955
rect 12585 18765 12645 18955
rect 12985 18765 13045 18955
rect -225 18760 -145 18765
rect -225 18700 -215 18760
rect -155 18700 -145 18760
rect -225 18650 -145 18700
rect -225 18590 -215 18650
rect -155 18590 -145 18650
rect -225 18585 -145 18590
rect 175 18760 255 18765
rect 175 18700 185 18760
rect 245 18700 255 18760
rect 175 18650 255 18700
rect 175 18590 185 18650
rect 245 18590 255 18650
rect 175 18585 255 18590
rect 575 18760 655 18765
rect 575 18700 585 18760
rect 645 18700 655 18760
rect 575 18650 655 18700
rect 575 18590 585 18650
rect 645 18590 655 18650
rect 575 18585 655 18590
rect 975 18760 1055 18765
rect 975 18700 985 18760
rect 1045 18700 1055 18760
rect 975 18650 1055 18700
rect 975 18590 985 18650
rect 1045 18590 1055 18650
rect 975 18585 1055 18590
rect 1375 18760 1455 18765
rect 1375 18700 1385 18760
rect 1445 18700 1455 18760
rect 1375 18650 1455 18700
rect 1375 18590 1385 18650
rect 1445 18590 1455 18650
rect 1375 18585 1455 18590
rect 1775 18760 1855 18765
rect 1775 18700 1785 18760
rect 1845 18700 1855 18760
rect 1775 18650 1855 18700
rect 1775 18590 1785 18650
rect 1845 18590 1855 18650
rect 1775 18585 1855 18590
rect 2175 18760 2255 18765
rect 2175 18700 2185 18760
rect 2245 18700 2255 18760
rect 2175 18650 2255 18700
rect 2175 18590 2185 18650
rect 2245 18590 2255 18650
rect 2175 18585 2255 18590
rect 2575 18760 2655 18765
rect 2575 18700 2585 18760
rect 2645 18700 2655 18760
rect 2575 18650 2655 18700
rect 2575 18590 2585 18650
rect 2645 18590 2655 18650
rect 2575 18585 2655 18590
rect 2975 18760 3055 18765
rect 2975 18700 2985 18760
rect 3045 18700 3055 18760
rect 2975 18650 3055 18700
rect 2975 18590 2985 18650
rect 3045 18590 3055 18650
rect 2975 18585 3055 18590
rect 3375 18760 3455 18765
rect 3375 18700 3385 18760
rect 3445 18700 3455 18760
rect 3375 18650 3455 18700
rect 3375 18590 3385 18650
rect 3445 18590 3455 18650
rect 3375 18585 3455 18590
rect 3775 18760 3855 18765
rect 3775 18700 3785 18760
rect 3845 18700 3855 18760
rect 3775 18650 3855 18700
rect 3775 18590 3785 18650
rect 3845 18590 3855 18650
rect 3775 18585 3855 18590
rect 4175 18760 4255 18765
rect 4175 18700 4185 18760
rect 4245 18700 4255 18760
rect 4175 18650 4255 18700
rect 4175 18590 4185 18650
rect 4245 18590 4255 18650
rect 4175 18585 4255 18590
rect 4575 18760 4655 18765
rect 4575 18700 4585 18760
rect 4645 18700 4655 18760
rect 4575 18650 4655 18700
rect 4575 18590 4585 18650
rect 4645 18590 4655 18650
rect 4575 18585 4655 18590
rect 4975 18760 5055 18765
rect 4975 18700 4985 18760
rect 5045 18700 5055 18760
rect 4975 18650 5055 18700
rect 4975 18590 4985 18650
rect 5045 18590 5055 18650
rect 4975 18585 5055 18590
rect 5375 18760 5455 18765
rect 5375 18700 5385 18760
rect 5445 18700 5455 18760
rect 5375 18650 5455 18700
rect 5375 18590 5385 18650
rect 5445 18590 5455 18650
rect 5375 18585 5455 18590
rect 5775 18760 5855 18765
rect 5775 18700 5785 18760
rect 5845 18700 5855 18760
rect 5775 18650 5855 18700
rect 5775 18590 5785 18650
rect 5845 18590 5855 18650
rect 5775 18585 5855 18590
rect 6175 18760 6255 18765
rect 6175 18700 6185 18760
rect 6245 18700 6255 18760
rect 6175 18650 6255 18700
rect 6175 18590 6185 18650
rect 6245 18590 6255 18650
rect 6175 18585 6255 18590
rect 6575 18760 6655 18765
rect 6575 18700 6585 18760
rect 6645 18700 6655 18760
rect 6575 18650 6655 18700
rect 6575 18590 6585 18650
rect 6645 18590 6655 18650
rect 6575 18585 6655 18590
rect 6975 18760 7055 18765
rect 6975 18700 6985 18760
rect 7045 18700 7055 18760
rect 6975 18650 7055 18700
rect 6975 18590 6985 18650
rect 7045 18590 7055 18650
rect 6975 18585 7055 18590
rect 7375 18760 7455 18765
rect 7375 18700 7385 18760
rect 7445 18700 7455 18760
rect 7375 18650 7455 18700
rect 7375 18590 7385 18650
rect 7445 18590 7455 18650
rect 7375 18585 7455 18590
rect 7775 18760 7855 18765
rect 7775 18700 7785 18760
rect 7845 18700 7855 18760
rect 7775 18650 7855 18700
rect 7775 18590 7785 18650
rect 7845 18590 7855 18650
rect 7775 18585 7855 18590
rect 8175 18760 8255 18765
rect 8175 18700 8185 18760
rect 8245 18700 8255 18760
rect 8175 18650 8255 18700
rect 8175 18590 8185 18650
rect 8245 18590 8255 18650
rect 8175 18585 8255 18590
rect 8575 18760 8655 18765
rect 8575 18700 8585 18760
rect 8645 18700 8655 18760
rect 8575 18650 8655 18700
rect 8575 18590 8585 18650
rect 8645 18590 8655 18650
rect 8575 18585 8655 18590
rect 8975 18760 9055 18765
rect 8975 18700 8985 18760
rect 9045 18700 9055 18760
rect 8975 18650 9055 18700
rect 8975 18590 8985 18650
rect 9045 18590 9055 18650
rect 8975 18585 9055 18590
rect 9375 18760 9455 18765
rect 9375 18700 9385 18760
rect 9445 18700 9455 18760
rect 9375 18650 9455 18700
rect 9375 18590 9385 18650
rect 9445 18590 9455 18650
rect 9375 18585 9455 18590
rect 9775 18760 9855 18765
rect 9775 18700 9785 18760
rect 9845 18700 9855 18760
rect 9775 18650 9855 18700
rect 9775 18590 9785 18650
rect 9845 18590 9855 18650
rect 9775 18585 9855 18590
rect 10175 18760 10255 18765
rect 10175 18700 10185 18760
rect 10245 18700 10255 18760
rect 10175 18650 10255 18700
rect 10175 18590 10185 18650
rect 10245 18590 10255 18650
rect 10175 18585 10255 18590
rect 10575 18760 10655 18765
rect 10575 18700 10585 18760
rect 10645 18700 10655 18760
rect 10575 18650 10655 18700
rect 10575 18590 10585 18650
rect 10645 18590 10655 18650
rect 10575 18585 10655 18590
rect 10975 18760 11055 18765
rect 10975 18700 10985 18760
rect 11045 18700 11055 18760
rect 10975 18650 11055 18700
rect 10975 18590 10985 18650
rect 11045 18590 11055 18650
rect 10975 18585 11055 18590
rect 11375 18760 11455 18765
rect 11375 18700 11385 18760
rect 11445 18700 11455 18760
rect 11375 18650 11455 18700
rect 11375 18590 11385 18650
rect 11445 18590 11455 18650
rect 11375 18585 11455 18590
rect 11775 18760 11855 18765
rect 11775 18700 11785 18760
rect 11845 18700 11855 18760
rect 11775 18650 11855 18700
rect 11775 18590 11785 18650
rect 11845 18590 11855 18650
rect 11775 18585 11855 18590
rect 12175 18760 12255 18765
rect 12175 18700 12185 18760
rect 12245 18700 12255 18760
rect 12175 18650 12255 18700
rect 12175 18590 12185 18650
rect 12245 18590 12255 18650
rect 12175 18585 12255 18590
rect 12575 18760 12655 18765
rect 12575 18700 12585 18760
rect 12645 18700 12655 18760
rect 12575 18650 12655 18700
rect 12575 18590 12585 18650
rect 12645 18590 12655 18650
rect 12575 18585 12655 18590
rect 12975 18760 13055 18765
rect 12975 18700 12985 18760
rect 13045 18700 13055 18760
rect 12975 18650 13055 18700
rect 12975 18590 12985 18650
rect 13045 18590 13055 18650
rect 12975 18585 13055 18590
rect -215 18395 -155 18585
rect 185 18395 245 18585
rect 585 18395 645 18585
rect 985 18395 1045 18585
rect 1385 18395 1445 18585
rect 1785 18395 1845 18585
rect 2185 18395 2245 18585
rect 2585 18395 2645 18585
rect 2985 18395 3045 18585
rect 3385 18395 3445 18585
rect 3785 18395 3845 18585
rect 4185 18395 4245 18585
rect 4585 18395 4645 18585
rect 4985 18395 5045 18585
rect 5385 18395 5445 18585
rect 5785 18395 5845 18585
rect 6185 18395 6245 18585
rect 6585 18395 6645 18585
rect 6985 18395 7045 18585
rect 7385 18395 7445 18585
rect 7785 18395 7845 18585
rect 8185 18395 8245 18585
rect 8585 18395 8645 18585
rect 8985 18395 9045 18585
rect 9385 18395 9445 18585
rect 9785 18395 9845 18585
rect 10185 18395 10245 18585
rect 10585 18395 10645 18585
rect 10985 18395 11045 18585
rect 11385 18395 11445 18585
rect 11785 18395 11845 18585
rect 12185 18395 12245 18585
rect 12585 18395 12645 18585
rect 12985 18395 13045 18585
rect -225 18390 -145 18395
rect -225 18330 -215 18390
rect -155 18330 -145 18390
rect -225 18280 -145 18330
rect -225 18220 -215 18280
rect -155 18220 -145 18280
rect -225 18215 -145 18220
rect 175 18390 255 18395
rect 175 18330 185 18390
rect 245 18330 255 18390
rect 175 18280 255 18330
rect 175 18220 185 18280
rect 245 18220 255 18280
rect 175 18215 255 18220
rect 575 18390 655 18395
rect 575 18330 585 18390
rect 645 18330 655 18390
rect 575 18280 655 18330
rect 575 18220 585 18280
rect 645 18220 655 18280
rect 575 18215 655 18220
rect 975 18390 1055 18395
rect 975 18330 985 18390
rect 1045 18330 1055 18390
rect 975 18280 1055 18330
rect 975 18220 985 18280
rect 1045 18220 1055 18280
rect 975 18215 1055 18220
rect 1375 18390 1455 18395
rect 1375 18330 1385 18390
rect 1445 18330 1455 18390
rect 1375 18280 1455 18330
rect 1375 18220 1385 18280
rect 1445 18220 1455 18280
rect 1375 18215 1455 18220
rect 1775 18390 1855 18395
rect 1775 18330 1785 18390
rect 1845 18330 1855 18390
rect 1775 18280 1855 18330
rect 1775 18220 1785 18280
rect 1845 18220 1855 18280
rect 1775 18215 1855 18220
rect 2175 18390 2255 18395
rect 2175 18330 2185 18390
rect 2245 18330 2255 18390
rect 2175 18280 2255 18330
rect 2175 18220 2185 18280
rect 2245 18220 2255 18280
rect 2175 18215 2255 18220
rect 2575 18390 2655 18395
rect 2575 18330 2585 18390
rect 2645 18330 2655 18390
rect 2575 18280 2655 18330
rect 2575 18220 2585 18280
rect 2645 18220 2655 18280
rect 2575 18215 2655 18220
rect 2975 18390 3055 18395
rect 2975 18330 2985 18390
rect 3045 18330 3055 18390
rect 2975 18280 3055 18330
rect 2975 18220 2985 18280
rect 3045 18220 3055 18280
rect 2975 18215 3055 18220
rect 3375 18390 3455 18395
rect 3375 18330 3385 18390
rect 3445 18330 3455 18390
rect 3375 18280 3455 18330
rect 3375 18220 3385 18280
rect 3445 18220 3455 18280
rect 3375 18215 3455 18220
rect 3775 18390 3855 18395
rect 3775 18330 3785 18390
rect 3845 18330 3855 18390
rect 3775 18280 3855 18330
rect 3775 18220 3785 18280
rect 3845 18220 3855 18280
rect 3775 18215 3855 18220
rect 4175 18390 4255 18395
rect 4175 18330 4185 18390
rect 4245 18330 4255 18390
rect 4175 18280 4255 18330
rect 4175 18220 4185 18280
rect 4245 18220 4255 18280
rect 4175 18215 4255 18220
rect 4575 18390 4655 18395
rect 4575 18330 4585 18390
rect 4645 18330 4655 18390
rect 4575 18280 4655 18330
rect 4575 18220 4585 18280
rect 4645 18220 4655 18280
rect 4575 18215 4655 18220
rect 4975 18390 5055 18395
rect 4975 18330 4985 18390
rect 5045 18330 5055 18390
rect 4975 18280 5055 18330
rect 4975 18220 4985 18280
rect 5045 18220 5055 18280
rect 4975 18215 5055 18220
rect 5375 18390 5455 18395
rect 5375 18330 5385 18390
rect 5445 18330 5455 18390
rect 5375 18280 5455 18330
rect 5375 18220 5385 18280
rect 5445 18220 5455 18280
rect 5375 18215 5455 18220
rect 5775 18390 5855 18395
rect 5775 18330 5785 18390
rect 5845 18330 5855 18390
rect 5775 18280 5855 18330
rect 5775 18220 5785 18280
rect 5845 18220 5855 18280
rect 5775 18215 5855 18220
rect 6175 18390 6255 18395
rect 6175 18330 6185 18390
rect 6245 18330 6255 18390
rect 6175 18280 6255 18330
rect 6175 18220 6185 18280
rect 6245 18220 6255 18280
rect 6175 18215 6255 18220
rect 6575 18390 6655 18395
rect 6575 18330 6585 18390
rect 6645 18330 6655 18390
rect 6575 18280 6655 18330
rect 6575 18220 6585 18280
rect 6645 18220 6655 18280
rect 6575 18215 6655 18220
rect 6975 18390 7055 18395
rect 6975 18330 6985 18390
rect 7045 18330 7055 18390
rect 6975 18280 7055 18330
rect 6975 18220 6985 18280
rect 7045 18220 7055 18280
rect 6975 18215 7055 18220
rect 7375 18390 7455 18395
rect 7375 18330 7385 18390
rect 7445 18330 7455 18390
rect 7375 18280 7455 18330
rect 7375 18220 7385 18280
rect 7445 18220 7455 18280
rect 7375 18215 7455 18220
rect 7775 18390 7855 18395
rect 7775 18330 7785 18390
rect 7845 18330 7855 18390
rect 7775 18280 7855 18330
rect 7775 18220 7785 18280
rect 7845 18220 7855 18280
rect 7775 18215 7855 18220
rect 8175 18390 8255 18395
rect 8175 18330 8185 18390
rect 8245 18330 8255 18390
rect 8175 18280 8255 18330
rect 8175 18220 8185 18280
rect 8245 18220 8255 18280
rect 8175 18215 8255 18220
rect 8575 18390 8655 18395
rect 8575 18330 8585 18390
rect 8645 18330 8655 18390
rect 8575 18280 8655 18330
rect 8575 18220 8585 18280
rect 8645 18220 8655 18280
rect 8575 18215 8655 18220
rect 8975 18390 9055 18395
rect 8975 18330 8985 18390
rect 9045 18330 9055 18390
rect 8975 18280 9055 18330
rect 8975 18220 8985 18280
rect 9045 18220 9055 18280
rect 8975 18215 9055 18220
rect 9375 18390 9455 18395
rect 9375 18330 9385 18390
rect 9445 18330 9455 18390
rect 9375 18280 9455 18330
rect 9375 18220 9385 18280
rect 9445 18220 9455 18280
rect 9375 18215 9455 18220
rect 9775 18390 9855 18395
rect 9775 18330 9785 18390
rect 9845 18330 9855 18390
rect 9775 18280 9855 18330
rect 9775 18220 9785 18280
rect 9845 18220 9855 18280
rect 9775 18215 9855 18220
rect 10175 18390 10255 18395
rect 10175 18330 10185 18390
rect 10245 18330 10255 18390
rect 10175 18280 10255 18330
rect 10175 18220 10185 18280
rect 10245 18220 10255 18280
rect 10175 18215 10255 18220
rect 10575 18390 10655 18395
rect 10575 18330 10585 18390
rect 10645 18330 10655 18390
rect 10575 18280 10655 18330
rect 10575 18220 10585 18280
rect 10645 18220 10655 18280
rect 10575 18215 10655 18220
rect 10975 18390 11055 18395
rect 10975 18330 10985 18390
rect 11045 18330 11055 18390
rect 10975 18280 11055 18330
rect 10975 18220 10985 18280
rect 11045 18220 11055 18280
rect 10975 18215 11055 18220
rect 11375 18390 11455 18395
rect 11375 18330 11385 18390
rect 11445 18330 11455 18390
rect 11375 18280 11455 18330
rect 11375 18220 11385 18280
rect 11445 18220 11455 18280
rect 11375 18215 11455 18220
rect 11775 18390 11855 18395
rect 11775 18330 11785 18390
rect 11845 18330 11855 18390
rect 11775 18280 11855 18330
rect 11775 18220 11785 18280
rect 11845 18220 11855 18280
rect 11775 18215 11855 18220
rect 12175 18390 12255 18395
rect 12175 18330 12185 18390
rect 12245 18330 12255 18390
rect 12175 18280 12255 18330
rect 12175 18220 12185 18280
rect 12245 18220 12255 18280
rect 12175 18215 12255 18220
rect 12575 18390 12655 18395
rect 12575 18330 12585 18390
rect 12645 18330 12655 18390
rect 12575 18280 12655 18330
rect 12575 18220 12585 18280
rect 12645 18220 12655 18280
rect 12575 18215 12655 18220
rect 12975 18390 13055 18395
rect 12975 18330 12985 18390
rect 13045 18330 13055 18390
rect 12975 18280 13055 18330
rect 12975 18220 12985 18280
rect 13045 18220 13055 18280
rect 12975 18215 13055 18220
rect -215 18025 -155 18215
rect 185 18025 245 18215
rect 585 18025 645 18215
rect 985 18025 1045 18215
rect 1385 18025 1445 18215
rect 1785 18025 1845 18215
rect 2185 18025 2245 18215
rect 2585 18025 2645 18215
rect 2985 18025 3045 18215
rect 3385 18025 3445 18215
rect 3785 18025 3845 18215
rect 4185 18025 4245 18215
rect 4585 18025 4645 18215
rect 4985 18025 5045 18215
rect 5385 18025 5445 18215
rect 5785 18025 5845 18215
rect 6185 18025 6245 18215
rect 6585 18025 6645 18215
rect 6985 18025 7045 18215
rect 7385 18025 7445 18215
rect 7785 18025 7845 18215
rect 8185 18025 8245 18215
rect 8585 18025 8645 18215
rect 8985 18025 9045 18215
rect 9385 18025 9445 18215
rect 9785 18025 9845 18215
rect 10185 18025 10245 18215
rect 10585 18025 10645 18215
rect 10985 18025 11045 18215
rect 11385 18025 11445 18215
rect 11785 18025 11845 18215
rect 12185 18025 12245 18215
rect 12585 18025 12645 18215
rect 12985 18025 13045 18215
rect -225 18020 -145 18025
rect -225 17960 -215 18020
rect -155 17960 -145 18020
rect -225 17910 -145 17960
rect -225 17850 -215 17910
rect -155 17850 -145 17910
rect -225 17845 -145 17850
rect 175 18020 255 18025
rect 175 17960 185 18020
rect 245 17960 255 18020
rect 175 17910 255 17960
rect 175 17850 185 17910
rect 245 17850 255 17910
rect 175 17845 255 17850
rect 575 18020 655 18025
rect 575 17960 585 18020
rect 645 17960 655 18020
rect 575 17910 655 17960
rect 575 17850 585 17910
rect 645 17850 655 17910
rect 575 17845 655 17850
rect 975 18020 1055 18025
rect 975 17960 985 18020
rect 1045 17960 1055 18020
rect 975 17910 1055 17960
rect 975 17850 985 17910
rect 1045 17850 1055 17910
rect 975 17845 1055 17850
rect 1375 18020 1455 18025
rect 1375 17960 1385 18020
rect 1445 17960 1455 18020
rect 1375 17910 1455 17960
rect 1375 17850 1385 17910
rect 1445 17850 1455 17910
rect 1375 17845 1455 17850
rect 1775 18020 1855 18025
rect 1775 17960 1785 18020
rect 1845 17960 1855 18020
rect 1775 17910 1855 17960
rect 1775 17850 1785 17910
rect 1845 17850 1855 17910
rect 1775 17845 1855 17850
rect 2175 18020 2255 18025
rect 2175 17960 2185 18020
rect 2245 17960 2255 18020
rect 2175 17910 2255 17960
rect 2175 17850 2185 17910
rect 2245 17850 2255 17910
rect 2175 17845 2255 17850
rect 2575 18020 2655 18025
rect 2575 17960 2585 18020
rect 2645 17960 2655 18020
rect 2575 17910 2655 17960
rect 2575 17850 2585 17910
rect 2645 17850 2655 17910
rect 2575 17845 2655 17850
rect 2975 18020 3055 18025
rect 2975 17960 2985 18020
rect 3045 17960 3055 18020
rect 2975 17910 3055 17960
rect 2975 17850 2985 17910
rect 3045 17850 3055 17910
rect 2975 17845 3055 17850
rect 3375 18020 3455 18025
rect 3375 17960 3385 18020
rect 3445 17960 3455 18020
rect 3375 17910 3455 17960
rect 3375 17850 3385 17910
rect 3445 17850 3455 17910
rect 3375 17845 3455 17850
rect 3775 18020 3855 18025
rect 3775 17960 3785 18020
rect 3845 17960 3855 18020
rect 3775 17910 3855 17960
rect 3775 17850 3785 17910
rect 3845 17850 3855 17910
rect 3775 17845 3855 17850
rect 4175 18020 4255 18025
rect 4175 17960 4185 18020
rect 4245 17960 4255 18020
rect 4175 17910 4255 17960
rect 4175 17850 4185 17910
rect 4245 17850 4255 17910
rect 4175 17845 4255 17850
rect 4575 18020 4655 18025
rect 4575 17960 4585 18020
rect 4645 17960 4655 18020
rect 4575 17910 4655 17960
rect 4575 17850 4585 17910
rect 4645 17850 4655 17910
rect 4575 17845 4655 17850
rect 4975 18020 5055 18025
rect 4975 17960 4985 18020
rect 5045 17960 5055 18020
rect 4975 17910 5055 17960
rect 4975 17850 4985 17910
rect 5045 17850 5055 17910
rect 4975 17845 5055 17850
rect 5375 18020 5455 18025
rect 5375 17960 5385 18020
rect 5445 17960 5455 18020
rect 5375 17910 5455 17960
rect 5375 17850 5385 17910
rect 5445 17850 5455 17910
rect 5375 17845 5455 17850
rect 5775 18020 5855 18025
rect 5775 17960 5785 18020
rect 5845 17960 5855 18020
rect 5775 17910 5855 17960
rect 5775 17850 5785 17910
rect 5845 17850 5855 17910
rect 5775 17845 5855 17850
rect 6175 18020 6255 18025
rect 6175 17960 6185 18020
rect 6245 17960 6255 18020
rect 6175 17910 6255 17960
rect 6175 17850 6185 17910
rect 6245 17850 6255 17910
rect 6175 17845 6255 17850
rect 6575 18020 6655 18025
rect 6575 17960 6585 18020
rect 6645 17960 6655 18020
rect 6575 17910 6655 17960
rect 6575 17850 6585 17910
rect 6645 17850 6655 17910
rect 6575 17845 6655 17850
rect 6975 18020 7055 18025
rect 6975 17960 6985 18020
rect 7045 17960 7055 18020
rect 6975 17910 7055 17960
rect 6975 17850 6985 17910
rect 7045 17850 7055 17910
rect 6975 17845 7055 17850
rect 7375 18020 7455 18025
rect 7375 17960 7385 18020
rect 7445 17960 7455 18020
rect 7375 17910 7455 17960
rect 7375 17850 7385 17910
rect 7445 17850 7455 17910
rect 7375 17845 7455 17850
rect 7775 18020 7855 18025
rect 7775 17960 7785 18020
rect 7845 17960 7855 18020
rect 7775 17910 7855 17960
rect 7775 17850 7785 17910
rect 7845 17850 7855 17910
rect 7775 17845 7855 17850
rect 8175 18020 8255 18025
rect 8175 17960 8185 18020
rect 8245 17960 8255 18020
rect 8175 17910 8255 17960
rect 8175 17850 8185 17910
rect 8245 17850 8255 17910
rect 8175 17845 8255 17850
rect 8575 18020 8655 18025
rect 8575 17960 8585 18020
rect 8645 17960 8655 18020
rect 8575 17910 8655 17960
rect 8575 17850 8585 17910
rect 8645 17850 8655 17910
rect 8575 17845 8655 17850
rect 8975 18020 9055 18025
rect 8975 17960 8985 18020
rect 9045 17960 9055 18020
rect 8975 17910 9055 17960
rect 8975 17850 8985 17910
rect 9045 17850 9055 17910
rect 8975 17845 9055 17850
rect 9375 18020 9455 18025
rect 9375 17960 9385 18020
rect 9445 17960 9455 18020
rect 9375 17910 9455 17960
rect 9375 17850 9385 17910
rect 9445 17850 9455 17910
rect 9375 17845 9455 17850
rect 9775 18020 9855 18025
rect 9775 17960 9785 18020
rect 9845 17960 9855 18020
rect 9775 17910 9855 17960
rect 9775 17850 9785 17910
rect 9845 17850 9855 17910
rect 9775 17845 9855 17850
rect 10175 18020 10255 18025
rect 10175 17960 10185 18020
rect 10245 17960 10255 18020
rect 10175 17910 10255 17960
rect 10175 17850 10185 17910
rect 10245 17850 10255 17910
rect 10175 17845 10255 17850
rect 10575 18020 10655 18025
rect 10575 17960 10585 18020
rect 10645 17960 10655 18020
rect 10575 17910 10655 17960
rect 10575 17850 10585 17910
rect 10645 17850 10655 17910
rect 10575 17845 10655 17850
rect 10975 18020 11055 18025
rect 10975 17960 10985 18020
rect 11045 17960 11055 18020
rect 10975 17910 11055 17960
rect 10975 17850 10985 17910
rect 11045 17850 11055 17910
rect 10975 17845 11055 17850
rect 11375 18020 11455 18025
rect 11375 17960 11385 18020
rect 11445 17960 11455 18020
rect 11375 17910 11455 17960
rect 11375 17850 11385 17910
rect 11445 17850 11455 17910
rect 11375 17845 11455 17850
rect 11775 18020 11855 18025
rect 11775 17960 11785 18020
rect 11845 17960 11855 18020
rect 11775 17910 11855 17960
rect 11775 17850 11785 17910
rect 11845 17850 11855 17910
rect 11775 17845 11855 17850
rect 12175 18020 12255 18025
rect 12175 17960 12185 18020
rect 12245 17960 12255 18020
rect 12175 17910 12255 17960
rect 12175 17850 12185 17910
rect 12245 17850 12255 17910
rect 12175 17845 12255 17850
rect 12575 18020 12655 18025
rect 12575 17960 12585 18020
rect 12645 17960 12655 18020
rect 12575 17910 12655 17960
rect 12575 17850 12585 17910
rect 12645 17850 12655 17910
rect 12575 17845 12655 17850
rect 12975 18020 13055 18025
rect 12975 17960 12985 18020
rect 13045 17960 13055 18020
rect 12975 17910 13055 17960
rect 12975 17850 12985 17910
rect 13045 17850 13055 17910
rect 12975 17845 13055 17850
rect -215 17655 -155 17845
rect 185 17655 245 17845
rect 585 17655 645 17845
rect 985 17655 1045 17845
rect 1385 17655 1445 17845
rect 1785 17655 1845 17845
rect 2185 17655 2245 17845
rect 2585 17655 2645 17845
rect 2985 17655 3045 17845
rect 3385 17655 3445 17845
rect 3785 17655 3845 17845
rect 4185 17655 4245 17845
rect 4585 17655 4645 17845
rect 4985 17655 5045 17845
rect 5385 17655 5445 17845
rect 5785 17655 5845 17845
rect 6185 17655 6245 17845
rect 6585 17655 6645 17845
rect 6985 17655 7045 17845
rect 7385 17655 7445 17845
rect 7785 17655 7845 17845
rect 8185 17655 8245 17845
rect 8585 17655 8645 17845
rect 8985 17655 9045 17845
rect 9385 17655 9445 17845
rect 9785 17655 9845 17845
rect 10185 17655 10245 17845
rect 10585 17655 10645 17845
rect 10985 17655 11045 17845
rect 11385 17655 11445 17845
rect 11785 17655 11845 17845
rect 12185 17655 12245 17845
rect 12585 17655 12645 17845
rect 12985 17655 13045 17845
rect -225 17650 -145 17655
rect -225 17590 -215 17650
rect -155 17590 -145 17650
rect -225 17540 -145 17590
rect -225 17480 -215 17540
rect -155 17480 -145 17540
rect -225 17475 -145 17480
rect 175 17650 255 17655
rect 175 17590 185 17650
rect 245 17590 255 17650
rect 175 17540 255 17590
rect 175 17480 185 17540
rect 245 17480 255 17540
rect 175 17475 255 17480
rect 575 17650 655 17655
rect 575 17590 585 17650
rect 645 17590 655 17650
rect 575 17540 655 17590
rect 575 17480 585 17540
rect 645 17480 655 17540
rect 575 17475 655 17480
rect 975 17650 1055 17655
rect 975 17590 985 17650
rect 1045 17590 1055 17650
rect 975 17540 1055 17590
rect 975 17480 985 17540
rect 1045 17480 1055 17540
rect 975 17475 1055 17480
rect 1375 17650 1455 17655
rect 1375 17590 1385 17650
rect 1445 17590 1455 17650
rect 1375 17540 1455 17590
rect 1375 17480 1385 17540
rect 1445 17480 1455 17540
rect 1375 17475 1455 17480
rect 1775 17650 1855 17655
rect 1775 17590 1785 17650
rect 1845 17590 1855 17650
rect 1775 17540 1855 17590
rect 1775 17480 1785 17540
rect 1845 17480 1855 17540
rect 1775 17475 1855 17480
rect 2175 17650 2255 17655
rect 2175 17590 2185 17650
rect 2245 17590 2255 17650
rect 2175 17540 2255 17590
rect 2175 17480 2185 17540
rect 2245 17480 2255 17540
rect 2175 17475 2255 17480
rect 2575 17650 2655 17655
rect 2575 17590 2585 17650
rect 2645 17590 2655 17650
rect 2575 17540 2655 17590
rect 2575 17480 2585 17540
rect 2645 17480 2655 17540
rect 2575 17475 2655 17480
rect 2975 17650 3055 17655
rect 2975 17590 2985 17650
rect 3045 17590 3055 17650
rect 2975 17540 3055 17590
rect 2975 17480 2985 17540
rect 3045 17480 3055 17540
rect 2975 17475 3055 17480
rect 3375 17650 3455 17655
rect 3375 17590 3385 17650
rect 3445 17590 3455 17650
rect 3375 17540 3455 17590
rect 3375 17480 3385 17540
rect 3445 17480 3455 17540
rect 3375 17475 3455 17480
rect 3775 17650 3855 17655
rect 3775 17590 3785 17650
rect 3845 17590 3855 17650
rect 3775 17540 3855 17590
rect 3775 17480 3785 17540
rect 3845 17480 3855 17540
rect 3775 17475 3855 17480
rect 4175 17650 4255 17655
rect 4175 17590 4185 17650
rect 4245 17590 4255 17650
rect 4175 17540 4255 17590
rect 4175 17480 4185 17540
rect 4245 17480 4255 17540
rect 4175 17475 4255 17480
rect 4575 17650 4655 17655
rect 4575 17590 4585 17650
rect 4645 17590 4655 17650
rect 4575 17540 4655 17590
rect 4575 17480 4585 17540
rect 4645 17480 4655 17540
rect 4575 17475 4655 17480
rect 4975 17650 5055 17655
rect 4975 17590 4985 17650
rect 5045 17590 5055 17650
rect 4975 17540 5055 17590
rect 4975 17480 4985 17540
rect 5045 17480 5055 17540
rect 4975 17475 5055 17480
rect 5375 17650 5455 17655
rect 5375 17590 5385 17650
rect 5445 17590 5455 17650
rect 5375 17540 5455 17590
rect 5375 17480 5385 17540
rect 5445 17480 5455 17540
rect 5375 17475 5455 17480
rect 5775 17650 5855 17655
rect 5775 17590 5785 17650
rect 5845 17590 5855 17650
rect 5775 17540 5855 17590
rect 5775 17480 5785 17540
rect 5845 17480 5855 17540
rect 5775 17475 5855 17480
rect 6175 17650 6255 17655
rect 6175 17590 6185 17650
rect 6245 17590 6255 17650
rect 6175 17540 6255 17590
rect 6175 17480 6185 17540
rect 6245 17480 6255 17540
rect 6175 17475 6255 17480
rect 6575 17650 6655 17655
rect 6575 17590 6585 17650
rect 6645 17590 6655 17650
rect 6575 17540 6655 17590
rect 6575 17480 6585 17540
rect 6645 17480 6655 17540
rect 6575 17475 6655 17480
rect 6975 17650 7055 17655
rect 6975 17590 6985 17650
rect 7045 17590 7055 17650
rect 6975 17540 7055 17590
rect 6975 17480 6985 17540
rect 7045 17480 7055 17540
rect 6975 17475 7055 17480
rect 7375 17650 7455 17655
rect 7375 17590 7385 17650
rect 7445 17590 7455 17650
rect 7375 17540 7455 17590
rect 7375 17480 7385 17540
rect 7445 17480 7455 17540
rect 7375 17475 7455 17480
rect 7775 17650 7855 17655
rect 7775 17590 7785 17650
rect 7845 17590 7855 17650
rect 7775 17540 7855 17590
rect 7775 17480 7785 17540
rect 7845 17480 7855 17540
rect 7775 17475 7855 17480
rect 8175 17650 8255 17655
rect 8175 17590 8185 17650
rect 8245 17590 8255 17650
rect 8175 17540 8255 17590
rect 8175 17480 8185 17540
rect 8245 17480 8255 17540
rect 8175 17475 8255 17480
rect 8575 17650 8655 17655
rect 8575 17590 8585 17650
rect 8645 17590 8655 17650
rect 8575 17540 8655 17590
rect 8575 17480 8585 17540
rect 8645 17480 8655 17540
rect 8575 17475 8655 17480
rect 8975 17650 9055 17655
rect 8975 17590 8985 17650
rect 9045 17590 9055 17650
rect 8975 17540 9055 17590
rect 8975 17480 8985 17540
rect 9045 17480 9055 17540
rect 8975 17475 9055 17480
rect 9375 17650 9455 17655
rect 9375 17590 9385 17650
rect 9445 17590 9455 17650
rect 9375 17540 9455 17590
rect 9375 17480 9385 17540
rect 9445 17480 9455 17540
rect 9375 17475 9455 17480
rect 9775 17650 9855 17655
rect 9775 17590 9785 17650
rect 9845 17590 9855 17650
rect 9775 17540 9855 17590
rect 9775 17480 9785 17540
rect 9845 17480 9855 17540
rect 9775 17475 9855 17480
rect 10175 17650 10255 17655
rect 10175 17590 10185 17650
rect 10245 17590 10255 17650
rect 10175 17540 10255 17590
rect 10175 17480 10185 17540
rect 10245 17480 10255 17540
rect 10175 17475 10255 17480
rect 10575 17650 10655 17655
rect 10575 17590 10585 17650
rect 10645 17590 10655 17650
rect 10575 17540 10655 17590
rect 10575 17480 10585 17540
rect 10645 17480 10655 17540
rect 10575 17475 10655 17480
rect 10975 17650 11055 17655
rect 10975 17590 10985 17650
rect 11045 17590 11055 17650
rect 10975 17540 11055 17590
rect 10975 17480 10985 17540
rect 11045 17480 11055 17540
rect 10975 17475 11055 17480
rect 11375 17650 11455 17655
rect 11375 17590 11385 17650
rect 11445 17590 11455 17650
rect 11375 17540 11455 17590
rect 11375 17480 11385 17540
rect 11445 17480 11455 17540
rect 11375 17475 11455 17480
rect 11775 17650 11855 17655
rect 11775 17590 11785 17650
rect 11845 17590 11855 17650
rect 11775 17540 11855 17590
rect 11775 17480 11785 17540
rect 11845 17480 11855 17540
rect 11775 17475 11855 17480
rect 12175 17650 12255 17655
rect 12175 17590 12185 17650
rect 12245 17590 12255 17650
rect 12175 17540 12255 17590
rect 12175 17480 12185 17540
rect 12245 17480 12255 17540
rect 12175 17475 12255 17480
rect 12575 17650 12655 17655
rect 12575 17590 12585 17650
rect 12645 17590 12655 17650
rect 12575 17540 12655 17590
rect 12575 17480 12585 17540
rect 12645 17480 12655 17540
rect 12575 17475 12655 17480
rect 12975 17650 13055 17655
rect 12975 17590 12985 17650
rect 13045 17590 13055 17650
rect 12975 17540 13055 17590
rect 12975 17480 12985 17540
rect 13045 17480 13055 17540
rect 12975 17475 13055 17480
rect -215 17285 -155 17475
rect 185 17285 245 17475
rect 585 17285 645 17475
rect 985 17285 1045 17475
rect 1385 17285 1445 17475
rect 1785 17285 1845 17475
rect 2185 17285 2245 17475
rect 2585 17285 2645 17475
rect 2985 17285 3045 17475
rect 3385 17285 3445 17475
rect 3785 17285 3845 17475
rect 4185 17285 4245 17475
rect 4585 17285 4645 17475
rect 4985 17285 5045 17475
rect 5385 17285 5445 17475
rect 5785 17285 5845 17475
rect 6185 17285 6245 17475
rect 6585 17285 6645 17475
rect 6985 17285 7045 17475
rect 7385 17285 7445 17475
rect 7785 17285 7845 17475
rect 8185 17285 8245 17475
rect 8585 17285 8645 17475
rect 8985 17285 9045 17475
rect 9385 17285 9445 17475
rect 9785 17285 9845 17475
rect 10185 17285 10245 17475
rect 10585 17285 10645 17475
rect 10985 17285 11045 17475
rect 11385 17285 11445 17475
rect 11785 17285 11845 17475
rect 12185 17285 12245 17475
rect 12585 17285 12645 17475
rect 12985 17285 13045 17475
rect -225 17280 -145 17285
rect -225 17220 -215 17280
rect -155 17220 -145 17280
rect -225 17170 -145 17220
rect -225 17110 -215 17170
rect -155 17110 -145 17170
rect -225 17105 -145 17110
rect 175 17280 255 17285
rect 175 17220 185 17280
rect 245 17220 255 17280
rect 175 17170 255 17220
rect 175 17110 185 17170
rect 245 17110 255 17170
rect 175 17105 255 17110
rect 575 17280 655 17285
rect 575 17220 585 17280
rect 645 17220 655 17280
rect 575 17170 655 17220
rect 575 17110 585 17170
rect 645 17110 655 17170
rect 575 17105 655 17110
rect 975 17280 1055 17285
rect 975 17220 985 17280
rect 1045 17220 1055 17280
rect 975 17170 1055 17220
rect 975 17110 985 17170
rect 1045 17110 1055 17170
rect 975 17105 1055 17110
rect 1375 17280 1455 17285
rect 1375 17220 1385 17280
rect 1445 17220 1455 17280
rect 1375 17170 1455 17220
rect 1375 17110 1385 17170
rect 1445 17110 1455 17170
rect 1375 17105 1455 17110
rect 1775 17280 1855 17285
rect 1775 17220 1785 17280
rect 1845 17220 1855 17280
rect 1775 17170 1855 17220
rect 1775 17110 1785 17170
rect 1845 17110 1855 17170
rect 1775 17105 1855 17110
rect 2175 17280 2255 17285
rect 2175 17220 2185 17280
rect 2245 17220 2255 17280
rect 2175 17170 2255 17220
rect 2175 17110 2185 17170
rect 2245 17110 2255 17170
rect 2175 17105 2255 17110
rect 2575 17280 2655 17285
rect 2575 17220 2585 17280
rect 2645 17220 2655 17280
rect 2575 17170 2655 17220
rect 2575 17110 2585 17170
rect 2645 17110 2655 17170
rect 2575 17105 2655 17110
rect 2975 17280 3055 17285
rect 2975 17220 2985 17280
rect 3045 17220 3055 17280
rect 2975 17170 3055 17220
rect 2975 17110 2985 17170
rect 3045 17110 3055 17170
rect 2975 17105 3055 17110
rect 3375 17280 3455 17285
rect 3375 17220 3385 17280
rect 3445 17220 3455 17280
rect 3375 17170 3455 17220
rect 3375 17110 3385 17170
rect 3445 17110 3455 17170
rect 3375 17105 3455 17110
rect 3775 17280 3855 17285
rect 3775 17220 3785 17280
rect 3845 17220 3855 17280
rect 3775 17170 3855 17220
rect 3775 17110 3785 17170
rect 3845 17110 3855 17170
rect 3775 17105 3855 17110
rect 4175 17280 4255 17285
rect 4175 17220 4185 17280
rect 4245 17220 4255 17280
rect 4175 17170 4255 17220
rect 4175 17110 4185 17170
rect 4245 17110 4255 17170
rect 4175 17105 4255 17110
rect 4575 17280 4655 17285
rect 4575 17220 4585 17280
rect 4645 17220 4655 17280
rect 4575 17170 4655 17220
rect 4575 17110 4585 17170
rect 4645 17110 4655 17170
rect 4575 17105 4655 17110
rect 4975 17280 5055 17285
rect 4975 17220 4985 17280
rect 5045 17220 5055 17280
rect 4975 17170 5055 17220
rect 4975 17110 4985 17170
rect 5045 17110 5055 17170
rect 4975 17105 5055 17110
rect 5375 17280 5455 17285
rect 5375 17220 5385 17280
rect 5445 17220 5455 17280
rect 5375 17170 5455 17220
rect 5375 17110 5385 17170
rect 5445 17110 5455 17170
rect 5375 17105 5455 17110
rect 5775 17280 5855 17285
rect 5775 17220 5785 17280
rect 5845 17220 5855 17280
rect 5775 17170 5855 17220
rect 5775 17110 5785 17170
rect 5845 17110 5855 17170
rect 5775 17105 5855 17110
rect 6175 17280 6255 17285
rect 6175 17220 6185 17280
rect 6245 17220 6255 17280
rect 6175 17170 6255 17220
rect 6175 17110 6185 17170
rect 6245 17110 6255 17170
rect 6175 17105 6255 17110
rect 6575 17280 6655 17285
rect 6575 17220 6585 17280
rect 6645 17220 6655 17280
rect 6575 17170 6655 17220
rect 6575 17110 6585 17170
rect 6645 17110 6655 17170
rect 6575 17105 6655 17110
rect 6975 17280 7055 17285
rect 6975 17220 6985 17280
rect 7045 17220 7055 17280
rect 6975 17170 7055 17220
rect 6975 17110 6985 17170
rect 7045 17110 7055 17170
rect 6975 17105 7055 17110
rect 7375 17280 7455 17285
rect 7375 17220 7385 17280
rect 7445 17220 7455 17280
rect 7375 17170 7455 17220
rect 7375 17110 7385 17170
rect 7445 17110 7455 17170
rect 7375 17105 7455 17110
rect 7775 17280 7855 17285
rect 7775 17220 7785 17280
rect 7845 17220 7855 17280
rect 7775 17170 7855 17220
rect 7775 17110 7785 17170
rect 7845 17110 7855 17170
rect 7775 17105 7855 17110
rect 8175 17280 8255 17285
rect 8175 17220 8185 17280
rect 8245 17220 8255 17280
rect 8175 17170 8255 17220
rect 8175 17110 8185 17170
rect 8245 17110 8255 17170
rect 8175 17105 8255 17110
rect 8575 17280 8655 17285
rect 8575 17220 8585 17280
rect 8645 17220 8655 17280
rect 8575 17170 8655 17220
rect 8575 17110 8585 17170
rect 8645 17110 8655 17170
rect 8575 17105 8655 17110
rect 8975 17280 9055 17285
rect 8975 17220 8985 17280
rect 9045 17220 9055 17280
rect 8975 17170 9055 17220
rect 8975 17110 8985 17170
rect 9045 17110 9055 17170
rect 8975 17105 9055 17110
rect 9375 17280 9455 17285
rect 9375 17220 9385 17280
rect 9445 17220 9455 17280
rect 9375 17170 9455 17220
rect 9375 17110 9385 17170
rect 9445 17110 9455 17170
rect 9375 17105 9455 17110
rect 9775 17280 9855 17285
rect 9775 17220 9785 17280
rect 9845 17220 9855 17280
rect 9775 17170 9855 17220
rect 9775 17110 9785 17170
rect 9845 17110 9855 17170
rect 9775 17105 9855 17110
rect 10175 17280 10255 17285
rect 10175 17220 10185 17280
rect 10245 17220 10255 17280
rect 10175 17170 10255 17220
rect 10175 17110 10185 17170
rect 10245 17110 10255 17170
rect 10175 17105 10255 17110
rect 10575 17280 10655 17285
rect 10575 17220 10585 17280
rect 10645 17220 10655 17280
rect 10575 17170 10655 17220
rect 10575 17110 10585 17170
rect 10645 17110 10655 17170
rect 10575 17105 10655 17110
rect 10975 17280 11055 17285
rect 10975 17220 10985 17280
rect 11045 17220 11055 17280
rect 10975 17170 11055 17220
rect 10975 17110 10985 17170
rect 11045 17110 11055 17170
rect 10975 17105 11055 17110
rect 11375 17280 11455 17285
rect 11375 17220 11385 17280
rect 11445 17220 11455 17280
rect 11375 17170 11455 17220
rect 11375 17110 11385 17170
rect 11445 17110 11455 17170
rect 11375 17105 11455 17110
rect 11775 17280 11855 17285
rect 11775 17220 11785 17280
rect 11845 17220 11855 17280
rect 11775 17170 11855 17220
rect 11775 17110 11785 17170
rect 11845 17110 11855 17170
rect 11775 17105 11855 17110
rect 12175 17280 12255 17285
rect 12175 17220 12185 17280
rect 12245 17220 12255 17280
rect 12175 17170 12255 17220
rect 12175 17110 12185 17170
rect 12245 17110 12255 17170
rect 12175 17105 12255 17110
rect 12575 17280 12655 17285
rect 12575 17220 12585 17280
rect 12645 17220 12655 17280
rect 12575 17170 12655 17220
rect 12575 17110 12585 17170
rect 12645 17110 12655 17170
rect 12575 17105 12655 17110
rect 12975 17280 13055 17285
rect 12975 17220 12985 17280
rect 13045 17220 13055 17280
rect 12975 17170 13055 17220
rect 12975 17110 12985 17170
rect 13045 17110 13055 17170
rect 12975 17105 13055 17110
rect -215 16915 -155 17105
rect 185 16915 245 17105
rect 585 16915 645 17105
rect 985 16915 1045 17105
rect 1385 16915 1445 17105
rect 1785 16915 1845 17105
rect 2185 16915 2245 17105
rect 2585 16915 2645 17105
rect 2985 16915 3045 17105
rect 3385 16915 3445 17105
rect 3785 16915 3845 17105
rect 4185 16915 4245 17105
rect 4585 16915 4645 17105
rect 4985 16915 5045 17105
rect 5385 16915 5445 17105
rect 5785 16915 5845 17105
rect 6185 16915 6245 17105
rect 6585 16915 6645 17105
rect 6985 16915 7045 17105
rect 7385 16915 7445 17105
rect 7785 16915 7845 17105
rect 8185 16915 8245 17105
rect 8585 16915 8645 17105
rect 8985 16915 9045 17105
rect 9385 16915 9445 17105
rect 9785 16915 9845 17105
rect 10185 16915 10245 17105
rect 10585 16915 10645 17105
rect 10985 16915 11045 17105
rect 11385 16915 11445 17105
rect 11785 16915 11845 17105
rect 12185 16915 12245 17105
rect 12585 16915 12645 17105
rect 12985 16915 13045 17105
rect -225 16910 -145 16915
rect -225 16850 -215 16910
rect -155 16850 -145 16910
rect -225 16800 -145 16850
rect -225 16740 -215 16800
rect -155 16740 -145 16800
rect -225 16735 -145 16740
rect 175 16910 255 16915
rect 175 16850 185 16910
rect 245 16850 255 16910
rect 175 16800 255 16850
rect 175 16740 185 16800
rect 245 16740 255 16800
rect 175 16735 255 16740
rect 575 16910 655 16915
rect 575 16850 585 16910
rect 645 16850 655 16910
rect 575 16800 655 16850
rect 575 16740 585 16800
rect 645 16740 655 16800
rect 575 16735 655 16740
rect 975 16910 1055 16915
rect 975 16850 985 16910
rect 1045 16850 1055 16910
rect 975 16800 1055 16850
rect 975 16740 985 16800
rect 1045 16740 1055 16800
rect 975 16735 1055 16740
rect 1375 16910 1455 16915
rect 1375 16850 1385 16910
rect 1445 16850 1455 16910
rect 1375 16800 1455 16850
rect 1375 16740 1385 16800
rect 1445 16740 1455 16800
rect 1375 16735 1455 16740
rect 1775 16910 1855 16915
rect 1775 16850 1785 16910
rect 1845 16850 1855 16910
rect 1775 16800 1855 16850
rect 1775 16740 1785 16800
rect 1845 16740 1855 16800
rect 1775 16735 1855 16740
rect 2175 16910 2255 16915
rect 2175 16850 2185 16910
rect 2245 16850 2255 16910
rect 2175 16800 2255 16850
rect 2175 16740 2185 16800
rect 2245 16740 2255 16800
rect 2175 16735 2255 16740
rect 2575 16910 2655 16915
rect 2575 16850 2585 16910
rect 2645 16850 2655 16910
rect 2575 16800 2655 16850
rect 2575 16740 2585 16800
rect 2645 16740 2655 16800
rect 2575 16735 2655 16740
rect 2975 16910 3055 16915
rect 2975 16850 2985 16910
rect 3045 16850 3055 16910
rect 2975 16800 3055 16850
rect 2975 16740 2985 16800
rect 3045 16740 3055 16800
rect 2975 16735 3055 16740
rect 3375 16910 3455 16915
rect 3375 16850 3385 16910
rect 3445 16850 3455 16910
rect 3375 16800 3455 16850
rect 3375 16740 3385 16800
rect 3445 16740 3455 16800
rect 3375 16735 3455 16740
rect 3775 16910 3855 16915
rect 3775 16850 3785 16910
rect 3845 16850 3855 16910
rect 3775 16800 3855 16850
rect 3775 16740 3785 16800
rect 3845 16740 3855 16800
rect 3775 16735 3855 16740
rect 4175 16910 4255 16915
rect 4175 16850 4185 16910
rect 4245 16850 4255 16910
rect 4175 16800 4255 16850
rect 4175 16740 4185 16800
rect 4245 16740 4255 16800
rect 4175 16735 4255 16740
rect 4575 16910 4655 16915
rect 4575 16850 4585 16910
rect 4645 16850 4655 16910
rect 4575 16800 4655 16850
rect 4575 16740 4585 16800
rect 4645 16740 4655 16800
rect 4575 16735 4655 16740
rect 4975 16910 5055 16915
rect 4975 16850 4985 16910
rect 5045 16850 5055 16910
rect 4975 16800 5055 16850
rect 4975 16740 4985 16800
rect 5045 16740 5055 16800
rect 4975 16735 5055 16740
rect 5375 16910 5455 16915
rect 5375 16850 5385 16910
rect 5445 16850 5455 16910
rect 5375 16800 5455 16850
rect 5375 16740 5385 16800
rect 5445 16740 5455 16800
rect 5375 16735 5455 16740
rect 5775 16910 5855 16915
rect 5775 16850 5785 16910
rect 5845 16850 5855 16910
rect 5775 16800 5855 16850
rect 5775 16740 5785 16800
rect 5845 16740 5855 16800
rect 5775 16735 5855 16740
rect 6175 16910 6255 16915
rect 6175 16850 6185 16910
rect 6245 16850 6255 16910
rect 6175 16800 6255 16850
rect 6175 16740 6185 16800
rect 6245 16740 6255 16800
rect 6175 16735 6255 16740
rect 6575 16910 6655 16915
rect 6575 16850 6585 16910
rect 6645 16850 6655 16910
rect 6575 16800 6655 16850
rect 6575 16740 6585 16800
rect 6645 16740 6655 16800
rect 6575 16735 6655 16740
rect 6975 16910 7055 16915
rect 6975 16850 6985 16910
rect 7045 16850 7055 16910
rect 6975 16800 7055 16850
rect 6975 16740 6985 16800
rect 7045 16740 7055 16800
rect 6975 16735 7055 16740
rect 7375 16910 7455 16915
rect 7375 16850 7385 16910
rect 7445 16850 7455 16910
rect 7375 16800 7455 16850
rect 7375 16740 7385 16800
rect 7445 16740 7455 16800
rect 7375 16735 7455 16740
rect 7775 16910 7855 16915
rect 7775 16850 7785 16910
rect 7845 16850 7855 16910
rect 7775 16800 7855 16850
rect 7775 16740 7785 16800
rect 7845 16740 7855 16800
rect 7775 16735 7855 16740
rect 8175 16910 8255 16915
rect 8175 16850 8185 16910
rect 8245 16850 8255 16910
rect 8175 16800 8255 16850
rect 8175 16740 8185 16800
rect 8245 16740 8255 16800
rect 8175 16735 8255 16740
rect 8575 16910 8655 16915
rect 8575 16850 8585 16910
rect 8645 16850 8655 16910
rect 8575 16800 8655 16850
rect 8575 16740 8585 16800
rect 8645 16740 8655 16800
rect 8575 16735 8655 16740
rect 8975 16910 9055 16915
rect 8975 16850 8985 16910
rect 9045 16850 9055 16910
rect 8975 16800 9055 16850
rect 8975 16740 8985 16800
rect 9045 16740 9055 16800
rect 8975 16735 9055 16740
rect 9375 16910 9455 16915
rect 9375 16850 9385 16910
rect 9445 16850 9455 16910
rect 9375 16800 9455 16850
rect 9375 16740 9385 16800
rect 9445 16740 9455 16800
rect 9375 16735 9455 16740
rect 9775 16910 9855 16915
rect 9775 16850 9785 16910
rect 9845 16850 9855 16910
rect 9775 16800 9855 16850
rect 9775 16740 9785 16800
rect 9845 16740 9855 16800
rect 9775 16735 9855 16740
rect 10175 16910 10255 16915
rect 10175 16850 10185 16910
rect 10245 16850 10255 16910
rect 10175 16800 10255 16850
rect 10175 16740 10185 16800
rect 10245 16740 10255 16800
rect 10175 16735 10255 16740
rect 10575 16910 10655 16915
rect 10575 16850 10585 16910
rect 10645 16850 10655 16910
rect 10575 16800 10655 16850
rect 10575 16740 10585 16800
rect 10645 16740 10655 16800
rect 10575 16735 10655 16740
rect 10975 16910 11055 16915
rect 10975 16850 10985 16910
rect 11045 16850 11055 16910
rect 10975 16800 11055 16850
rect 10975 16740 10985 16800
rect 11045 16740 11055 16800
rect 10975 16735 11055 16740
rect 11375 16910 11455 16915
rect 11375 16850 11385 16910
rect 11445 16850 11455 16910
rect 11375 16800 11455 16850
rect 11375 16740 11385 16800
rect 11445 16740 11455 16800
rect 11375 16735 11455 16740
rect 11775 16910 11855 16915
rect 11775 16850 11785 16910
rect 11845 16850 11855 16910
rect 11775 16800 11855 16850
rect 11775 16740 11785 16800
rect 11845 16740 11855 16800
rect 11775 16735 11855 16740
rect 12175 16910 12255 16915
rect 12175 16850 12185 16910
rect 12245 16850 12255 16910
rect 12175 16800 12255 16850
rect 12175 16740 12185 16800
rect 12245 16740 12255 16800
rect 12175 16735 12255 16740
rect 12575 16910 12655 16915
rect 12575 16850 12585 16910
rect 12645 16850 12655 16910
rect 12575 16800 12655 16850
rect 12575 16740 12585 16800
rect 12645 16740 12655 16800
rect 12575 16735 12655 16740
rect 12975 16910 13055 16915
rect 12975 16850 12985 16910
rect 13045 16850 13055 16910
rect 12975 16800 13055 16850
rect 12975 16740 12985 16800
rect 13045 16740 13055 16800
rect 12975 16735 13055 16740
rect -215 16545 -155 16735
rect 185 16545 245 16735
rect 585 16545 645 16735
rect 985 16545 1045 16735
rect 1385 16545 1445 16735
rect 1785 16545 1845 16735
rect 2185 16545 2245 16735
rect 2585 16545 2645 16735
rect 2985 16545 3045 16735
rect 3385 16545 3445 16735
rect 3785 16545 3845 16735
rect 4185 16545 4245 16735
rect 4585 16545 4645 16735
rect 4985 16545 5045 16735
rect 5385 16545 5445 16735
rect 5785 16545 5845 16735
rect 6185 16545 6245 16735
rect 6585 16545 6645 16735
rect 6985 16545 7045 16735
rect 7385 16545 7445 16735
rect 7785 16545 7845 16735
rect 8185 16545 8245 16735
rect 8585 16545 8645 16735
rect 8985 16545 9045 16735
rect 9385 16545 9445 16735
rect 9785 16545 9845 16735
rect 10185 16545 10245 16735
rect 10585 16545 10645 16735
rect 10985 16545 11045 16735
rect 11385 16545 11445 16735
rect 11785 16545 11845 16735
rect 12185 16545 12245 16735
rect 12585 16545 12645 16735
rect 12985 16545 13045 16735
rect -225 16540 -145 16545
rect -225 16480 -215 16540
rect -155 16480 -145 16540
rect -225 16430 -145 16480
rect -225 16370 -215 16430
rect -155 16370 -145 16430
rect -225 16365 -145 16370
rect 175 16540 255 16545
rect 175 16480 185 16540
rect 245 16480 255 16540
rect 175 16430 255 16480
rect 175 16370 185 16430
rect 245 16370 255 16430
rect 175 16365 255 16370
rect 575 16540 655 16545
rect 575 16480 585 16540
rect 645 16480 655 16540
rect 575 16430 655 16480
rect 575 16370 585 16430
rect 645 16370 655 16430
rect 575 16365 655 16370
rect 975 16540 1055 16545
rect 975 16480 985 16540
rect 1045 16480 1055 16540
rect 975 16430 1055 16480
rect 975 16370 985 16430
rect 1045 16370 1055 16430
rect 975 16365 1055 16370
rect 1375 16540 1455 16545
rect 1375 16480 1385 16540
rect 1445 16480 1455 16540
rect 1375 16430 1455 16480
rect 1375 16370 1385 16430
rect 1445 16370 1455 16430
rect 1375 16365 1455 16370
rect 1775 16540 1855 16545
rect 1775 16480 1785 16540
rect 1845 16480 1855 16540
rect 1775 16430 1855 16480
rect 1775 16370 1785 16430
rect 1845 16370 1855 16430
rect 1775 16365 1855 16370
rect 2175 16540 2255 16545
rect 2175 16480 2185 16540
rect 2245 16480 2255 16540
rect 2175 16430 2255 16480
rect 2175 16370 2185 16430
rect 2245 16370 2255 16430
rect 2175 16365 2255 16370
rect 2575 16540 2655 16545
rect 2575 16480 2585 16540
rect 2645 16480 2655 16540
rect 2575 16430 2655 16480
rect 2575 16370 2585 16430
rect 2645 16370 2655 16430
rect 2575 16365 2655 16370
rect 2975 16540 3055 16545
rect 2975 16480 2985 16540
rect 3045 16480 3055 16540
rect 2975 16430 3055 16480
rect 2975 16370 2985 16430
rect 3045 16370 3055 16430
rect 2975 16365 3055 16370
rect 3375 16540 3455 16545
rect 3375 16480 3385 16540
rect 3445 16480 3455 16540
rect 3375 16430 3455 16480
rect 3375 16370 3385 16430
rect 3445 16370 3455 16430
rect 3375 16365 3455 16370
rect 3775 16540 3855 16545
rect 3775 16480 3785 16540
rect 3845 16480 3855 16540
rect 3775 16430 3855 16480
rect 3775 16370 3785 16430
rect 3845 16370 3855 16430
rect 3775 16365 3855 16370
rect 4175 16540 4255 16545
rect 4175 16480 4185 16540
rect 4245 16480 4255 16540
rect 4175 16430 4255 16480
rect 4175 16370 4185 16430
rect 4245 16370 4255 16430
rect 4175 16365 4255 16370
rect 4575 16540 4655 16545
rect 4575 16480 4585 16540
rect 4645 16480 4655 16540
rect 4575 16430 4655 16480
rect 4575 16370 4585 16430
rect 4645 16370 4655 16430
rect 4575 16365 4655 16370
rect 4975 16540 5055 16545
rect 4975 16480 4985 16540
rect 5045 16480 5055 16540
rect 4975 16430 5055 16480
rect 4975 16370 4985 16430
rect 5045 16370 5055 16430
rect 4975 16365 5055 16370
rect 5375 16540 5455 16545
rect 5375 16480 5385 16540
rect 5445 16480 5455 16540
rect 5375 16430 5455 16480
rect 5375 16370 5385 16430
rect 5445 16370 5455 16430
rect 5375 16365 5455 16370
rect 5775 16540 5855 16545
rect 5775 16480 5785 16540
rect 5845 16480 5855 16540
rect 5775 16430 5855 16480
rect 5775 16370 5785 16430
rect 5845 16370 5855 16430
rect 5775 16365 5855 16370
rect 6175 16540 6255 16545
rect 6175 16480 6185 16540
rect 6245 16480 6255 16540
rect 6175 16430 6255 16480
rect 6175 16370 6185 16430
rect 6245 16370 6255 16430
rect 6175 16365 6255 16370
rect 6575 16540 6655 16545
rect 6575 16480 6585 16540
rect 6645 16480 6655 16540
rect 6575 16430 6655 16480
rect 6575 16370 6585 16430
rect 6645 16370 6655 16430
rect 6575 16365 6655 16370
rect 6975 16540 7055 16545
rect 6975 16480 6985 16540
rect 7045 16480 7055 16540
rect 6975 16430 7055 16480
rect 6975 16370 6985 16430
rect 7045 16370 7055 16430
rect 6975 16365 7055 16370
rect 7375 16540 7455 16545
rect 7375 16480 7385 16540
rect 7445 16480 7455 16540
rect 7375 16430 7455 16480
rect 7375 16370 7385 16430
rect 7445 16370 7455 16430
rect 7375 16365 7455 16370
rect 7775 16540 7855 16545
rect 7775 16480 7785 16540
rect 7845 16480 7855 16540
rect 7775 16430 7855 16480
rect 7775 16370 7785 16430
rect 7845 16370 7855 16430
rect 7775 16365 7855 16370
rect 8175 16540 8255 16545
rect 8175 16480 8185 16540
rect 8245 16480 8255 16540
rect 8175 16430 8255 16480
rect 8175 16370 8185 16430
rect 8245 16370 8255 16430
rect 8175 16365 8255 16370
rect 8575 16540 8655 16545
rect 8575 16480 8585 16540
rect 8645 16480 8655 16540
rect 8575 16430 8655 16480
rect 8575 16370 8585 16430
rect 8645 16370 8655 16430
rect 8575 16365 8655 16370
rect 8975 16540 9055 16545
rect 8975 16480 8985 16540
rect 9045 16480 9055 16540
rect 8975 16430 9055 16480
rect 8975 16370 8985 16430
rect 9045 16370 9055 16430
rect 8975 16365 9055 16370
rect 9375 16540 9455 16545
rect 9375 16480 9385 16540
rect 9445 16480 9455 16540
rect 9375 16430 9455 16480
rect 9375 16370 9385 16430
rect 9445 16370 9455 16430
rect 9375 16365 9455 16370
rect 9775 16540 9855 16545
rect 9775 16480 9785 16540
rect 9845 16480 9855 16540
rect 9775 16430 9855 16480
rect 9775 16370 9785 16430
rect 9845 16370 9855 16430
rect 9775 16365 9855 16370
rect 10175 16540 10255 16545
rect 10175 16480 10185 16540
rect 10245 16480 10255 16540
rect 10175 16430 10255 16480
rect 10175 16370 10185 16430
rect 10245 16370 10255 16430
rect 10175 16365 10255 16370
rect 10575 16540 10655 16545
rect 10575 16480 10585 16540
rect 10645 16480 10655 16540
rect 10575 16430 10655 16480
rect 10575 16370 10585 16430
rect 10645 16370 10655 16430
rect 10575 16365 10655 16370
rect 10975 16540 11055 16545
rect 10975 16480 10985 16540
rect 11045 16480 11055 16540
rect 10975 16430 11055 16480
rect 10975 16370 10985 16430
rect 11045 16370 11055 16430
rect 10975 16365 11055 16370
rect 11375 16540 11455 16545
rect 11375 16480 11385 16540
rect 11445 16480 11455 16540
rect 11375 16430 11455 16480
rect 11375 16370 11385 16430
rect 11445 16370 11455 16430
rect 11375 16365 11455 16370
rect 11775 16540 11855 16545
rect 11775 16480 11785 16540
rect 11845 16480 11855 16540
rect 11775 16430 11855 16480
rect 11775 16370 11785 16430
rect 11845 16370 11855 16430
rect 11775 16365 11855 16370
rect 12175 16540 12255 16545
rect 12175 16480 12185 16540
rect 12245 16480 12255 16540
rect 12175 16430 12255 16480
rect 12175 16370 12185 16430
rect 12245 16370 12255 16430
rect 12175 16365 12255 16370
rect 12575 16540 12655 16545
rect 12575 16480 12585 16540
rect 12645 16480 12655 16540
rect 12575 16430 12655 16480
rect 12575 16370 12585 16430
rect 12645 16370 12655 16430
rect 12575 16365 12655 16370
rect 12975 16540 13055 16545
rect 12975 16480 12985 16540
rect 13045 16480 13055 16540
rect 12975 16430 13055 16480
rect 12975 16370 12985 16430
rect 13045 16370 13055 16430
rect 12975 16365 13055 16370
rect -215 16175 -155 16365
rect 185 16175 245 16365
rect 585 16175 645 16365
rect 985 16175 1045 16365
rect 1385 16175 1445 16365
rect 1785 16175 1845 16365
rect 2185 16175 2245 16365
rect 2585 16175 2645 16365
rect 2985 16175 3045 16365
rect 3385 16175 3445 16365
rect 3785 16175 3845 16365
rect 4185 16175 4245 16365
rect 4585 16175 4645 16365
rect 4985 16175 5045 16365
rect 5385 16175 5445 16365
rect 5785 16175 5845 16365
rect 6185 16175 6245 16365
rect 6585 16175 6645 16365
rect 6985 16175 7045 16365
rect 7385 16175 7445 16365
rect 7785 16175 7845 16365
rect 8185 16175 8245 16365
rect 8585 16175 8645 16365
rect 8985 16175 9045 16365
rect 9385 16175 9445 16365
rect 9785 16175 9845 16365
rect 10185 16175 10245 16365
rect 10585 16175 10645 16365
rect 10985 16175 11045 16365
rect 11385 16175 11445 16365
rect 11785 16175 11845 16365
rect 12185 16175 12245 16365
rect 12585 16175 12645 16365
rect 12985 16175 13045 16365
rect -225 16170 -145 16175
rect -225 16110 -215 16170
rect -155 16110 -145 16170
rect -225 16060 -145 16110
rect -225 16000 -215 16060
rect -155 16000 -145 16060
rect -225 15995 -145 16000
rect 175 16170 255 16175
rect 175 16110 185 16170
rect 245 16110 255 16170
rect 175 16060 255 16110
rect 175 16000 185 16060
rect 245 16000 255 16060
rect 175 15995 255 16000
rect 575 16170 655 16175
rect 575 16110 585 16170
rect 645 16110 655 16170
rect 575 16060 655 16110
rect 575 16000 585 16060
rect 645 16000 655 16060
rect 575 15995 655 16000
rect 975 16170 1055 16175
rect 975 16110 985 16170
rect 1045 16110 1055 16170
rect 975 16060 1055 16110
rect 975 16000 985 16060
rect 1045 16000 1055 16060
rect 975 15995 1055 16000
rect 1375 16170 1455 16175
rect 1375 16110 1385 16170
rect 1445 16110 1455 16170
rect 1375 16060 1455 16110
rect 1375 16000 1385 16060
rect 1445 16000 1455 16060
rect 1375 15995 1455 16000
rect 1775 16170 1855 16175
rect 1775 16110 1785 16170
rect 1845 16110 1855 16170
rect 1775 16060 1855 16110
rect 1775 16000 1785 16060
rect 1845 16000 1855 16060
rect 1775 15995 1855 16000
rect 2175 16170 2255 16175
rect 2175 16110 2185 16170
rect 2245 16110 2255 16170
rect 2175 16060 2255 16110
rect 2175 16000 2185 16060
rect 2245 16000 2255 16060
rect 2175 15995 2255 16000
rect 2575 16170 2655 16175
rect 2575 16110 2585 16170
rect 2645 16110 2655 16170
rect 2575 16060 2655 16110
rect 2575 16000 2585 16060
rect 2645 16000 2655 16060
rect 2575 15995 2655 16000
rect 2975 16170 3055 16175
rect 2975 16110 2985 16170
rect 3045 16110 3055 16170
rect 2975 16060 3055 16110
rect 2975 16000 2985 16060
rect 3045 16000 3055 16060
rect 2975 15995 3055 16000
rect 3375 16170 3455 16175
rect 3375 16110 3385 16170
rect 3445 16110 3455 16170
rect 3375 16060 3455 16110
rect 3375 16000 3385 16060
rect 3445 16000 3455 16060
rect 3375 15995 3455 16000
rect 3775 16170 3855 16175
rect 3775 16110 3785 16170
rect 3845 16110 3855 16170
rect 3775 16060 3855 16110
rect 3775 16000 3785 16060
rect 3845 16000 3855 16060
rect 3775 15995 3855 16000
rect 4175 16170 4255 16175
rect 4175 16110 4185 16170
rect 4245 16110 4255 16170
rect 4175 16060 4255 16110
rect 4175 16000 4185 16060
rect 4245 16000 4255 16060
rect 4175 15995 4255 16000
rect 4575 16170 4655 16175
rect 4575 16110 4585 16170
rect 4645 16110 4655 16170
rect 4575 16060 4655 16110
rect 4575 16000 4585 16060
rect 4645 16000 4655 16060
rect 4575 15995 4655 16000
rect 4975 16170 5055 16175
rect 4975 16110 4985 16170
rect 5045 16110 5055 16170
rect 4975 16060 5055 16110
rect 4975 16000 4985 16060
rect 5045 16000 5055 16060
rect 4975 15995 5055 16000
rect 5375 16170 5455 16175
rect 5375 16110 5385 16170
rect 5445 16110 5455 16170
rect 5375 16060 5455 16110
rect 5375 16000 5385 16060
rect 5445 16000 5455 16060
rect 5375 15995 5455 16000
rect 5775 16170 5855 16175
rect 5775 16110 5785 16170
rect 5845 16110 5855 16170
rect 5775 16060 5855 16110
rect 5775 16000 5785 16060
rect 5845 16000 5855 16060
rect 5775 15995 5855 16000
rect 6175 16170 6255 16175
rect 6175 16110 6185 16170
rect 6245 16110 6255 16170
rect 6175 16060 6255 16110
rect 6175 16000 6185 16060
rect 6245 16000 6255 16060
rect 6175 15995 6255 16000
rect 6575 16170 6655 16175
rect 6575 16110 6585 16170
rect 6645 16110 6655 16170
rect 6575 16060 6655 16110
rect 6575 16000 6585 16060
rect 6645 16000 6655 16060
rect 6575 15995 6655 16000
rect 6975 16170 7055 16175
rect 6975 16110 6985 16170
rect 7045 16110 7055 16170
rect 6975 16060 7055 16110
rect 6975 16000 6985 16060
rect 7045 16000 7055 16060
rect 6975 15995 7055 16000
rect 7375 16170 7455 16175
rect 7375 16110 7385 16170
rect 7445 16110 7455 16170
rect 7375 16060 7455 16110
rect 7375 16000 7385 16060
rect 7445 16000 7455 16060
rect 7375 15995 7455 16000
rect 7775 16170 7855 16175
rect 7775 16110 7785 16170
rect 7845 16110 7855 16170
rect 7775 16060 7855 16110
rect 7775 16000 7785 16060
rect 7845 16000 7855 16060
rect 7775 15995 7855 16000
rect 8175 16170 8255 16175
rect 8175 16110 8185 16170
rect 8245 16110 8255 16170
rect 8175 16060 8255 16110
rect 8175 16000 8185 16060
rect 8245 16000 8255 16060
rect 8175 15995 8255 16000
rect 8575 16170 8655 16175
rect 8575 16110 8585 16170
rect 8645 16110 8655 16170
rect 8575 16060 8655 16110
rect 8575 16000 8585 16060
rect 8645 16000 8655 16060
rect 8575 15995 8655 16000
rect 8975 16170 9055 16175
rect 8975 16110 8985 16170
rect 9045 16110 9055 16170
rect 8975 16060 9055 16110
rect 8975 16000 8985 16060
rect 9045 16000 9055 16060
rect 8975 15995 9055 16000
rect 9375 16170 9455 16175
rect 9375 16110 9385 16170
rect 9445 16110 9455 16170
rect 9375 16060 9455 16110
rect 9375 16000 9385 16060
rect 9445 16000 9455 16060
rect 9375 15995 9455 16000
rect 9775 16170 9855 16175
rect 9775 16110 9785 16170
rect 9845 16110 9855 16170
rect 9775 16060 9855 16110
rect 9775 16000 9785 16060
rect 9845 16000 9855 16060
rect 9775 15995 9855 16000
rect 10175 16170 10255 16175
rect 10175 16110 10185 16170
rect 10245 16110 10255 16170
rect 10175 16060 10255 16110
rect 10175 16000 10185 16060
rect 10245 16000 10255 16060
rect 10175 15995 10255 16000
rect 10575 16170 10655 16175
rect 10575 16110 10585 16170
rect 10645 16110 10655 16170
rect 10575 16060 10655 16110
rect 10575 16000 10585 16060
rect 10645 16000 10655 16060
rect 10575 15995 10655 16000
rect 10975 16170 11055 16175
rect 10975 16110 10985 16170
rect 11045 16110 11055 16170
rect 10975 16060 11055 16110
rect 10975 16000 10985 16060
rect 11045 16000 11055 16060
rect 10975 15995 11055 16000
rect 11375 16170 11455 16175
rect 11375 16110 11385 16170
rect 11445 16110 11455 16170
rect 11375 16060 11455 16110
rect 11375 16000 11385 16060
rect 11445 16000 11455 16060
rect 11375 15995 11455 16000
rect 11775 16170 11855 16175
rect 11775 16110 11785 16170
rect 11845 16110 11855 16170
rect 11775 16060 11855 16110
rect 11775 16000 11785 16060
rect 11845 16000 11855 16060
rect 11775 15995 11855 16000
rect 12175 16170 12255 16175
rect 12175 16110 12185 16170
rect 12245 16110 12255 16170
rect 12175 16060 12255 16110
rect 12175 16000 12185 16060
rect 12245 16000 12255 16060
rect 12175 15995 12255 16000
rect 12575 16170 12655 16175
rect 12575 16110 12585 16170
rect 12645 16110 12655 16170
rect 12575 16060 12655 16110
rect 12575 16000 12585 16060
rect 12645 16000 12655 16060
rect 12575 15995 12655 16000
rect 12975 16170 13055 16175
rect 12975 16110 12985 16170
rect 13045 16110 13055 16170
rect 12975 16060 13055 16110
rect 12975 16000 12985 16060
rect 13045 16000 13055 16060
rect 12975 15995 13055 16000
rect -215 15805 -155 15995
rect 185 15805 245 15995
rect 585 15805 645 15995
rect 985 15805 1045 15995
rect 1385 15805 1445 15995
rect 1785 15805 1845 15995
rect 2185 15805 2245 15995
rect 2585 15805 2645 15995
rect 2985 15805 3045 15995
rect 3385 15805 3445 15995
rect 3785 15805 3845 15995
rect 4185 15805 4245 15995
rect 4585 15805 4645 15995
rect 4985 15805 5045 15995
rect 5385 15805 5445 15995
rect 5785 15805 5845 15995
rect 6185 15805 6245 15995
rect 6585 15805 6645 15995
rect 6985 15805 7045 15995
rect 7385 15805 7445 15995
rect 7785 15805 7845 15995
rect 8185 15805 8245 15995
rect 8585 15805 8645 15995
rect 8985 15805 9045 15995
rect 9385 15805 9445 15995
rect 9785 15805 9845 15995
rect 10185 15805 10245 15995
rect 10585 15805 10645 15995
rect 10985 15805 11045 15995
rect 11385 15805 11445 15995
rect 11785 15805 11845 15995
rect 12185 15805 12245 15995
rect 12585 15805 12645 15995
rect 12985 15805 13045 15995
rect -225 15800 -145 15805
rect -225 15740 -215 15800
rect -155 15740 -145 15800
rect -225 15690 -145 15740
rect -225 15630 -215 15690
rect -155 15630 -145 15690
rect -225 15625 -145 15630
rect 175 15800 255 15805
rect 175 15740 185 15800
rect 245 15740 255 15800
rect 175 15690 255 15740
rect 175 15630 185 15690
rect 245 15630 255 15690
rect 175 15625 255 15630
rect 575 15800 655 15805
rect 575 15740 585 15800
rect 645 15740 655 15800
rect 575 15690 655 15740
rect 575 15630 585 15690
rect 645 15630 655 15690
rect 575 15625 655 15630
rect 975 15800 1055 15805
rect 975 15740 985 15800
rect 1045 15740 1055 15800
rect 975 15690 1055 15740
rect 975 15630 985 15690
rect 1045 15630 1055 15690
rect 975 15625 1055 15630
rect 1375 15800 1455 15805
rect 1375 15740 1385 15800
rect 1445 15740 1455 15800
rect 1375 15690 1455 15740
rect 1375 15630 1385 15690
rect 1445 15630 1455 15690
rect 1375 15625 1455 15630
rect 1775 15800 1855 15805
rect 1775 15740 1785 15800
rect 1845 15740 1855 15800
rect 1775 15690 1855 15740
rect 1775 15630 1785 15690
rect 1845 15630 1855 15690
rect 1775 15625 1855 15630
rect 2175 15800 2255 15805
rect 2175 15740 2185 15800
rect 2245 15740 2255 15800
rect 2175 15690 2255 15740
rect 2175 15630 2185 15690
rect 2245 15630 2255 15690
rect 2175 15625 2255 15630
rect 2575 15800 2655 15805
rect 2575 15740 2585 15800
rect 2645 15740 2655 15800
rect 2575 15690 2655 15740
rect 2575 15630 2585 15690
rect 2645 15630 2655 15690
rect 2575 15625 2655 15630
rect 2975 15800 3055 15805
rect 2975 15740 2985 15800
rect 3045 15740 3055 15800
rect 2975 15690 3055 15740
rect 2975 15630 2985 15690
rect 3045 15630 3055 15690
rect 2975 15625 3055 15630
rect 3375 15800 3455 15805
rect 3375 15740 3385 15800
rect 3445 15740 3455 15800
rect 3375 15690 3455 15740
rect 3375 15630 3385 15690
rect 3445 15630 3455 15690
rect 3375 15625 3455 15630
rect 3775 15800 3855 15805
rect 3775 15740 3785 15800
rect 3845 15740 3855 15800
rect 3775 15690 3855 15740
rect 3775 15630 3785 15690
rect 3845 15630 3855 15690
rect 3775 15625 3855 15630
rect 4175 15800 4255 15805
rect 4175 15740 4185 15800
rect 4245 15740 4255 15800
rect 4175 15690 4255 15740
rect 4175 15630 4185 15690
rect 4245 15630 4255 15690
rect 4175 15625 4255 15630
rect 4575 15800 4655 15805
rect 4575 15740 4585 15800
rect 4645 15740 4655 15800
rect 4575 15690 4655 15740
rect 4575 15630 4585 15690
rect 4645 15630 4655 15690
rect 4575 15625 4655 15630
rect 4975 15800 5055 15805
rect 4975 15740 4985 15800
rect 5045 15740 5055 15800
rect 4975 15690 5055 15740
rect 4975 15630 4985 15690
rect 5045 15630 5055 15690
rect 4975 15625 5055 15630
rect 5375 15800 5455 15805
rect 5375 15740 5385 15800
rect 5445 15740 5455 15800
rect 5375 15690 5455 15740
rect 5375 15630 5385 15690
rect 5445 15630 5455 15690
rect 5375 15625 5455 15630
rect 5775 15800 5855 15805
rect 5775 15740 5785 15800
rect 5845 15740 5855 15800
rect 5775 15690 5855 15740
rect 5775 15630 5785 15690
rect 5845 15630 5855 15690
rect 5775 15625 5855 15630
rect 6175 15800 6255 15805
rect 6175 15740 6185 15800
rect 6245 15740 6255 15800
rect 6175 15690 6255 15740
rect 6175 15630 6185 15690
rect 6245 15630 6255 15690
rect 6175 15625 6255 15630
rect 6575 15800 6655 15805
rect 6575 15740 6585 15800
rect 6645 15740 6655 15800
rect 6575 15690 6655 15740
rect 6575 15630 6585 15690
rect 6645 15630 6655 15690
rect 6575 15625 6655 15630
rect 6975 15800 7055 15805
rect 6975 15740 6985 15800
rect 7045 15740 7055 15800
rect 6975 15690 7055 15740
rect 6975 15630 6985 15690
rect 7045 15630 7055 15690
rect 6975 15625 7055 15630
rect 7375 15800 7455 15805
rect 7375 15740 7385 15800
rect 7445 15740 7455 15800
rect 7375 15690 7455 15740
rect 7375 15630 7385 15690
rect 7445 15630 7455 15690
rect 7375 15625 7455 15630
rect 7775 15800 7855 15805
rect 7775 15740 7785 15800
rect 7845 15740 7855 15800
rect 7775 15690 7855 15740
rect 7775 15630 7785 15690
rect 7845 15630 7855 15690
rect 7775 15625 7855 15630
rect 8175 15800 8255 15805
rect 8175 15740 8185 15800
rect 8245 15740 8255 15800
rect 8175 15690 8255 15740
rect 8175 15630 8185 15690
rect 8245 15630 8255 15690
rect 8175 15625 8255 15630
rect 8575 15800 8655 15805
rect 8575 15740 8585 15800
rect 8645 15740 8655 15800
rect 8575 15690 8655 15740
rect 8575 15630 8585 15690
rect 8645 15630 8655 15690
rect 8575 15625 8655 15630
rect 8975 15800 9055 15805
rect 8975 15740 8985 15800
rect 9045 15740 9055 15800
rect 8975 15690 9055 15740
rect 8975 15630 8985 15690
rect 9045 15630 9055 15690
rect 8975 15625 9055 15630
rect 9375 15800 9455 15805
rect 9375 15740 9385 15800
rect 9445 15740 9455 15800
rect 9375 15690 9455 15740
rect 9375 15630 9385 15690
rect 9445 15630 9455 15690
rect 9375 15625 9455 15630
rect 9775 15800 9855 15805
rect 9775 15740 9785 15800
rect 9845 15740 9855 15800
rect 9775 15690 9855 15740
rect 9775 15630 9785 15690
rect 9845 15630 9855 15690
rect 9775 15625 9855 15630
rect 10175 15800 10255 15805
rect 10175 15740 10185 15800
rect 10245 15740 10255 15800
rect 10175 15690 10255 15740
rect 10175 15630 10185 15690
rect 10245 15630 10255 15690
rect 10175 15625 10255 15630
rect 10575 15800 10655 15805
rect 10575 15740 10585 15800
rect 10645 15740 10655 15800
rect 10575 15690 10655 15740
rect 10575 15630 10585 15690
rect 10645 15630 10655 15690
rect 10575 15625 10655 15630
rect 10975 15800 11055 15805
rect 10975 15740 10985 15800
rect 11045 15740 11055 15800
rect 10975 15690 11055 15740
rect 10975 15630 10985 15690
rect 11045 15630 11055 15690
rect 10975 15625 11055 15630
rect 11375 15800 11455 15805
rect 11375 15740 11385 15800
rect 11445 15740 11455 15800
rect 11375 15690 11455 15740
rect 11375 15630 11385 15690
rect 11445 15630 11455 15690
rect 11375 15625 11455 15630
rect 11775 15800 11855 15805
rect 11775 15740 11785 15800
rect 11845 15740 11855 15800
rect 11775 15690 11855 15740
rect 11775 15630 11785 15690
rect 11845 15630 11855 15690
rect 11775 15625 11855 15630
rect 12175 15800 12255 15805
rect 12175 15740 12185 15800
rect 12245 15740 12255 15800
rect 12175 15690 12255 15740
rect 12175 15630 12185 15690
rect 12245 15630 12255 15690
rect 12175 15625 12255 15630
rect 12575 15800 12655 15805
rect 12575 15740 12585 15800
rect 12645 15740 12655 15800
rect 12575 15690 12655 15740
rect 12575 15630 12585 15690
rect 12645 15630 12655 15690
rect 12575 15625 12655 15630
rect 12975 15800 13055 15805
rect 12975 15740 12985 15800
rect 13045 15740 13055 15800
rect 12975 15690 13055 15740
rect 12975 15630 12985 15690
rect 13045 15630 13055 15690
rect 12975 15625 13055 15630
rect -215 15435 -155 15625
rect 185 15435 245 15625
rect 585 15435 645 15625
rect 985 15435 1045 15625
rect 1385 15435 1445 15625
rect 1785 15435 1845 15625
rect 2185 15435 2245 15625
rect 2585 15435 2645 15625
rect 2985 15435 3045 15625
rect 3385 15435 3445 15625
rect 3785 15435 3845 15625
rect 4185 15435 4245 15625
rect 4585 15435 4645 15625
rect 4985 15435 5045 15625
rect 5385 15435 5445 15625
rect 5785 15435 5845 15625
rect 6185 15435 6245 15625
rect 6585 15435 6645 15625
rect 6985 15435 7045 15625
rect 7385 15435 7445 15625
rect 7785 15435 7845 15625
rect 8185 15435 8245 15625
rect 8585 15435 8645 15625
rect 8985 15435 9045 15625
rect 9385 15435 9445 15625
rect 9785 15435 9845 15625
rect 10185 15435 10245 15625
rect 10585 15435 10645 15625
rect 10985 15435 11045 15625
rect 11385 15435 11445 15625
rect 11785 15435 11845 15625
rect 12185 15435 12245 15625
rect 12585 15435 12645 15625
rect 12985 15435 13045 15625
rect -225 15430 -145 15435
rect -225 15370 -215 15430
rect -155 15370 -145 15430
rect -225 15320 -145 15370
rect -225 15260 -215 15320
rect -155 15260 -145 15320
rect -225 15255 -145 15260
rect 175 15430 255 15435
rect 175 15370 185 15430
rect 245 15370 255 15430
rect 175 15320 255 15370
rect 175 15260 185 15320
rect 245 15260 255 15320
rect 175 15255 255 15260
rect 575 15430 655 15435
rect 575 15370 585 15430
rect 645 15370 655 15430
rect 575 15320 655 15370
rect 575 15260 585 15320
rect 645 15260 655 15320
rect 575 15255 655 15260
rect 975 15430 1055 15435
rect 975 15370 985 15430
rect 1045 15370 1055 15430
rect 975 15320 1055 15370
rect 975 15260 985 15320
rect 1045 15260 1055 15320
rect 975 15255 1055 15260
rect 1375 15430 1455 15435
rect 1375 15370 1385 15430
rect 1445 15370 1455 15430
rect 1375 15320 1455 15370
rect 1375 15260 1385 15320
rect 1445 15260 1455 15320
rect 1375 15255 1455 15260
rect 1775 15430 1855 15435
rect 1775 15370 1785 15430
rect 1845 15370 1855 15430
rect 1775 15320 1855 15370
rect 1775 15260 1785 15320
rect 1845 15260 1855 15320
rect 1775 15255 1855 15260
rect 2175 15430 2255 15435
rect 2175 15370 2185 15430
rect 2245 15370 2255 15430
rect 2175 15320 2255 15370
rect 2175 15260 2185 15320
rect 2245 15260 2255 15320
rect 2175 15255 2255 15260
rect 2575 15430 2655 15435
rect 2575 15370 2585 15430
rect 2645 15370 2655 15430
rect 2575 15320 2655 15370
rect 2575 15260 2585 15320
rect 2645 15260 2655 15320
rect 2575 15255 2655 15260
rect 2975 15430 3055 15435
rect 2975 15370 2985 15430
rect 3045 15370 3055 15430
rect 2975 15320 3055 15370
rect 2975 15260 2985 15320
rect 3045 15260 3055 15320
rect 2975 15255 3055 15260
rect 3375 15430 3455 15435
rect 3375 15370 3385 15430
rect 3445 15370 3455 15430
rect 3375 15320 3455 15370
rect 3375 15260 3385 15320
rect 3445 15260 3455 15320
rect 3375 15255 3455 15260
rect 3775 15430 3855 15435
rect 3775 15370 3785 15430
rect 3845 15370 3855 15430
rect 3775 15320 3855 15370
rect 3775 15260 3785 15320
rect 3845 15260 3855 15320
rect 3775 15255 3855 15260
rect 4175 15430 4255 15435
rect 4175 15370 4185 15430
rect 4245 15370 4255 15430
rect 4175 15320 4255 15370
rect 4175 15260 4185 15320
rect 4245 15260 4255 15320
rect 4175 15255 4255 15260
rect 4575 15430 4655 15435
rect 4575 15370 4585 15430
rect 4645 15370 4655 15430
rect 4575 15320 4655 15370
rect 4575 15260 4585 15320
rect 4645 15260 4655 15320
rect 4575 15255 4655 15260
rect 4975 15430 5055 15435
rect 4975 15370 4985 15430
rect 5045 15370 5055 15430
rect 4975 15320 5055 15370
rect 4975 15260 4985 15320
rect 5045 15260 5055 15320
rect 4975 15255 5055 15260
rect 5375 15430 5455 15435
rect 5375 15370 5385 15430
rect 5445 15370 5455 15430
rect 5375 15320 5455 15370
rect 5375 15260 5385 15320
rect 5445 15260 5455 15320
rect 5375 15255 5455 15260
rect 5775 15430 5855 15435
rect 5775 15370 5785 15430
rect 5845 15370 5855 15430
rect 5775 15320 5855 15370
rect 5775 15260 5785 15320
rect 5845 15260 5855 15320
rect 5775 15255 5855 15260
rect 6175 15430 6255 15435
rect 6175 15370 6185 15430
rect 6245 15370 6255 15430
rect 6175 15320 6255 15370
rect 6175 15260 6185 15320
rect 6245 15260 6255 15320
rect 6175 15255 6255 15260
rect 6575 15430 6655 15435
rect 6575 15370 6585 15430
rect 6645 15370 6655 15430
rect 6575 15320 6655 15370
rect 6575 15260 6585 15320
rect 6645 15260 6655 15320
rect 6575 15255 6655 15260
rect 6975 15430 7055 15435
rect 6975 15370 6985 15430
rect 7045 15370 7055 15430
rect 6975 15320 7055 15370
rect 6975 15260 6985 15320
rect 7045 15260 7055 15320
rect 6975 15255 7055 15260
rect 7375 15430 7455 15435
rect 7375 15370 7385 15430
rect 7445 15370 7455 15430
rect 7375 15320 7455 15370
rect 7375 15260 7385 15320
rect 7445 15260 7455 15320
rect 7375 15255 7455 15260
rect 7775 15430 7855 15435
rect 7775 15370 7785 15430
rect 7845 15370 7855 15430
rect 7775 15320 7855 15370
rect 7775 15260 7785 15320
rect 7845 15260 7855 15320
rect 7775 15255 7855 15260
rect 8175 15430 8255 15435
rect 8175 15370 8185 15430
rect 8245 15370 8255 15430
rect 8175 15320 8255 15370
rect 8175 15260 8185 15320
rect 8245 15260 8255 15320
rect 8175 15255 8255 15260
rect 8575 15430 8655 15435
rect 8575 15370 8585 15430
rect 8645 15370 8655 15430
rect 8575 15320 8655 15370
rect 8575 15260 8585 15320
rect 8645 15260 8655 15320
rect 8575 15255 8655 15260
rect 8975 15430 9055 15435
rect 8975 15370 8985 15430
rect 9045 15370 9055 15430
rect 8975 15320 9055 15370
rect 8975 15260 8985 15320
rect 9045 15260 9055 15320
rect 8975 15255 9055 15260
rect 9375 15430 9455 15435
rect 9375 15370 9385 15430
rect 9445 15370 9455 15430
rect 9375 15320 9455 15370
rect 9375 15260 9385 15320
rect 9445 15260 9455 15320
rect 9375 15255 9455 15260
rect 9775 15430 9855 15435
rect 9775 15370 9785 15430
rect 9845 15370 9855 15430
rect 9775 15320 9855 15370
rect 9775 15260 9785 15320
rect 9845 15260 9855 15320
rect 9775 15255 9855 15260
rect 10175 15430 10255 15435
rect 10175 15370 10185 15430
rect 10245 15370 10255 15430
rect 10175 15320 10255 15370
rect 10175 15260 10185 15320
rect 10245 15260 10255 15320
rect 10175 15255 10255 15260
rect 10575 15430 10655 15435
rect 10575 15370 10585 15430
rect 10645 15370 10655 15430
rect 10575 15320 10655 15370
rect 10575 15260 10585 15320
rect 10645 15260 10655 15320
rect 10575 15255 10655 15260
rect 10975 15430 11055 15435
rect 10975 15370 10985 15430
rect 11045 15370 11055 15430
rect 10975 15320 11055 15370
rect 10975 15260 10985 15320
rect 11045 15260 11055 15320
rect 10975 15255 11055 15260
rect 11375 15430 11455 15435
rect 11375 15370 11385 15430
rect 11445 15370 11455 15430
rect 11375 15320 11455 15370
rect 11375 15260 11385 15320
rect 11445 15260 11455 15320
rect 11375 15255 11455 15260
rect 11775 15430 11855 15435
rect 11775 15370 11785 15430
rect 11845 15370 11855 15430
rect 11775 15320 11855 15370
rect 11775 15260 11785 15320
rect 11845 15260 11855 15320
rect 11775 15255 11855 15260
rect 12175 15430 12255 15435
rect 12175 15370 12185 15430
rect 12245 15370 12255 15430
rect 12175 15320 12255 15370
rect 12175 15260 12185 15320
rect 12245 15260 12255 15320
rect 12175 15255 12255 15260
rect 12575 15430 12655 15435
rect 12575 15370 12585 15430
rect 12645 15370 12655 15430
rect 12575 15320 12655 15370
rect 12575 15260 12585 15320
rect 12645 15260 12655 15320
rect 12575 15255 12655 15260
rect 12975 15430 13055 15435
rect 12975 15370 12985 15430
rect 13045 15370 13055 15430
rect 12975 15320 13055 15370
rect 12975 15260 12985 15320
rect 13045 15260 13055 15320
rect 12975 15255 13055 15260
rect -215 15065 -155 15255
rect 185 15065 245 15255
rect 585 15065 645 15255
rect 985 15065 1045 15255
rect 1385 15065 1445 15255
rect 1785 15065 1845 15255
rect 2185 15065 2245 15255
rect 2585 15065 2645 15255
rect 2985 15065 3045 15255
rect 3385 15065 3445 15255
rect 3785 15065 3845 15255
rect 4185 15065 4245 15255
rect 4585 15065 4645 15255
rect 4985 15065 5045 15255
rect 5385 15065 5445 15255
rect 5785 15065 5845 15255
rect 6185 15065 6245 15255
rect 6585 15065 6645 15255
rect 6985 15065 7045 15255
rect 7385 15065 7445 15255
rect 7785 15065 7845 15255
rect 8185 15065 8245 15255
rect 8585 15065 8645 15255
rect 8985 15065 9045 15255
rect 9385 15065 9445 15255
rect 9785 15065 9845 15255
rect 10185 15065 10245 15255
rect 10585 15065 10645 15255
rect 10985 15065 11045 15255
rect 11385 15065 11445 15255
rect 11785 15065 11845 15255
rect 12185 15065 12245 15255
rect 12585 15065 12645 15255
rect 12985 15065 13045 15255
rect -225 15060 -145 15065
rect -225 15000 -215 15060
rect -155 15000 -145 15060
rect -225 14950 -145 15000
rect -225 14890 -215 14950
rect -155 14890 -145 14950
rect -225 14885 -145 14890
rect 175 15060 255 15065
rect 175 15000 185 15060
rect 245 15000 255 15060
rect 175 14950 255 15000
rect 175 14890 185 14950
rect 245 14890 255 14950
rect 175 14885 255 14890
rect 575 15060 655 15065
rect 575 15000 585 15060
rect 645 15000 655 15060
rect 575 14950 655 15000
rect 575 14890 585 14950
rect 645 14890 655 14950
rect 575 14885 655 14890
rect 975 15060 1055 15065
rect 975 15000 985 15060
rect 1045 15000 1055 15060
rect 975 14950 1055 15000
rect 975 14890 985 14950
rect 1045 14890 1055 14950
rect 975 14885 1055 14890
rect 1375 15060 1455 15065
rect 1375 15000 1385 15060
rect 1445 15000 1455 15060
rect 1375 14950 1455 15000
rect 1375 14890 1385 14950
rect 1445 14890 1455 14950
rect 1375 14885 1455 14890
rect 1775 15060 1855 15065
rect 1775 15000 1785 15060
rect 1845 15000 1855 15060
rect 1775 14950 1855 15000
rect 1775 14890 1785 14950
rect 1845 14890 1855 14950
rect 1775 14885 1855 14890
rect 2175 15060 2255 15065
rect 2175 15000 2185 15060
rect 2245 15000 2255 15060
rect 2175 14950 2255 15000
rect 2175 14890 2185 14950
rect 2245 14890 2255 14950
rect 2175 14885 2255 14890
rect 2575 15060 2655 15065
rect 2575 15000 2585 15060
rect 2645 15000 2655 15060
rect 2575 14950 2655 15000
rect 2575 14890 2585 14950
rect 2645 14890 2655 14950
rect 2575 14885 2655 14890
rect 2975 15060 3055 15065
rect 2975 15000 2985 15060
rect 3045 15000 3055 15060
rect 2975 14950 3055 15000
rect 2975 14890 2985 14950
rect 3045 14890 3055 14950
rect 2975 14885 3055 14890
rect 3375 15060 3455 15065
rect 3375 15000 3385 15060
rect 3445 15000 3455 15060
rect 3375 14950 3455 15000
rect 3375 14890 3385 14950
rect 3445 14890 3455 14950
rect 3375 14885 3455 14890
rect 3775 15060 3855 15065
rect 3775 15000 3785 15060
rect 3845 15000 3855 15060
rect 3775 14950 3855 15000
rect 3775 14890 3785 14950
rect 3845 14890 3855 14950
rect 3775 14885 3855 14890
rect 4175 15060 4255 15065
rect 4175 15000 4185 15060
rect 4245 15000 4255 15060
rect 4175 14950 4255 15000
rect 4175 14890 4185 14950
rect 4245 14890 4255 14950
rect 4175 14885 4255 14890
rect 4575 15060 4655 15065
rect 4575 15000 4585 15060
rect 4645 15000 4655 15060
rect 4575 14950 4655 15000
rect 4575 14890 4585 14950
rect 4645 14890 4655 14950
rect 4575 14885 4655 14890
rect 4975 15060 5055 15065
rect 4975 15000 4985 15060
rect 5045 15000 5055 15060
rect 4975 14950 5055 15000
rect 4975 14890 4985 14950
rect 5045 14890 5055 14950
rect 4975 14885 5055 14890
rect 5375 15060 5455 15065
rect 5375 15000 5385 15060
rect 5445 15000 5455 15060
rect 5375 14950 5455 15000
rect 5375 14890 5385 14950
rect 5445 14890 5455 14950
rect 5375 14885 5455 14890
rect 5775 15060 5855 15065
rect 5775 15000 5785 15060
rect 5845 15000 5855 15060
rect 5775 14950 5855 15000
rect 5775 14890 5785 14950
rect 5845 14890 5855 14950
rect 5775 14885 5855 14890
rect 6175 15060 6255 15065
rect 6175 15000 6185 15060
rect 6245 15000 6255 15060
rect 6175 14950 6255 15000
rect 6175 14890 6185 14950
rect 6245 14890 6255 14950
rect 6175 14885 6255 14890
rect 6575 15060 6655 15065
rect 6575 15000 6585 15060
rect 6645 15000 6655 15060
rect 6575 14950 6655 15000
rect 6575 14890 6585 14950
rect 6645 14890 6655 14950
rect 6575 14885 6655 14890
rect 6975 15060 7055 15065
rect 6975 15000 6985 15060
rect 7045 15000 7055 15060
rect 6975 14950 7055 15000
rect 6975 14890 6985 14950
rect 7045 14890 7055 14950
rect 6975 14885 7055 14890
rect 7375 15060 7455 15065
rect 7375 15000 7385 15060
rect 7445 15000 7455 15060
rect 7375 14950 7455 15000
rect 7375 14890 7385 14950
rect 7445 14890 7455 14950
rect 7375 14885 7455 14890
rect 7775 15060 7855 15065
rect 7775 15000 7785 15060
rect 7845 15000 7855 15060
rect 7775 14950 7855 15000
rect 7775 14890 7785 14950
rect 7845 14890 7855 14950
rect 7775 14885 7855 14890
rect 8175 15060 8255 15065
rect 8175 15000 8185 15060
rect 8245 15000 8255 15060
rect 8175 14950 8255 15000
rect 8175 14890 8185 14950
rect 8245 14890 8255 14950
rect 8175 14885 8255 14890
rect 8575 15060 8655 15065
rect 8575 15000 8585 15060
rect 8645 15000 8655 15060
rect 8575 14950 8655 15000
rect 8575 14890 8585 14950
rect 8645 14890 8655 14950
rect 8575 14885 8655 14890
rect 8975 15060 9055 15065
rect 8975 15000 8985 15060
rect 9045 15000 9055 15060
rect 8975 14950 9055 15000
rect 8975 14890 8985 14950
rect 9045 14890 9055 14950
rect 8975 14885 9055 14890
rect 9375 15060 9455 15065
rect 9375 15000 9385 15060
rect 9445 15000 9455 15060
rect 9375 14950 9455 15000
rect 9375 14890 9385 14950
rect 9445 14890 9455 14950
rect 9375 14885 9455 14890
rect 9775 15060 9855 15065
rect 9775 15000 9785 15060
rect 9845 15000 9855 15060
rect 9775 14950 9855 15000
rect 9775 14890 9785 14950
rect 9845 14890 9855 14950
rect 9775 14885 9855 14890
rect 10175 15060 10255 15065
rect 10175 15000 10185 15060
rect 10245 15000 10255 15060
rect 10175 14950 10255 15000
rect 10175 14890 10185 14950
rect 10245 14890 10255 14950
rect 10175 14885 10255 14890
rect 10575 15060 10655 15065
rect 10575 15000 10585 15060
rect 10645 15000 10655 15060
rect 10575 14950 10655 15000
rect 10575 14890 10585 14950
rect 10645 14890 10655 14950
rect 10575 14885 10655 14890
rect 10975 15060 11055 15065
rect 10975 15000 10985 15060
rect 11045 15000 11055 15060
rect 10975 14950 11055 15000
rect 10975 14890 10985 14950
rect 11045 14890 11055 14950
rect 10975 14885 11055 14890
rect 11375 15060 11455 15065
rect 11375 15000 11385 15060
rect 11445 15000 11455 15060
rect 11375 14950 11455 15000
rect 11375 14890 11385 14950
rect 11445 14890 11455 14950
rect 11375 14885 11455 14890
rect 11775 15060 11855 15065
rect 11775 15000 11785 15060
rect 11845 15000 11855 15060
rect 11775 14950 11855 15000
rect 11775 14890 11785 14950
rect 11845 14890 11855 14950
rect 11775 14885 11855 14890
rect 12175 15060 12255 15065
rect 12175 15000 12185 15060
rect 12245 15000 12255 15060
rect 12175 14950 12255 15000
rect 12175 14890 12185 14950
rect 12245 14890 12255 14950
rect 12175 14885 12255 14890
rect 12575 15060 12655 15065
rect 12575 15000 12585 15060
rect 12645 15000 12655 15060
rect 12575 14950 12655 15000
rect 12575 14890 12585 14950
rect 12645 14890 12655 14950
rect 12575 14885 12655 14890
rect 12975 15060 13055 15065
rect 12975 15000 12985 15060
rect 13045 15000 13055 15060
rect 12975 14950 13055 15000
rect 12975 14890 12985 14950
rect 13045 14890 13055 14950
rect 12975 14885 13055 14890
rect -215 14695 -155 14885
rect 185 14695 245 14885
rect 585 14695 645 14885
rect 985 14695 1045 14885
rect 1385 14695 1445 14885
rect 1785 14695 1845 14885
rect 2185 14695 2245 14885
rect 2585 14695 2645 14885
rect 2985 14695 3045 14885
rect 3385 14695 3445 14885
rect 3785 14695 3845 14885
rect 4185 14695 4245 14885
rect 4585 14695 4645 14885
rect 4985 14695 5045 14885
rect 5385 14695 5445 14885
rect 5785 14695 5845 14885
rect 6185 14695 6245 14885
rect 6585 14695 6645 14885
rect 6985 14695 7045 14885
rect 7385 14695 7445 14885
rect 7785 14695 7845 14885
rect 8185 14695 8245 14885
rect 8585 14695 8645 14885
rect 8985 14695 9045 14885
rect 9385 14695 9445 14885
rect 9785 14695 9845 14885
rect 10185 14695 10245 14885
rect 10585 14695 10645 14885
rect 10985 14695 11045 14885
rect 11385 14695 11445 14885
rect 11785 14695 11845 14885
rect 12185 14695 12245 14885
rect 12585 14695 12645 14885
rect 12985 14695 13045 14885
rect -225 14690 -145 14695
rect -225 14630 -215 14690
rect -155 14630 -145 14690
rect -225 14580 -145 14630
rect -225 14520 -215 14580
rect -155 14520 -145 14580
rect -225 14515 -145 14520
rect 175 14690 255 14695
rect 175 14630 185 14690
rect 245 14630 255 14690
rect 175 14580 255 14630
rect 175 14520 185 14580
rect 245 14520 255 14580
rect 175 14515 255 14520
rect 575 14690 655 14695
rect 575 14630 585 14690
rect 645 14630 655 14690
rect 575 14580 655 14630
rect 575 14520 585 14580
rect 645 14520 655 14580
rect 575 14515 655 14520
rect 975 14690 1055 14695
rect 975 14630 985 14690
rect 1045 14630 1055 14690
rect 975 14580 1055 14630
rect 975 14520 985 14580
rect 1045 14520 1055 14580
rect 975 14515 1055 14520
rect 1375 14690 1455 14695
rect 1375 14630 1385 14690
rect 1445 14630 1455 14690
rect 1375 14580 1455 14630
rect 1375 14520 1385 14580
rect 1445 14520 1455 14580
rect 1375 14515 1455 14520
rect 1775 14690 1855 14695
rect 1775 14630 1785 14690
rect 1845 14630 1855 14690
rect 1775 14580 1855 14630
rect 1775 14520 1785 14580
rect 1845 14520 1855 14580
rect 1775 14515 1855 14520
rect 2175 14690 2255 14695
rect 2175 14630 2185 14690
rect 2245 14630 2255 14690
rect 2175 14580 2255 14630
rect 2175 14520 2185 14580
rect 2245 14520 2255 14580
rect 2175 14515 2255 14520
rect 2575 14690 2655 14695
rect 2575 14630 2585 14690
rect 2645 14630 2655 14690
rect 2575 14580 2655 14630
rect 2575 14520 2585 14580
rect 2645 14520 2655 14580
rect 2575 14515 2655 14520
rect 2975 14690 3055 14695
rect 2975 14630 2985 14690
rect 3045 14630 3055 14690
rect 2975 14580 3055 14630
rect 2975 14520 2985 14580
rect 3045 14520 3055 14580
rect 2975 14515 3055 14520
rect 3375 14690 3455 14695
rect 3375 14630 3385 14690
rect 3445 14630 3455 14690
rect 3375 14580 3455 14630
rect 3375 14520 3385 14580
rect 3445 14520 3455 14580
rect 3375 14515 3455 14520
rect 3775 14690 3855 14695
rect 3775 14630 3785 14690
rect 3845 14630 3855 14690
rect 3775 14580 3855 14630
rect 3775 14520 3785 14580
rect 3845 14520 3855 14580
rect 3775 14515 3855 14520
rect 4175 14690 4255 14695
rect 4175 14630 4185 14690
rect 4245 14630 4255 14690
rect 4175 14580 4255 14630
rect 4175 14520 4185 14580
rect 4245 14520 4255 14580
rect 4175 14515 4255 14520
rect 4575 14690 4655 14695
rect 4575 14630 4585 14690
rect 4645 14630 4655 14690
rect 4575 14580 4655 14630
rect 4575 14520 4585 14580
rect 4645 14520 4655 14580
rect 4575 14515 4655 14520
rect 4975 14690 5055 14695
rect 4975 14630 4985 14690
rect 5045 14630 5055 14690
rect 4975 14580 5055 14630
rect 4975 14520 4985 14580
rect 5045 14520 5055 14580
rect 4975 14515 5055 14520
rect 5375 14690 5455 14695
rect 5375 14630 5385 14690
rect 5445 14630 5455 14690
rect 5375 14580 5455 14630
rect 5375 14520 5385 14580
rect 5445 14520 5455 14580
rect 5375 14515 5455 14520
rect 5775 14690 5855 14695
rect 5775 14630 5785 14690
rect 5845 14630 5855 14690
rect 5775 14580 5855 14630
rect 5775 14520 5785 14580
rect 5845 14520 5855 14580
rect 5775 14515 5855 14520
rect 6175 14690 6255 14695
rect 6175 14630 6185 14690
rect 6245 14630 6255 14690
rect 6175 14580 6255 14630
rect 6175 14520 6185 14580
rect 6245 14520 6255 14580
rect 6175 14515 6255 14520
rect 6575 14690 6655 14695
rect 6575 14630 6585 14690
rect 6645 14630 6655 14690
rect 6575 14580 6655 14630
rect 6575 14520 6585 14580
rect 6645 14520 6655 14580
rect 6575 14515 6655 14520
rect 6975 14690 7055 14695
rect 6975 14630 6985 14690
rect 7045 14630 7055 14690
rect 6975 14580 7055 14630
rect 6975 14520 6985 14580
rect 7045 14520 7055 14580
rect 6975 14515 7055 14520
rect 7375 14690 7455 14695
rect 7375 14630 7385 14690
rect 7445 14630 7455 14690
rect 7375 14580 7455 14630
rect 7375 14520 7385 14580
rect 7445 14520 7455 14580
rect 7375 14515 7455 14520
rect 7775 14690 7855 14695
rect 7775 14630 7785 14690
rect 7845 14630 7855 14690
rect 7775 14580 7855 14630
rect 7775 14520 7785 14580
rect 7845 14520 7855 14580
rect 7775 14515 7855 14520
rect 8175 14690 8255 14695
rect 8175 14630 8185 14690
rect 8245 14630 8255 14690
rect 8175 14580 8255 14630
rect 8175 14520 8185 14580
rect 8245 14520 8255 14580
rect 8175 14515 8255 14520
rect 8575 14690 8655 14695
rect 8575 14630 8585 14690
rect 8645 14630 8655 14690
rect 8575 14580 8655 14630
rect 8575 14520 8585 14580
rect 8645 14520 8655 14580
rect 8575 14515 8655 14520
rect 8975 14690 9055 14695
rect 8975 14630 8985 14690
rect 9045 14630 9055 14690
rect 8975 14580 9055 14630
rect 8975 14520 8985 14580
rect 9045 14520 9055 14580
rect 8975 14515 9055 14520
rect 9375 14690 9455 14695
rect 9375 14630 9385 14690
rect 9445 14630 9455 14690
rect 9375 14580 9455 14630
rect 9375 14520 9385 14580
rect 9445 14520 9455 14580
rect 9375 14515 9455 14520
rect 9775 14690 9855 14695
rect 9775 14630 9785 14690
rect 9845 14630 9855 14690
rect 9775 14580 9855 14630
rect 9775 14520 9785 14580
rect 9845 14520 9855 14580
rect 9775 14515 9855 14520
rect 10175 14690 10255 14695
rect 10175 14630 10185 14690
rect 10245 14630 10255 14690
rect 10175 14580 10255 14630
rect 10175 14520 10185 14580
rect 10245 14520 10255 14580
rect 10175 14515 10255 14520
rect 10575 14690 10655 14695
rect 10575 14630 10585 14690
rect 10645 14630 10655 14690
rect 10575 14580 10655 14630
rect 10575 14520 10585 14580
rect 10645 14520 10655 14580
rect 10575 14515 10655 14520
rect 10975 14690 11055 14695
rect 10975 14630 10985 14690
rect 11045 14630 11055 14690
rect 10975 14580 11055 14630
rect 10975 14520 10985 14580
rect 11045 14520 11055 14580
rect 10975 14515 11055 14520
rect 11375 14690 11455 14695
rect 11375 14630 11385 14690
rect 11445 14630 11455 14690
rect 11375 14580 11455 14630
rect 11375 14520 11385 14580
rect 11445 14520 11455 14580
rect 11375 14515 11455 14520
rect 11775 14690 11855 14695
rect 11775 14630 11785 14690
rect 11845 14630 11855 14690
rect 11775 14580 11855 14630
rect 11775 14520 11785 14580
rect 11845 14520 11855 14580
rect 11775 14515 11855 14520
rect 12175 14690 12255 14695
rect 12175 14630 12185 14690
rect 12245 14630 12255 14690
rect 12175 14580 12255 14630
rect 12175 14520 12185 14580
rect 12245 14520 12255 14580
rect 12175 14515 12255 14520
rect 12575 14690 12655 14695
rect 12575 14630 12585 14690
rect 12645 14630 12655 14690
rect 12575 14580 12655 14630
rect 12575 14520 12585 14580
rect 12645 14520 12655 14580
rect 12575 14515 12655 14520
rect 12975 14690 13055 14695
rect 12975 14630 12985 14690
rect 13045 14630 13055 14690
rect 12975 14580 13055 14630
rect 12975 14520 12985 14580
rect 13045 14520 13055 14580
rect 12975 14515 13055 14520
rect -215 14325 -155 14515
rect 185 14325 245 14515
rect 585 14325 645 14515
rect 985 14325 1045 14515
rect 1385 14325 1445 14515
rect 1785 14325 1845 14515
rect 2185 14325 2245 14515
rect 2585 14325 2645 14515
rect 2985 14325 3045 14515
rect 3385 14325 3445 14515
rect 3785 14325 3845 14515
rect 4185 14325 4245 14515
rect 4585 14325 4645 14515
rect 4985 14325 5045 14515
rect 5385 14325 5445 14515
rect 5785 14325 5845 14515
rect 6185 14325 6245 14515
rect 6585 14325 6645 14515
rect 6985 14325 7045 14515
rect 7385 14325 7445 14515
rect 7785 14325 7845 14515
rect 8185 14325 8245 14515
rect 8585 14325 8645 14515
rect 8985 14325 9045 14515
rect 9385 14325 9445 14515
rect 9785 14325 9845 14515
rect 10185 14325 10245 14515
rect 10585 14325 10645 14515
rect 10985 14325 11045 14515
rect 11385 14325 11445 14515
rect 11785 14325 11845 14515
rect 12185 14325 12245 14515
rect 12585 14325 12645 14515
rect 12985 14325 13045 14515
rect -225 14320 -145 14325
rect -225 14260 -215 14320
rect -155 14260 -145 14320
rect -225 14210 -145 14260
rect -225 14150 -215 14210
rect -155 14150 -145 14210
rect -225 14145 -145 14150
rect 175 14320 255 14325
rect 175 14260 185 14320
rect 245 14260 255 14320
rect 175 14210 255 14260
rect 175 14150 185 14210
rect 245 14150 255 14210
rect 175 14145 255 14150
rect 575 14320 655 14325
rect 575 14260 585 14320
rect 645 14260 655 14320
rect 575 14210 655 14260
rect 575 14150 585 14210
rect 645 14150 655 14210
rect 575 14145 655 14150
rect 975 14320 1055 14325
rect 975 14260 985 14320
rect 1045 14260 1055 14320
rect 975 14210 1055 14260
rect 975 14150 985 14210
rect 1045 14150 1055 14210
rect 975 14145 1055 14150
rect 1375 14320 1455 14325
rect 1375 14260 1385 14320
rect 1445 14260 1455 14320
rect 1375 14210 1455 14260
rect 1375 14150 1385 14210
rect 1445 14150 1455 14210
rect 1375 14145 1455 14150
rect 1775 14320 1855 14325
rect 1775 14260 1785 14320
rect 1845 14260 1855 14320
rect 1775 14210 1855 14260
rect 1775 14150 1785 14210
rect 1845 14150 1855 14210
rect 1775 14145 1855 14150
rect 2175 14320 2255 14325
rect 2175 14260 2185 14320
rect 2245 14260 2255 14320
rect 2175 14210 2255 14260
rect 2175 14150 2185 14210
rect 2245 14150 2255 14210
rect 2175 14145 2255 14150
rect 2575 14320 2655 14325
rect 2575 14260 2585 14320
rect 2645 14260 2655 14320
rect 2575 14210 2655 14260
rect 2575 14150 2585 14210
rect 2645 14150 2655 14210
rect 2575 14145 2655 14150
rect 2975 14320 3055 14325
rect 2975 14260 2985 14320
rect 3045 14260 3055 14320
rect 2975 14210 3055 14260
rect 2975 14150 2985 14210
rect 3045 14150 3055 14210
rect 2975 14145 3055 14150
rect 3375 14320 3455 14325
rect 3375 14260 3385 14320
rect 3445 14260 3455 14320
rect 3375 14210 3455 14260
rect 3375 14150 3385 14210
rect 3445 14150 3455 14210
rect 3375 14145 3455 14150
rect 3775 14320 3855 14325
rect 3775 14260 3785 14320
rect 3845 14260 3855 14320
rect 3775 14210 3855 14260
rect 3775 14150 3785 14210
rect 3845 14150 3855 14210
rect 3775 14145 3855 14150
rect 4175 14320 4255 14325
rect 4175 14260 4185 14320
rect 4245 14260 4255 14320
rect 4175 14210 4255 14260
rect 4175 14150 4185 14210
rect 4245 14150 4255 14210
rect 4175 14145 4255 14150
rect 4575 14320 4655 14325
rect 4575 14260 4585 14320
rect 4645 14260 4655 14320
rect 4575 14210 4655 14260
rect 4575 14150 4585 14210
rect 4645 14150 4655 14210
rect 4575 14145 4655 14150
rect 4975 14320 5055 14325
rect 4975 14260 4985 14320
rect 5045 14260 5055 14320
rect 4975 14210 5055 14260
rect 4975 14150 4985 14210
rect 5045 14150 5055 14210
rect 4975 14145 5055 14150
rect 5375 14320 5455 14325
rect 5375 14260 5385 14320
rect 5445 14260 5455 14320
rect 5375 14210 5455 14260
rect 5375 14150 5385 14210
rect 5445 14150 5455 14210
rect 5375 14145 5455 14150
rect 5775 14320 5855 14325
rect 5775 14260 5785 14320
rect 5845 14260 5855 14320
rect 5775 14210 5855 14260
rect 5775 14150 5785 14210
rect 5845 14150 5855 14210
rect 5775 14145 5855 14150
rect 6175 14320 6255 14325
rect 6175 14260 6185 14320
rect 6245 14260 6255 14320
rect 6175 14210 6255 14260
rect 6175 14150 6185 14210
rect 6245 14150 6255 14210
rect 6175 14145 6255 14150
rect 6575 14320 6655 14325
rect 6575 14260 6585 14320
rect 6645 14260 6655 14320
rect 6575 14210 6655 14260
rect 6575 14150 6585 14210
rect 6645 14150 6655 14210
rect 6575 14145 6655 14150
rect 6975 14320 7055 14325
rect 6975 14260 6985 14320
rect 7045 14260 7055 14320
rect 6975 14210 7055 14260
rect 6975 14150 6985 14210
rect 7045 14150 7055 14210
rect 6975 14145 7055 14150
rect 7375 14320 7455 14325
rect 7375 14260 7385 14320
rect 7445 14260 7455 14320
rect 7375 14210 7455 14260
rect 7375 14150 7385 14210
rect 7445 14150 7455 14210
rect 7375 14145 7455 14150
rect 7775 14320 7855 14325
rect 7775 14260 7785 14320
rect 7845 14260 7855 14320
rect 7775 14210 7855 14260
rect 7775 14150 7785 14210
rect 7845 14150 7855 14210
rect 7775 14145 7855 14150
rect 8175 14320 8255 14325
rect 8175 14260 8185 14320
rect 8245 14260 8255 14320
rect 8175 14210 8255 14260
rect 8175 14150 8185 14210
rect 8245 14150 8255 14210
rect 8175 14145 8255 14150
rect 8575 14320 8655 14325
rect 8575 14260 8585 14320
rect 8645 14260 8655 14320
rect 8575 14210 8655 14260
rect 8575 14150 8585 14210
rect 8645 14150 8655 14210
rect 8575 14145 8655 14150
rect 8975 14320 9055 14325
rect 8975 14260 8985 14320
rect 9045 14260 9055 14320
rect 8975 14210 9055 14260
rect 8975 14150 8985 14210
rect 9045 14150 9055 14210
rect 8975 14145 9055 14150
rect 9375 14320 9455 14325
rect 9375 14260 9385 14320
rect 9445 14260 9455 14320
rect 9375 14210 9455 14260
rect 9375 14150 9385 14210
rect 9445 14150 9455 14210
rect 9375 14145 9455 14150
rect 9775 14320 9855 14325
rect 9775 14260 9785 14320
rect 9845 14260 9855 14320
rect 9775 14210 9855 14260
rect 9775 14150 9785 14210
rect 9845 14150 9855 14210
rect 9775 14145 9855 14150
rect 10175 14320 10255 14325
rect 10175 14260 10185 14320
rect 10245 14260 10255 14320
rect 10175 14210 10255 14260
rect 10175 14150 10185 14210
rect 10245 14150 10255 14210
rect 10175 14145 10255 14150
rect 10575 14320 10655 14325
rect 10575 14260 10585 14320
rect 10645 14260 10655 14320
rect 10575 14210 10655 14260
rect 10575 14150 10585 14210
rect 10645 14150 10655 14210
rect 10575 14145 10655 14150
rect 10975 14320 11055 14325
rect 10975 14260 10985 14320
rect 11045 14260 11055 14320
rect 10975 14210 11055 14260
rect 10975 14150 10985 14210
rect 11045 14150 11055 14210
rect 10975 14145 11055 14150
rect 11375 14320 11455 14325
rect 11375 14260 11385 14320
rect 11445 14260 11455 14320
rect 11375 14210 11455 14260
rect 11375 14150 11385 14210
rect 11445 14150 11455 14210
rect 11375 14145 11455 14150
rect 11775 14320 11855 14325
rect 11775 14260 11785 14320
rect 11845 14260 11855 14320
rect 11775 14210 11855 14260
rect 11775 14150 11785 14210
rect 11845 14150 11855 14210
rect 11775 14145 11855 14150
rect 12175 14320 12255 14325
rect 12175 14260 12185 14320
rect 12245 14260 12255 14320
rect 12175 14210 12255 14260
rect 12175 14150 12185 14210
rect 12245 14150 12255 14210
rect 12175 14145 12255 14150
rect 12575 14320 12655 14325
rect 12575 14260 12585 14320
rect 12645 14260 12655 14320
rect 12575 14210 12655 14260
rect 12575 14150 12585 14210
rect 12645 14150 12655 14210
rect 12575 14145 12655 14150
rect 12975 14320 13055 14325
rect 12975 14260 12985 14320
rect 13045 14260 13055 14320
rect 12975 14210 13055 14260
rect 12975 14150 12985 14210
rect 13045 14150 13055 14210
rect 12975 14145 13055 14150
rect -215 13955 -155 14145
rect 185 13955 245 14145
rect 585 13955 645 14145
rect 985 13955 1045 14145
rect 1385 13955 1445 14145
rect 1785 13955 1845 14145
rect 2185 13955 2245 14145
rect 2585 13955 2645 14145
rect 2985 13955 3045 14145
rect 3385 13955 3445 14145
rect 3785 13955 3845 14145
rect 4185 13955 4245 14145
rect 4585 13955 4645 14145
rect 4985 13955 5045 14145
rect 5385 13955 5445 14145
rect 5785 13955 5845 14145
rect 6185 13955 6245 14145
rect 6585 13955 6645 14145
rect 6985 13955 7045 14145
rect 7385 13955 7445 14145
rect 7785 13955 7845 14145
rect 8185 13955 8245 14145
rect 8585 13955 8645 14145
rect 8985 13955 9045 14145
rect 9385 13955 9445 14145
rect 9785 13955 9845 14145
rect 10185 13955 10245 14145
rect 10585 13955 10645 14145
rect 10985 13955 11045 14145
rect 11385 13955 11445 14145
rect 11785 13955 11845 14145
rect 12185 13955 12245 14145
rect 12585 13955 12645 14145
rect 12985 13955 13045 14145
rect -225 13950 -145 13955
rect -225 13890 -215 13950
rect -155 13890 -145 13950
rect -225 13840 -145 13890
rect -225 13780 -215 13840
rect -155 13780 -145 13840
rect -225 13775 -145 13780
rect 175 13950 255 13955
rect 175 13890 185 13950
rect 245 13890 255 13950
rect 175 13840 255 13890
rect 175 13780 185 13840
rect 245 13780 255 13840
rect 175 13775 255 13780
rect 575 13950 655 13955
rect 575 13890 585 13950
rect 645 13890 655 13950
rect 575 13840 655 13890
rect 575 13780 585 13840
rect 645 13780 655 13840
rect 575 13775 655 13780
rect 975 13950 1055 13955
rect 975 13890 985 13950
rect 1045 13890 1055 13950
rect 975 13840 1055 13890
rect 975 13780 985 13840
rect 1045 13780 1055 13840
rect 975 13775 1055 13780
rect 1375 13950 1455 13955
rect 1375 13890 1385 13950
rect 1445 13890 1455 13950
rect 1375 13840 1455 13890
rect 1375 13780 1385 13840
rect 1445 13780 1455 13840
rect 1375 13775 1455 13780
rect 1775 13950 1855 13955
rect 1775 13890 1785 13950
rect 1845 13890 1855 13950
rect 1775 13840 1855 13890
rect 1775 13780 1785 13840
rect 1845 13780 1855 13840
rect 1775 13775 1855 13780
rect 2175 13950 2255 13955
rect 2175 13890 2185 13950
rect 2245 13890 2255 13950
rect 2175 13840 2255 13890
rect 2175 13780 2185 13840
rect 2245 13780 2255 13840
rect 2175 13775 2255 13780
rect 2575 13950 2655 13955
rect 2575 13890 2585 13950
rect 2645 13890 2655 13950
rect 2575 13840 2655 13890
rect 2575 13780 2585 13840
rect 2645 13780 2655 13840
rect 2575 13775 2655 13780
rect 2975 13950 3055 13955
rect 2975 13890 2985 13950
rect 3045 13890 3055 13950
rect 2975 13840 3055 13890
rect 2975 13780 2985 13840
rect 3045 13780 3055 13840
rect 2975 13775 3055 13780
rect 3375 13950 3455 13955
rect 3375 13890 3385 13950
rect 3445 13890 3455 13950
rect 3375 13840 3455 13890
rect 3375 13780 3385 13840
rect 3445 13780 3455 13840
rect 3375 13775 3455 13780
rect 3775 13950 3855 13955
rect 3775 13890 3785 13950
rect 3845 13890 3855 13950
rect 3775 13840 3855 13890
rect 3775 13780 3785 13840
rect 3845 13780 3855 13840
rect 3775 13775 3855 13780
rect 4175 13950 4255 13955
rect 4175 13890 4185 13950
rect 4245 13890 4255 13950
rect 4175 13840 4255 13890
rect 4175 13780 4185 13840
rect 4245 13780 4255 13840
rect 4175 13775 4255 13780
rect 4575 13950 4655 13955
rect 4575 13890 4585 13950
rect 4645 13890 4655 13950
rect 4575 13840 4655 13890
rect 4575 13780 4585 13840
rect 4645 13780 4655 13840
rect 4575 13775 4655 13780
rect 4975 13950 5055 13955
rect 4975 13890 4985 13950
rect 5045 13890 5055 13950
rect 4975 13840 5055 13890
rect 4975 13780 4985 13840
rect 5045 13780 5055 13840
rect 4975 13775 5055 13780
rect 5375 13950 5455 13955
rect 5375 13890 5385 13950
rect 5445 13890 5455 13950
rect 5375 13840 5455 13890
rect 5375 13780 5385 13840
rect 5445 13780 5455 13840
rect 5375 13775 5455 13780
rect 5775 13950 5855 13955
rect 5775 13890 5785 13950
rect 5845 13890 5855 13950
rect 5775 13840 5855 13890
rect 5775 13780 5785 13840
rect 5845 13780 5855 13840
rect 5775 13775 5855 13780
rect 6175 13950 6255 13955
rect 6175 13890 6185 13950
rect 6245 13890 6255 13950
rect 6175 13840 6255 13890
rect 6175 13780 6185 13840
rect 6245 13780 6255 13840
rect 6175 13775 6255 13780
rect 6575 13950 6655 13955
rect 6575 13890 6585 13950
rect 6645 13890 6655 13950
rect 6575 13840 6655 13890
rect 6575 13780 6585 13840
rect 6645 13780 6655 13840
rect 6575 13775 6655 13780
rect 6975 13950 7055 13955
rect 6975 13890 6985 13950
rect 7045 13890 7055 13950
rect 6975 13840 7055 13890
rect 6975 13780 6985 13840
rect 7045 13780 7055 13840
rect 6975 13775 7055 13780
rect 7375 13950 7455 13955
rect 7375 13890 7385 13950
rect 7445 13890 7455 13950
rect 7375 13840 7455 13890
rect 7375 13780 7385 13840
rect 7445 13780 7455 13840
rect 7375 13775 7455 13780
rect 7775 13950 7855 13955
rect 7775 13890 7785 13950
rect 7845 13890 7855 13950
rect 7775 13840 7855 13890
rect 7775 13780 7785 13840
rect 7845 13780 7855 13840
rect 7775 13775 7855 13780
rect 8175 13950 8255 13955
rect 8175 13890 8185 13950
rect 8245 13890 8255 13950
rect 8175 13840 8255 13890
rect 8175 13780 8185 13840
rect 8245 13780 8255 13840
rect 8175 13775 8255 13780
rect 8575 13950 8655 13955
rect 8575 13890 8585 13950
rect 8645 13890 8655 13950
rect 8575 13840 8655 13890
rect 8575 13780 8585 13840
rect 8645 13780 8655 13840
rect 8575 13775 8655 13780
rect 8975 13950 9055 13955
rect 8975 13890 8985 13950
rect 9045 13890 9055 13950
rect 8975 13840 9055 13890
rect 8975 13780 8985 13840
rect 9045 13780 9055 13840
rect 8975 13775 9055 13780
rect 9375 13950 9455 13955
rect 9375 13890 9385 13950
rect 9445 13890 9455 13950
rect 9375 13840 9455 13890
rect 9375 13780 9385 13840
rect 9445 13780 9455 13840
rect 9375 13775 9455 13780
rect 9775 13950 9855 13955
rect 9775 13890 9785 13950
rect 9845 13890 9855 13950
rect 9775 13840 9855 13890
rect 9775 13780 9785 13840
rect 9845 13780 9855 13840
rect 9775 13775 9855 13780
rect 10175 13950 10255 13955
rect 10175 13890 10185 13950
rect 10245 13890 10255 13950
rect 10175 13840 10255 13890
rect 10175 13780 10185 13840
rect 10245 13780 10255 13840
rect 10175 13775 10255 13780
rect 10575 13950 10655 13955
rect 10575 13890 10585 13950
rect 10645 13890 10655 13950
rect 10575 13840 10655 13890
rect 10575 13780 10585 13840
rect 10645 13780 10655 13840
rect 10575 13775 10655 13780
rect 10975 13950 11055 13955
rect 10975 13890 10985 13950
rect 11045 13890 11055 13950
rect 10975 13840 11055 13890
rect 10975 13780 10985 13840
rect 11045 13780 11055 13840
rect 10975 13775 11055 13780
rect 11375 13950 11455 13955
rect 11375 13890 11385 13950
rect 11445 13890 11455 13950
rect 11375 13840 11455 13890
rect 11375 13780 11385 13840
rect 11445 13780 11455 13840
rect 11375 13775 11455 13780
rect 11775 13950 11855 13955
rect 11775 13890 11785 13950
rect 11845 13890 11855 13950
rect 11775 13840 11855 13890
rect 11775 13780 11785 13840
rect 11845 13780 11855 13840
rect 11775 13775 11855 13780
rect 12175 13950 12255 13955
rect 12175 13890 12185 13950
rect 12245 13890 12255 13950
rect 12175 13840 12255 13890
rect 12175 13780 12185 13840
rect 12245 13780 12255 13840
rect 12175 13775 12255 13780
rect 12575 13950 12655 13955
rect 12575 13890 12585 13950
rect 12645 13890 12655 13950
rect 12575 13840 12655 13890
rect 12575 13780 12585 13840
rect 12645 13780 12655 13840
rect 12575 13775 12655 13780
rect 12975 13950 13055 13955
rect 12975 13890 12985 13950
rect 13045 13890 13055 13950
rect 12975 13840 13055 13890
rect 12975 13780 12985 13840
rect 13045 13780 13055 13840
rect 12975 13775 13055 13780
rect -215 13585 -155 13775
rect 185 13585 245 13775
rect 585 13585 645 13775
rect 985 13585 1045 13775
rect 1385 13585 1445 13775
rect 1785 13585 1845 13775
rect 2185 13585 2245 13775
rect 2585 13585 2645 13775
rect 2985 13585 3045 13775
rect 3385 13585 3445 13775
rect 3785 13585 3845 13775
rect 4185 13585 4245 13775
rect 4585 13585 4645 13775
rect 4985 13585 5045 13775
rect 5385 13585 5445 13775
rect 5785 13585 5845 13775
rect 6185 13585 6245 13775
rect 6585 13585 6645 13775
rect 6985 13585 7045 13775
rect 7385 13585 7445 13775
rect 7785 13585 7845 13775
rect 8185 13585 8245 13775
rect 8585 13585 8645 13775
rect 8985 13585 9045 13775
rect 9385 13585 9445 13775
rect 9785 13585 9845 13775
rect 10185 13585 10245 13775
rect 10585 13585 10645 13775
rect 10985 13585 11045 13775
rect 11385 13585 11445 13775
rect 11785 13585 11845 13775
rect 12185 13585 12245 13775
rect 12585 13585 12645 13775
rect 12985 13585 13045 13775
rect -225 13580 -145 13585
rect -225 13520 -215 13580
rect -155 13520 -145 13580
rect -225 13470 -145 13520
rect -225 13410 -215 13470
rect -155 13410 -145 13470
rect -225 13405 -145 13410
rect 175 13580 255 13585
rect 175 13520 185 13580
rect 245 13520 255 13580
rect 175 13470 255 13520
rect 175 13410 185 13470
rect 245 13410 255 13470
rect 175 13405 255 13410
rect 575 13580 655 13585
rect 575 13520 585 13580
rect 645 13520 655 13580
rect 575 13470 655 13520
rect 575 13410 585 13470
rect 645 13410 655 13470
rect 575 13405 655 13410
rect 975 13580 1055 13585
rect 975 13520 985 13580
rect 1045 13520 1055 13580
rect 975 13470 1055 13520
rect 975 13410 985 13470
rect 1045 13410 1055 13470
rect 975 13405 1055 13410
rect 1375 13580 1455 13585
rect 1375 13520 1385 13580
rect 1445 13520 1455 13580
rect 1375 13470 1455 13520
rect 1375 13410 1385 13470
rect 1445 13410 1455 13470
rect 1375 13405 1455 13410
rect 1775 13580 1855 13585
rect 1775 13520 1785 13580
rect 1845 13520 1855 13580
rect 1775 13470 1855 13520
rect 1775 13410 1785 13470
rect 1845 13410 1855 13470
rect 1775 13405 1855 13410
rect 2175 13580 2255 13585
rect 2175 13520 2185 13580
rect 2245 13520 2255 13580
rect 2175 13470 2255 13520
rect 2175 13410 2185 13470
rect 2245 13410 2255 13470
rect 2175 13405 2255 13410
rect 2575 13580 2655 13585
rect 2575 13520 2585 13580
rect 2645 13520 2655 13580
rect 2575 13470 2655 13520
rect 2575 13410 2585 13470
rect 2645 13410 2655 13470
rect 2575 13405 2655 13410
rect 2975 13580 3055 13585
rect 2975 13520 2985 13580
rect 3045 13520 3055 13580
rect 2975 13470 3055 13520
rect 2975 13410 2985 13470
rect 3045 13410 3055 13470
rect 2975 13405 3055 13410
rect 3375 13580 3455 13585
rect 3375 13520 3385 13580
rect 3445 13520 3455 13580
rect 3375 13470 3455 13520
rect 3375 13410 3385 13470
rect 3445 13410 3455 13470
rect 3375 13405 3455 13410
rect 3775 13580 3855 13585
rect 3775 13520 3785 13580
rect 3845 13520 3855 13580
rect 3775 13470 3855 13520
rect 3775 13410 3785 13470
rect 3845 13410 3855 13470
rect 3775 13405 3855 13410
rect 4175 13580 4255 13585
rect 4175 13520 4185 13580
rect 4245 13520 4255 13580
rect 4175 13470 4255 13520
rect 4175 13410 4185 13470
rect 4245 13410 4255 13470
rect 4175 13405 4255 13410
rect 4575 13580 4655 13585
rect 4575 13520 4585 13580
rect 4645 13520 4655 13580
rect 4575 13470 4655 13520
rect 4575 13410 4585 13470
rect 4645 13410 4655 13470
rect 4575 13405 4655 13410
rect 4975 13580 5055 13585
rect 4975 13520 4985 13580
rect 5045 13520 5055 13580
rect 4975 13470 5055 13520
rect 4975 13410 4985 13470
rect 5045 13410 5055 13470
rect 4975 13405 5055 13410
rect 5375 13580 5455 13585
rect 5375 13520 5385 13580
rect 5445 13520 5455 13580
rect 5375 13470 5455 13520
rect 5375 13410 5385 13470
rect 5445 13410 5455 13470
rect 5375 13405 5455 13410
rect 5775 13580 5855 13585
rect 5775 13520 5785 13580
rect 5845 13520 5855 13580
rect 5775 13470 5855 13520
rect 5775 13410 5785 13470
rect 5845 13410 5855 13470
rect 5775 13405 5855 13410
rect 6175 13580 6255 13585
rect 6175 13520 6185 13580
rect 6245 13520 6255 13580
rect 6175 13470 6255 13520
rect 6175 13410 6185 13470
rect 6245 13410 6255 13470
rect 6175 13405 6255 13410
rect 6575 13580 6655 13585
rect 6575 13520 6585 13580
rect 6645 13520 6655 13580
rect 6575 13470 6655 13520
rect 6575 13410 6585 13470
rect 6645 13410 6655 13470
rect 6575 13405 6655 13410
rect 6975 13580 7055 13585
rect 6975 13520 6985 13580
rect 7045 13520 7055 13580
rect 6975 13470 7055 13520
rect 6975 13410 6985 13470
rect 7045 13410 7055 13470
rect 6975 13405 7055 13410
rect 7375 13580 7455 13585
rect 7375 13520 7385 13580
rect 7445 13520 7455 13580
rect 7375 13470 7455 13520
rect 7375 13410 7385 13470
rect 7445 13410 7455 13470
rect 7375 13405 7455 13410
rect 7775 13580 7855 13585
rect 7775 13520 7785 13580
rect 7845 13520 7855 13580
rect 7775 13470 7855 13520
rect 7775 13410 7785 13470
rect 7845 13410 7855 13470
rect 7775 13405 7855 13410
rect 8175 13580 8255 13585
rect 8175 13520 8185 13580
rect 8245 13520 8255 13580
rect 8175 13470 8255 13520
rect 8175 13410 8185 13470
rect 8245 13410 8255 13470
rect 8175 13405 8255 13410
rect 8575 13580 8655 13585
rect 8575 13520 8585 13580
rect 8645 13520 8655 13580
rect 8575 13470 8655 13520
rect 8575 13410 8585 13470
rect 8645 13410 8655 13470
rect 8575 13405 8655 13410
rect 8975 13580 9055 13585
rect 8975 13520 8985 13580
rect 9045 13520 9055 13580
rect 8975 13470 9055 13520
rect 8975 13410 8985 13470
rect 9045 13410 9055 13470
rect 8975 13405 9055 13410
rect 9375 13580 9455 13585
rect 9375 13520 9385 13580
rect 9445 13520 9455 13580
rect 9375 13470 9455 13520
rect 9375 13410 9385 13470
rect 9445 13410 9455 13470
rect 9375 13405 9455 13410
rect 9775 13580 9855 13585
rect 9775 13520 9785 13580
rect 9845 13520 9855 13580
rect 9775 13470 9855 13520
rect 9775 13410 9785 13470
rect 9845 13410 9855 13470
rect 9775 13405 9855 13410
rect 10175 13580 10255 13585
rect 10175 13520 10185 13580
rect 10245 13520 10255 13580
rect 10175 13470 10255 13520
rect 10175 13410 10185 13470
rect 10245 13410 10255 13470
rect 10175 13405 10255 13410
rect 10575 13580 10655 13585
rect 10575 13520 10585 13580
rect 10645 13520 10655 13580
rect 10575 13470 10655 13520
rect 10575 13410 10585 13470
rect 10645 13410 10655 13470
rect 10575 13405 10655 13410
rect 10975 13580 11055 13585
rect 10975 13520 10985 13580
rect 11045 13520 11055 13580
rect 10975 13470 11055 13520
rect 10975 13410 10985 13470
rect 11045 13410 11055 13470
rect 10975 13405 11055 13410
rect 11375 13580 11455 13585
rect 11375 13520 11385 13580
rect 11445 13520 11455 13580
rect 11375 13470 11455 13520
rect 11375 13410 11385 13470
rect 11445 13410 11455 13470
rect 11375 13405 11455 13410
rect 11775 13580 11855 13585
rect 11775 13520 11785 13580
rect 11845 13520 11855 13580
rect 11775 13470 11855 13520
rect 11775 13410 11785 13470
rect 11845 13410 11855 13470
rect 11775 13405 11855 13410
rect 12175 13580 12255 13585
rect 12175 13520 12185 13580
rect 12245 13520 12255 13580
rect 12175 13470 12255 13520
rect 12175 13410 12185 13470
rect 12245 13410 12255 13470
rect 12175 13405 12255 13410
rect 12575 13580 12655 13585
rect 12575 13520 12585 13580
rect 12645 13520 12655 13580
rect 12575 13470 12655 13520
rect 12575 13410 12585 13470
rect 12645 13410 12655 13470
rect 12575 13405 12655 13410
rect 12975 13580 13055 13585
rect 12975 13520 12985 13580
rect 13045 13520 13055 13580
rect 12975 13470 13055 13520
rect 12975 13410 12985 13470
rect 13045 13410 13055 13470
rect 12975 13405 13055 13410
rect -215 13215 -155 13405
rect 185 13215 245 13405
rect 585 13215 645 13405
rect 985 13215 1045 13405
rect 1385 13215 1445 13405
rect 1785 13215 1845 13405
rect 2185 13215 2245 13405
rect 2585 13215 2645 13405
rect 2985 13215 3045 13405
rect 3385 13215 3445 13405
rect 3785 13215 3845 13405
rect 4185 13215 4245 13405
rect 4585 13215 4645 13405
rect 4985 13215 5045 13405
rect 5385 13215 5445 13405
rect 5785 13215 5845 13405
rect 6185 13215 6245 13405
rect 6585 13215 6645 13405
rect 6985 13215 7045 13405
rect 7385 13215 7445 13405
rect 7785 13215 7845 13405
rect 8185 13215 8245 13405
rect 8585 13215 8645 13405
rect 8985 13215 9045 13405
rect 9385 13215 9445 13405
rect 9785 13215 9845 13405
rect 10185 13215 10245 13405
rect 10585 13215 10645 13405
rect 10985 13215 11045 13405
rect 11385 13215 11445 13405
rect 11785 13215 11845 13405
rect 12185 13215 12245 13405
rect 12585 13215 12645 13405
rect 12985 13215 13045 13405
rect -225 13210 -145 13215
rect -225 13150 -215 13210
rect -155 13150 -145 13210
rect -225 13100 -145 13150
rect -225 13040 -215 13100
rect -155 13040 -145 13100
rect -225 13035 -145 13040
rect 175 13210 255 13215
rect 175 13150 185 13210
rect 245 13150 255 13210
rect 175 13100 255 13150
rect 175 13040 185 13100
rect 245 13040 255 13100
rect 175 13035 255 13040
rect 575 13210 655 13215
rect 575 13150 585 13210
rect 645 13150 655 13210
rect 575 13100 655 13150
rect 575 13040 585 13100
rect 645 13040 655 13100
rect 575 13035 655 13040
rect 975 13210 1055 13215
rect 975 13150 985 13210
rect 1045 13150 1055 13210
rect 975 13100 1055 13150
rect 975 13040 985 13100
rect 1045 13040 1055 13100
rect 975 13035 1055 13040
rect 1375 13210 1455 13215
rect 1375 13150 1385 13210
rect 1445 13150 1455 13210
rect 1375 13100 1455 13150
rect 1375 13040 1385 13100
rect 1445 13040 1455 13100
rect 1375 13035 1455 13040
rect 1775 13210 1855 13215
rect 1775 13150 1785 13210
rect 1845 13150 1855 13210
rect 1775 13100 1855 13150
rect 1775 13040 1785 13100
rect 1845 13040 1855 13100
rect 1775 13035 1855 13040
rect 2175 13210 2255 13215
rect 2175 13150 2185 13210
rect 2245 13150 2255 13210
rect 2175 13100 2255 13150
rect 2175 13040 2185 13100
rect 2245 13040 2255 13100
rect 2175 13035 2255 13040
rect 2575 13210 2655 13215
rect 2575 13150 2585 13210
rect 2645 13150 2655 13210
rect 2575 13100 2655 13150
rect 2575 13040 2585 13100
rect 2645 13040 2655 13100
rect 2575 13035 2655 13040
rect 2975 13210 3055 13215
rect 2975 13150 2985 13210
rect 3045 13150 3055 13210
rect 2975 13100 3055 13150
rect 2975 13040 2985 13100
rect 3045 13040 3055 13100
rect 2975 13035 3055 13040
rect 3375 13210 3455 13215
rect 3375 13150 3385 13210
rect 3445 13150 3455 13210
rect 3375 13100 3455 13150
rect 3375 13040 3385 13100
rect 3445 13040 3455 13100
rect 3375 13035 3455 13040
rect 3775 13210 3855 13215
rect 3775 13150 3785 13210
rect 3845 13150 3855 13210
rect 3775 13100 3855 13150
rect 3775 13040 3785 13100
rect 3845 13040 3855 13100
rect 3775 13035 3855 13040
rect 4175 13210 4255 13215
rect 4175 13150 4185 13210
rect 4245 13150 4255 13210
rect 4175 13100 4255 13150
rect 4175 13040 4185 13100
rect 4245 13040 4255 13100
rect 4175 13035 4255 13040
rect 4575 13210 4655 13215
rect 4575 13150 4585 13210
rect 4645 13150 4655 13210
rect 4575 13100 4655 13150
rect 4575 13040 4585 13100
rect 4645 13040 4655 13100
rect 4575 13035 4655 13040
rect 4975 13210 5055 13215
rect 4975 13150 4985 13210
rect 5045 13150 5055 13210
rect 4975 13100 5055 13150
rect 4975 13040 4985 13100
rect 5045 13040 5055 13100
rect 4975 13035 5055 13040
rect 5375 13210 5455 13215
rect 5375 13150 5385 13210
rect 5445 13150 5455 13210
rect 5375 13100 5455 13150
rect 5375 13040 5385 13100
rect 5445 13040 5455 13100
rect 5375 13035 5455 13040
rect 5775 13210 5855 13215
rect 5775 13150 5785 13210
rect 5845 13150 5855 13210
rect 5775 13100 5855 13150
rect 5775 13040 5785 13100
rect 5845 13040 5855 13100
rect 5775 13035 5855 13040
rect 6175 13210 6255 13215
rect 6175 13150 6185 13210
rect 6245 13150 6255 13210
rect 6175 13100 6255 13150
rect 6175 13040 6185 13100
rect 6245 13040 6255 13100
rect 6175 13035 6255 13040
rect 6575 13210 6655 13215
rect 6575 13150 6585 13210
rect 6645 13150 6655 13210
rect 6575 13100 6655 13150
rect 6575 13040 6585 13100
rect 6645 13040 6655 13100
rect 6575 13035 6655 13040
rect 6975 13210 7055 13215
rect 6975 13150 6985 13210
rect 7045 13150 7055 13210
rect 6975 13100 7055 13150
rect 6975 13040 6985 13100
rect 7045 13040 7055 13100
rect 6975 13035 7055 13040
rect 7375 13210 7455 13215
rect 7375 13150 7385 13210
rect 7445 13150 7455 13210
rect 7375 13100 7455 13150
rect 7375 13040 7385 13100
rect 7445 13040 7455 13100
rect 7375 13035 7455 13040
rect 7775 13210 7855 13215
rect 7775 13150 7785 13210
rect 7845 13150 7855 13210
rect 7775 13100 7855 13150
rect 7775 13040 7785 13100
rect 7845 13040 7855 13100
rect 7775 13035 7855 13040
rect 8175 13210 8255 13215
rect 8175 13150 8185 13210
rect 8245 13150 8255 13210
rect 8175 13100 8255 13150
rect 8175 13040 8185 13100
rect 8245 13040 8255 13100
rect 8175 13035 8255 13040
rect 8575 13210 8655 13215
rect 8575 13150 8585 13210
rect 8645 13150 8655 13210
rect 8575 13100 8655 13150
rect 8575 13040 8585 13100
rect 8645 13040 8655 13100
rect 8575 13035 8655 13040
rect 8975 13210 9055 13215
rect 8975 13150 8985 13210
rect 9045 13150 9055 13210
rect 8975 13100 9055 13150
rect 8975 13040 8985 13100
rect 9045 13040 9055 13100
rect 8975 13035 9055 13040
rect 9375 13210 9455 13215
rect 9375 13150 9385 13210
rect 9445 13150 9455 13210
rect 9375 13100 9455 13150
rect 9375 13040 9385 13100
rect 9445 13040 9455 13100
rect 9375 13035 9455 13040
rect 9775 13210 9855 13215
rect 9775 13150 9785 13210
rect 9845 13150 9855 13210
rect 9775 13100 9855 13150
rect 9775 13040 9785 13100
rect 9845 13040 9855 13100
rect 9775 13035 9855 13040
rect 10175 13210 10255 13215
rect 10175 13150 10185 13210
rect 10245 13150 10255 13210
rect 10175 13100 10255 13150
rect 10175 13040 10185 13100
rect 10245 13040 10255 13100
rect 10175 13035 10255 13040
rect 10575 13210 10655 13215
rect 10575 13150 10585 13210
rect 10645 13150 10655 13210
rect 10575 13100 10655 13150
rect 10575 13040 10585 13100
rect 10645 13040 10655 13100
rect 10575 13035 10655 13040
rect 10975 13210 11055 13215
rect 10975 13150 10985 13210
rect 11045 13150 11055 13210
rect 10975 13100 11055 13150
rect 10975 13040 10985 13100
rect 11045 13040 11055 13100
rect 10975 13035 11055 13040
rect 11375 13210 11455 13215
rect 11375 13150 11385 13210
rect 11445 13150 11455 13210
rect 11375 13100 11455 13150
rect 11375 13040 11385 13100
rect 11445 13040 11455 13100
rect 11375 13035 11455 13040
rect 11775 13210 11855 13215
rect 11775 13150 11785 13210
rect 11845 13150 11855 13210
rect 11775 13100 11855 13150
rect 11775 13040 11785 13100
rect 11845 13040 11855 13100
rect 11775 13035 11855 13040
rect 12175 13210 12255 13215
rect 12175 13150 12185 13210
rect 12245 13150 12255 13210
rect 12175 13100 12255 13150
rect 12175 13040 12185 13100
rect 12245 13040 12255 13100
rect 12175 13035 12255 13040
rect 12575 13210 12655 13215
rect 12575 13150 12585 13210
rect 12645 13150 12655 13210
rect 12575 13100 12655 13150
rect 12575 13040 12585 13100
rect 12645 13040 12655 13100
rect 12575 13035 12655 13040
rect 12975 13210 13055 13215
rect 12975 13150 12985 13210
rect 13045 13150 13055 13210
rect 12975 13100 13055 13150
rect 12975 13040 12985 13100
rect 13045 13040 13055 13100
rect 12975 13035 13055 13040
rect -215 12845 -155 13035
rect 185 12845 245 13035
rect 585 12845 645 13035
rect 985 12845 1045 13035
rect 1385 12845 1445 13035
rect 1785 12845 1845 13035
rect 2185 12845 2245 13035
rect 2585 12845 2645 13035
rect 2985 12845 3045 13035
rect 3385 12845 3445 13035
rect 3785 12845 3845 13035
rect 4185 12845 4245 13035
rect 4585 12845 4645 13035
rect 4985 12845 5045 13035
rect 5385 12845 5445 13035
rect 5785 12845 5845 13035
rect 6185 12845 6245 13035
rect 6585 12845 6645 13035
rect 6985 12845 7045 13035
rect 7385 12845 7445 13035
rect 7785 12845 7845 13035
rect 8185 12845 8245 13035
rect 8585 12845 8645 13035
rect 8985 12845 9045 13035
rect 9385 12845 9445 13035
rect 9785 12845 9845 13035
rect 10185 12845 10245 13035
rect 10585 12845 10645 13035
rect 10985 12845 11045 13035
rect 11385 12845 11445 13035
rect 11785 12845 11845 13035
rect 12185 12845 12245 13035
rect 12585 12845 12645 13035
rect 12985 12845 13045 13035
rect -225 12840 -145 12845
rect -225 12780 -215 12840
rect -155 12780 -145 12840
rect -225 12730 -145 12780
rect -225 12670 -215 12730
rect -155 12670 -145 12730
rect -225 12665 -145 12670
rect 175 12840 255 12845
rect 175 12780 185 12840
rect 245 12780 255 12840
rect 175 12730 255 12780
rect 175 12670 185 12730
rect 245 12670 255 12730
rect 175 12665 255 12670
rect 575 12840 655 12845
rect 575 12780 585 12840
rect 645 12780 655 12840
rect 575 12730 655 12780
rect 575 12670 585 12730
rect 645 12670 655 12730
rect 575 12665 655 12670
rect 975 12840 1055 12845
rect 975 12780 985 12840
rect 1045 12780 1055 12840
rect 975 12730 1055 12780
rect 975 12670 985 12730
rect 1045 12670 1055 12730
rect 975 12665 1055 12670
rect 1375 12840 1455 12845
rect 1375 12780 1385 12840
rect 1445 12780 1455 12840
rect 1375 12730 1455 12780
rect 1375 12670 1385 12730
rect 1445 12670 1455 12730
rect 1375 12665 1455 12670
rect 1775 12840 1855 12845
rect 1775 12780 1785 12840
rect 1845 12780 1855 12840
rect 1775 12730 1855 12780
rect 1775 12670 1785 12730
rect 1845 12670 1855 12730
rect 1775 12665 1855 12670
rect 2175 12840 2255 12845
rect 2175 12780 2185 12840
rect 2245 12780 2255 12840
rect 2175 12730 2255 12780
rect 2175 12670 2185 12730
rect 2245 12670 2255 12730
rect 2175 12665 2255 12670
rect 2575 12840 2655 12845
rect 2575 12780 2585 12840
rect 2645 12780 2655 12840
rect 2575 12730 2655 12780
rect 2575 12670 2585 12730
rect 2645 12670 2655 12730
rect 2575 12665 2655 12670
rect 2975 12840 3055 12845
rect 2975 12780 2985 12840
rect 3045 12780 3055 12840
rect 2975 12730 3055 12780
rect 2975 12670 2985 12730
rect 3045 12670 3055 12730
rect 2975 12665 3055 12670
rect 3375 12840 3455 12845
rect 3375 12780 3385 12840
rect 3445 12780 3455 12840
rect 3375 12730 3455 12780
rect 3375 12670 3385 12730
rect 3445 12670 3455 12730
rect 3375 12665 3455 12670
rect 3775 12840 3855 12845
rect 3775 12780 3785 12840
rect 3845 12780 3855 12840
rect 3775 12730 3855 12780
rect 3775 12670 3785 12730
rect 3845 12670 3855 12730
rect 3775 12665 3855 12670
rect 4175 12840 4255 12845
rect 4175 12780 4185 12840
rect 4245 12780 4255 12840
rect 4175 12730 4255 12780
rect 4175 12670 4185 12730
rect 4245 12670 4255 12730
rect 4175 12665 4255 12670
rect 4575 12840 4655 12845
rect 4575 12780 4585 12840
rect 4645 12780 4655 12840
rect 4575 12730 4655 12780
rect 4575 12670 4585 12730
rect 4645 12670 4655 12730
rect 4575 12665 4655 12670
rect 4975 12840 5055 12845
rect 4975 12780 4985 12840
rect 5045 12780 5055 12840
rect 4975 12730 5055 12780
rect 4975 12670 4985 12730
rect 5045 12670 5055 12730
rect 4975 12665 5055 12670
rect 5375 12840 5455 12845
rect 5375 12780 5385 12840
rect 5445 12780 5455 12840
rect 5375 12730 5455 12780
rect 5375 12670 5385 12730
rect 5445 12670 5455 12730
rect 5375 12665 5455 12670
rect 5775 12840 5855 12845
rect 5775 12780 5785 12840
rect 5845 12780 5855 12840
rect 5775 12730 5855 12780
rect 5775 12670 5785 12730
rect 5845 12670 5855 12730
rect 5775 12665 5855 12670
rect 6175 12840 6255 12845
rect 6175 12780 6185 12840
rect 6245 12780 6255 12840
rect 6175 12730 6255 12780
rect 6175 12670 6185 12730
rect 6245 12670 6255 12730
rect 6175 12665 6255 12670
rect 6575 12840 6655 12845
rect 6575 12780 6585 12840
rect 6645 12780 6655 12840
rect 6575 12730 6655 12780
rect 6575 12670 6585 12730
rect 6645 12670 6655 12730
rect 6575 12665 6655 12670
rect 6975 12840 7055 12845
rect 6975 12780 6985 12840
rect 7045 12780 7055 12840
rect 6975 12730 7055 12780
rect 6975 12670 6985 12730
rect 7045 12670 7055 12730
rect 6975 12665 7055 12670
rect 7375 12840 7455 12845
rect 7375 12780 7385 12840
rect 7445 12780 7455 12840
rect 7375 12730 7455 12780
rect 7375 12670 7385 12730
rect 7445 12670 7455 12730
rect 7375 12665 7455 12670
rect 7775 12840 7855 12845
rect 7775 12780 7785 12840
rect 7845 12780 7855 12840
rect 7775 12730 7855 12780
rect 7775 12670 7785 12730
rect 7845 12670 7855 12730
rect 7775 12665 7855 12670
rect 8175 12840 8255 12845
rect 8175 12780 8185 12840
rect 8245 12780 8255 12840
rect 8175 12730 8255 12780
rect 8175 12670 8185 12730
rect 8245 12670 8255 12730
rect 8175 12665 8255 12670
rect 8575 12840 8655 12845
rect 8575 12780 8585 12840
rect 8645 12780 8655 12840
rect 8575 12730 8655 12780
rect 8575 12670 8585 12730
rect 8645 12670 8655 12730
rect 8575 12665 8655 12670
rect 8975 12840 9055 12845
rect 8975 12780 8985 12840
rect 9045 12780 9055 12840
rect 8975 12730 9055 12780
rect 8975 12670 8985 12730
rect 9045 12670 9055 12730
rect 8975 12665 9055 12670
rect 9375 12840 9455 12845
rect 9375 12780 9385 12840
rect 9445 12780 9455 12840
rect 9375 12730 9455 12780
rect 9375 12670 9385 12730
rect 9445 12670 9455 12730
rect 9375 12665 9455 12670
rect 9775 12840 9855 12845
rect 9775 12780 9785 12840
rect 9845 12780 9855 12840
rect 9775 12730 9855 12780
rect 9775 12670 9785 12730
rect 9845 12670 9855 12730
rect 9775 12665 9855 12670
rect 10175 12840 10255 12845
rect 10175 12780 10185 12840
rect 10245 12780 10255 12840
rect 10175 12730 10255 12780
rect 10175 12670 10185 12730
rect 10245 12670 10255 12730
rect 10175 12665 10255 12670
rect 10575 12840 10655 12845
rect 10575 12780 10585 12840
rect 10645 12780 10655 12840
rect 10575 12730 10655 12780
rect 10575 12670 10585 12730
rect 10645 12670 10655 12730
rect 10575 12665 10655 12670
rect 10975 12840 11055 12845
rect 10975 12780 10985 12840
rect 11045 12780 11055 12840
rect 10975 12730 11055 12780
rect 10975 12670 10985 12730
rect 11045 12670 11055 12730
rect 10975 12665 11055 12670
rect 11375 12840 11455 12845
rect 11375 12780 11385 12840
rect 11445 12780 11455 12840
rect 11375 12730 11455 12780
rect 11375 12670 11385 12730
rect 11445 12670 11455 12730
rect 11375 12665 11455 12670
rect 11775 12840 11855 12845
rect 11775 12780 11785 12840
rect 11845 12780 11855 12840
rect 11775 12730 11855 12780
rect 11775 12670 11785 12730
rect 11845 12670 11855 12730
rect 11775 12665 11855 12670
rect 12175 12840 12255 12845
rect 12175 12780 12185 12840
rect 12245 12780 12255 12840
rect 12175 12730 12255 12780
rect 12175 12670 12185 12730
rect 12245 12670 12255 12730
rect 12175 12665 12255 12670
rect 12575 12840 12655 12845
rect 12575 12780 12585 12840
rect 12645 12780 12655 12840
rect 12575 12730 12655 12780
rect 12575 12670 12585 12730
rect 12645 12670 12655 12730
rect 12575 12665 12655 12670
rect 12975 12840 13055 12845
rect 12975 12780 12985 12840
rect 13045 12780 13055 12840
rect 12975 12730 13055 12780
rect 12975 12670 12985 12730
rect 13045 12670 13055 12730
rect 12975 12665 13055 12670
rect -215 12475 -155 12665
rect 185 12475 245 12665
rect 585 12475 645 12665
rect 985 12475 1045 12665
rect 1385 12475 1445 12665
rect 1785 12475 1845 12665
rect 2185 12475 2245 12665
rect 2585 12475 2645 12665
rect 2985 12475 3045 12665
rect 3385 12475 3445 12665
rect 3785 12475 3845 12665
rect 4185 12475 4245 12665
rect 4585 12475 4645 12665
rect 4985 12475 5045 12665
rect 5385 12475 5445 12665
rect 5785 12475 5845 12665
rect 6185 12475 6245 12665
rect 6585 12475 6645 12665
rect 6985 12475 7045 12665
rect 7385 12475 7445 12665
rect 7785 12475 7845 12665
rect 8185 12475 8245 12665
rect 8585 12475 8645 12665
rect 8985 12475 9045 12665
rect 9385 12475 9445 12665
rect 9785 12475 9845 12665
rect 10185 12475 10245 12665
rect 10585 12475 10645 12665
rect 10985 12475 11045 12665
rect 11385 12475 11445 12665
rect 11785 12475 11845 12665
rect 12185 12475 12245 12665
rect 12585 12475 12645 12665
rect 12985 12475 13045 12665
rect -225 12470 -145 12475
rect -225 12410 -215 12470
rect -155 12410 -145 12470
rect -225 12360 -145 12410
rect -225 12300 -215 12360
rect -155 12300 -145 12360
rect -225 12295 -145 12300
rect 175 12470 255 12475
rect 175 12410 185 12470
rect 245 12410 255 12470
rect 175 12360 255 12410
rect 175 12300 185 12360
rect 245 12300 255 12360
rect 175 12295 255 12300
rect 575 12470 655 12475
rect 575 12410 585 12470
rect 645 12410 655 12470
rect 575 12360 655 12410
rect 575 12300 585 12360
rect 645 12300 655 12360
rect 575 12295 655 12300
rect 975 12470 1055 12475
rect 975 12410 985 12470
rect 1045 12410 1055 12470
rect 975 12360 1055 12410
rect 975 12300 985 12360
rect 1045 12300 1055 12360
rect 975 12295 1055 12300
rect 1375 12470 1455 12475
rect 1375 12410 1385 12470
rect 1445 12410 1455 12470
rect 1375 12360 1455 12410
rect 1375 12300 1385 12360
rect 1445 12300 1455 12360
rect 1375 12295 1455 12300
rect 1775 12470 1855 12475
rect 1775 12410 1785 12470
rect 1845 12410 1855 12470
rect 1775 12360 1855 12410
rect 1775 12300 1785 12360
rect 1845 12300 1855 12360
rect 1775 12295 1855 12300
rect 2175 12470 2255 12475
rect 2175 12410 2185 12470
rect 2245 12410 2255 12470
rect 2175 12360 2255 12410
rect 2175 12300 2185 12360
rect 2245 12300 2255 12360
rect 2175 12295 2255 12300
rect 2575 12470 2655 12475
rect 2575 12410 2585 12470
rect 2645 12410 2655 12470
rect 2575 12360 2655 12410
rect 2575 12300 2585 12360
rect 2645 12300 2655 12360
rect 2575 12295 2655 12300
rect 2975 12470 3055 12475
rect 2975 12410 2985 12470
rect 3045 12410 3055 12470
rect 2975 12360 3055 12410
rect 2975 12300 2985 12360
rect 3045 12300 3055 12360
rect 2975 12295 3055 12300
rect 3375 12470 3455 12475
rect 3375 12410 3385 12470
rect 3445 12410 3455 12470
rect 3375 12360 3455 12410
rect 3375 12300 3385 12360
rect 3445 12300 3455 12360
rect 3375 12295 3455 12300
rect 3775 12470 3855 12475
rect 3775 12410 3785 12470
rect 3845 12410 3855 12470
rect 3775 12360 3855 12410
rect 3775 12300 3785 12360
rect 3845 12300 3855 12360
rect 3775 12295 3855 12300
rect 4175 12470 4255 12475
rect 4175 12410 4185 12470
rect 4245 12410 4255 12470
rect 4175 12360 4255 12410
rect 4175 12300 4185 12360
rect 4245 12300 4255 12360
rect 4175 12295 4255 12300
rect 4575 12470 4655 12475
rect 4575 12410 4585 12470
rect 4645 12410 4655 12470
rect 4575 12360 4655 12410
rect 4575 12300 4585 12360
rect 4645 12300 4655 12360
rect 4575 12295 4655 12300
rect 4975 12470 5055 12475
rect 4975 12410 4985 12470
rect 5045 12410 5055 12470
rect 4975 12360 5055 12410
rect 4975 12300 4985 12360
rect 5045 12300 5055 12360
rect 4975 12295 5055 12300
rect 5375 12470 5455 12475
rect 5375 12410 5385 12470
rect 5445 12410 5455 12470
rect 5375 12360 5455 12410
rect 5375 12300 5385 12360
rect 5445 12300 5455 12360
rect 5375 12295 5455 12300
rect 5775 12470 5855 12475
rect 5775 12410 5785 12470
rect 5845 12410 5855 12470
rect 5775 12360 5855 12410
rect 5775 12300 5785 12360
rect 5845 12300 5855 12360
rect 5775 12295 5855 12300
rect 6175 12470 6255 12475
rect 6175 12410 6185 12470
rect 6245 12410 6255 12470
rect 6175 12360 6255 12410
rect 6175 12300 6185 12360
rect 6245 12300 6255 12360
rect 6175 12295 6255 12300
rect 6575 12470 6655 12475
rect 6575 12410 6585 12470
rect 6645 12410 6655 12470
rect 6575 12360 6655 12410
rect 6575 12300 6585 12360
rect 6645 12300 6655 12360
rect 6575 12295 6655 12300
rect 6975 12470 7055 12475
rect 6975 12410 6985 12470
rect 7045 12410 7055 12470
rect 6975 12360 7055 12410
rect 6975 12300 6985 12360
rect 7045 12300 7055 12360
rect 6975 12295 7055 12300
rect 7375 12470 7455 12475
rect 7375 12410 7385 12470
rect 7445 12410 7455 12470
rect 7375 12360 7455 12410
rect 7375 12300 7385 12360
rect 7445 12300 7455 12360
rect 7375 12295 7455 12300
rect 7775 12470 7855 12475
rect 7775 12410 7785 12470
rect 7845 12410 7855 12470
rect 7775 12360 7855 12410
rect 7775 12300 7785 12360
rect 7845 12300 7855 12360
rect 7775 12295 7855 12300
rect 8175 12470 8255 12475
rect 8175 12410 8185 12470
rect 8245 12410 8255 12470
rect 8175 12360 8255 12410
rect 8175 12300 8185 12360
rect 8245 12300 8255 12360
rect 8175 12295 8255 12300
rect 8575 12470 8655 12475
rect 8575 12410 8585 12470
rect 8645 12410 8655 12470
rect 8575 12360 8655 12410
rect 8575 12300 8585 12360
rect 8645 12300 8655 12360
rect 8575 12295 8655 12300
rect 8975 12470 9055 12475
rect 8975 12410 8985 12470
rect 9045 12410 9055 12470
rect 8975 12360 9055 12410
rect 8975 12300 8985 12360
rect 9045 12300 9055 12360
rect 8975 12295 9055 12300
rect 9375 12470 9455 12475
rect 9375 12410 9385 12470
rect 9445 12410 9455 12470
rect 9375 12360 9455 12410
rect 9375 12300 9385 12360
rect 9445 12300 9455 12360
rect 9375 12295 9455 12300
rect 9775 12470 9855 12475
rect 9775 12410 9785 12470
rect 9845 12410 9855 12470
rect 9775 12360 9855 12410
rect 9775 12300 9785 12360
rect 9845 12300 9855 12360
rect 9775 12295 9855 12300
rect 10175 12470 10255 12475
rect 10175 12410 10185 12470
rect 10245 12410 10255 12470
rect 10175 12360 10255 12410
rect 10175 12300 10185 12360
rect 10245 12300 10255 12360
rect 10175 12295 10255 12300
rect 10575 12470 10655 12475
rect 10575 12410 10585 12470
rect 10645 12410 10655 12470
rect 10575 12360 10655 12410
rect 10575 12300 10585 12360
rect 10645 12300 10655 12360
rect 10575 12295 10655 12300
rect 10975 12470 11055 12475
rect 10975 12410 10985 12470
rect 11045 12410 11055 12470
rect 10975 12360 11055 12410
rect 10975 12300 10985 12360
rect 11045 12300 11055 12360
rect 10975 12295 11055 12300
rect 11375 12470 11455 12475
rect 11375 12410 11385 12470
rect 11445 12410 11455 12470
rect 11375 12360 11455 12410
rect 11375 12300 11385 12360
rect 11445 12300 11455 12360
rect 11375 12295 11455 12300
rect 11775 12470 11855 12475
rect 11775 12410 11785 12470
rect 11845 12410 11855 12470
rect 11775 12360 11855 12410
rect 11775 12300 11785 12360
rect 11845 12300 11855 12360
rect 11775 12295 11855 12300
rect 12175 12470 12255 12475
rect 12175 12410 12185 12470
rect 12245 12410 12255 12470
rect 12175 12360 12255 12410
rect 12175 12300 12185 12360
rect 12245 12300 12255 12360
rect 12175 12295 12255 12300
rect 12575 12470 12655 12475
rect 12575 12410 12585 12470
rect 12645 12410 12655 12470
rect 12575 12360 12655 12410
rect 12575 12300 12585 12360
rect 12645 12300 12655 12360
rect 12575 12295 12655 12300
rect 12975 12470 13055 12475
rect 12975 12410 12985 12470
rect 13045 12410 13055 12470
rect 12975 12360 13055 12410
rect 12975 12300 12985 12360
rect 13045 12300 13055 12360
rect 12975 12295 13055 12300
rect -215 12105 -155 12295
rect 185 12105 245 12295
rect 585 12105 645 12295
rect 985 12105 1045 12295
rect 1385 12105 1445 12295
rect 1785 12105 1845 12295
rect 2185 12105 2245 12295
rect 2585 12105 2645 12295
rect 2985 12105 3045 12295
rect 3385 12105 3445 12295
rect 3785 12105 3845 12295
rect 4185 12105 4245 12295
rect 4585 12105 4645 12295
rect 4985 12105 5045 12295
rect 5385 12105 5445 12295
rect 5785 12105 5845 12295
rect 6185 12105 6245 12295
rect 6585 12105 6645 12295
rect 6985 12105 7045 12295
rect 7385 12105 7445 12295
rect 7785 12105 7845 12295
rect 8185 12105 8245 12295
rect 8585 12105 8645 12295
rect 8985 12105 9045 12295
rect 9385 12105 9445 12295
rect 9785 12105 9845 12295
rect 10185 12105 10245 12295
rect 10585 12105 10645 12295
rect 10985 12105 11045 12295
rect 11385 12105 11445 12295
rect 11785 12105 11845 12295
rect 12185 12105 12245 12295
rect 12585 12105 12645 12295
rect 12985 12105 13045 12295
rect -225 12100 -145 12105
rect -225 12040 -215 12100
rect -155 12040 -145 12100
rect -225 11990 -145 12040
rect -225 11930 -215 11990
rect -155 11930 -145 11990
rect -225 11925 -145 11930
rect 175 12100 255 12105
rect 175 12040 185 12100
rect 245 12040 255 12100
rect 175 11990 255 12040
rect 175 11930 185 11990
rect 245 11930 255 11990
rect 175 11925 255 11930
rect 575 12100 655 12105
rect 575 12040 585 12100
rect 645 12040 655 12100
rect 575 11990 655 12040
rect 575 11930 585 11990
rect 645 11930 655 11990
rect 575 11925 655 11930
rect 975 12100 1055 12105
rect 975 12040 985 12100
rect 1045 12040 1055 12100
rect 975 11990 1055 12040
rect 975 11930 985 11990
rect 1045 11930 1055 11990
rect 975 11925 1055 11930
rect 1375 12100 1455 12105
rect 1375 12040 1385 12100
rect 1445 12040 1455 12100
rect 1375 11990 1455 12040
rect 1375 11930 1385 11990
rect 1445 11930 1455 11990
rect 1375 11925 1455 11930
rect 1775 12100 1855 12105
rect 1775 12040 1785 12100
rect 1845 12040 1855 12100
rect 1775 11990 1855 12040
rect 1775 11930 1785 11990
rect 1845 11930 1855 11990
rect 1775 11925 1855 11930
rect 2175 12100 2255 12105
rect 2175 12040 2185 12100
rect 2245 12040 2255 12100
rect 2175 11990 2255 12040
rect 2175 11930 2185 11990
rect 2245 11930 2255 11990
rect 2175 11925 2255 11930
rect 2575 12100 2655 12105
rect 2575 12040 2585 12100
rect 2645 12040 2655 12100
rect 2575 11990 2655 12040
rect 2575 11930 2585 11990
rect 2645 11930 2655 11990
rect 2575 11925 2655 11930
rect 2975 12100 3055 12105
rect 2975 12040 2985 12100
rect 3045 12040 3055 12100
rect 2975 11990 3055 12040
rect 2975 11930 2985 11990
rect 3045 11930 3055 11990
rect 2975 11925 3055 11930
rect 3375 12100 3455 12105
rect 3375 12040 3385 12100
rect 3445 12040 3455 12100
rect 3375 11990 3455 12040
rect 3375 11930 3385 11990
rect 3445 11930 3455 11990
rect 3375 11925 3455 11930
rect 3775 12100 3855 12105
rect 3775 12040 3785 12100
rect 3845 12040 3855 12100
rect 3775 11990 3855 12040
rect 3775 11930 3785 11990
rect 3845 11930 3855 11990
rect 3775 11925 3855 11930
rect 4175 12100 4255 12105
rect 4175 12040 4185 12100
rect 4245 12040 4255 12100
rect 4175 11990 4255 12040
rect 4175 11930 4185 11990
rect 4245 11930 4255 11990
rect 4175 11925 4255 11930
rect 4575 12100 4655 12105
rect 4575 12040 4585 12100
rect 4645 12040 4655 12100
rect 4575 11990 4655 12040
rect 4575 11930 4585 11990
rect 4645 11930 4655 11990
rect 4575 11925 4655 11930
rect 4975 12100 5055 12105
rect 4975 12040 4985 12100
rect 5045 12040 5055 12100
rect 4975 11990 5055 12040
rect 4975 11930 4985 11990
rect 5045 11930 5055 11990
rect 4975 11925 5055 11930
rect 5375 12100 5455 12105
rect 5375 12040 5385 12100
rect 5445 12040 5455 12100
rect 5375 11990 5455 12040
rect 5375 11930 5385 11990
rect 5445 11930 5455 11990
rect 5375 11925 5455 11930
rect 5775 12100 5855 12105
rect 5775 12040 5785 12100
rect 5845 12040 5855 12100
rect 5775 11990 5855 12040
rect 5775 11930 5785 11990
rect 5845 11930 5855 11990
rect 5775 11925 5855 11930
rect 6175 12100 6255 12105
rect 6175 12040 6185 12100
rect 6245 12040 6255 12100
rect 6175 11990 6255 12040
rect 6175 11930 6185 11990
rect 6245 11930 6255 11990
rect 6175 11925 6255 11930
rect 6575 12100 6655 12105
rect 6575 12040 6585 12100
rect 6645 12040 6655 12100
rect 6575 11990 6655 12040
rect 6575 11930 6585 11990
rect 6645 11930 6655 11990
rect 6575 11925 6655 11930
rect 6975 12100 7055 12105
rect 6975 12040 6985 12100
rect 7045 12040 7055 12100
rect 6975 11990 7055 12040
rect 6975 11930 6985 11990
rect 7045 11930 7055 11990
rect 6975 11925 7055 11930
rect 7375 12100 7455 12105
rect 7375 12040 7385 12100
rect 7445 12040 7455 12100
rect 7375 11990 7455 12040
rect 7375 11930 7385 11990
rect 7445 11930 7455 11990
rect 7375 11925 7455 11930
rect 7775 12100 7855 12105
rect 7775 12040 7785 12100
rect 7845 12040 7855 12100
rect 7775 11990 7855 12040
rect 7775 11930 7785 11990
rect 7845 11930 7855 11990
rect 7775 11925 7855 11930
rect 8175 12100 8255 12105
rect 8175 12040 8185 12100
rect 8245 12040 8255 12100
rect 8175 11990 8255 12040
rect 8175 11930 8185 11990
rect 8245 11930 8255 11990
rect 8175 11925 8255 11930
rect 8575 12100 8655 12105
rect 8575 12040 8585 12100
rect 8645 12040 8655 12100
rect 8575 11990 8655 12040
rect 8575 11930 8585 11990
rect 8645 11930 8655 11990
rect 8575 11925 8655 11930
rect 8975 12100 9055 12105
rect 8975 12040 8985 12100
rect 9045 12040 9055 12100
rect 8975 11990 9055 12040
rect 8975 11930 8985 11990
rect 9045 11930 9055 11990
rect 8975 11925 9055 11930
rect 9375 12100 9455 12105
rect 9375 12040 9385 12100
rect 9445 12040 9455 12100
rect 9375 11990 9455 12040
rect 9375 11930 9385 11990
rect 9445 11930 9455 11990
rect 9375 11925 9455 11930
rect 9775 12100 9855 12105
rect 9775 12040 9785 12100
rect 9845 12040 9855 12100
rect 9775 11990 9855 12040
rect 9775 11930 9785 11990
rect 9845 11930 9855 11990
rect 9775 11925 9855 11930
rect 10175 12100 10255 12105
rect 10175 12040 10185 12100
rect 10245 12040 10255 12100
rect 10175 11990 10255 12040
rect 10175 11930 10185 11990
rect 10245 11930 10255 11990
rect 10175 11925 10255 11930
rect 10575 12100 10655 12105
rect 10575 12040 10585 12100
rect 10645 12040 10655 12100
rect 10575 11990 10655 12040
rect 10575 11930 10585 11990
rect 10645 11930 10655 11990
rect 10575 11925 10655 11930
rect 10975 12100 11055 12105
rect 10975 12040 10985 12100
rect 11045 12040 11055 12100
rect 10975 11990 11055 12040
rect 10975 11930 10985 11990
rect 11045 11930 11055 11990
rect 10975 11925 11055 11930
rect 11375 12100 11455 12105
rect 11375 12040 11385 12100
rect 11445 12040 11455 12100
rect 11375 11990 11455 12040
rect 11375 11930 11385 11990
rect 11445 11930 11455 11990
rect 11375 11925 11455 11930
rect 11775 12100 11855 12105
rect 11775 12040 11785 12100
rect 11845 12040 11855 12100
rect 11775 11990 11855 12040
rect 11775 11930 11785 11990
rect 11845 11930 11855 11990
rect 11775 11925 11855 11930
rect 12175 12100 12255 12105
rect 12175 12040 12185 12100
rect 12245 12040 12255 12100
rect 12175 11990 12255 12040
rect 12175 11930 12185 11990
rect 12245 11930 12255 11990
rect 12175 11925 12255 11930
rect 12575 12100 12655 12105
rect 12575 12040 12585 12100
rect 12645 12040 12655 12100
rect 12575 11990 12655 12040
rect 12575 11930 12585 11990
rect 12645 11930 12655 11990
rect 12575 11925 12655 11930
rect 12975 12100 13055 12105
rect 12975 12040 12985 12100
rect 13045 12040 13055 12100
rect 12975 11990 13055 12040
rect 12975 11930 12985 11990
rect 13045 11930 13055 11990
rect 12975 11925 13055 11930
rect -215 11735 -155 11925
rect 185 11735 245 11925
rect 585 11735 645 11925
rect 985 11735 1045 11925
rect 1385 11735 1445 11925
rect 1785 11735 1845 11925
rect 2185 11735 2245 11925
rect 2585 11735 2645 11925
rect 2985 11735 3045 11925
rect 3385 11735 3445 11925
rect 3785 11735 3845 11925
rect 4185 11735 4245 11925
rect 4585 11735 4645 11925
rect 4985 11735 5045 11925
rect 5385 11735 5445 11925
rect 5785 11735 5845 11925
rect 6185 11735 6245 11925
rect 6585 11735 6645 11925
rect 6985 11735 7045 11925
rect 7385 11735 7445 11925
rect 7785 11735 7845 11925
rect 8185 11735 8245 11925
rect 8585 11735 8645 11925
rect 8985 11735 9045 11925
rect 9385 11735 9445 11925
rect 9785 11735 9845 11925
rect 10185 11735 10245 11925
rect 10585 11735 10645 11925
rect 10985 11735 11045 11925
rect 11385 11735 11445 11925
rect 11785 11735 11845 11925
rect 12185 11735 12245 11925
rect 12585 11735 12645 11925
rect 12985 11735 13045 11925
rect -225 11730 -145 11735
rect -225 11670 -215 11730
rect -155 11670 -145 11730
rect -225 11620 -145 11670
rect -225 11560 -215 11620
rect -155 11560 -145 11620
rect -225 11555 -145 11560
rect 175 11730 255 11735
rect 175 11670 185 11730
rect 245 11670 255 11730
rect 175 11620 255 11670
rect 175 11560 185 11620
rect 245 11560 255 11620
rect 175 11555 255 11560
rect 575 11730 655 11735
rect 575 11670 585 11730
rect 645 11670 655 11730
rect 575 11620 655 11670
rect 575 11560 585 11620
rect 645 11560 655 11620
rect 575 11555 655 11560
rect 975 11730 1055 11735
rect 975 11670 985 11730
rect 1045 11670 1055 11730
rect 975 11620 1055 11670
rect 975 11560 985 11620
rect 1045 11560 1055 11620
rect 975 11555 1055 11560
rect 1375 11730 1455 11735
rect 1375 11670 1385 11730
rect 1445 11670 1455 11730
rect 1375 11620 1455 11670
rect 1375 11560 1385 11620
rect 1445 11560 1455 11620
rect 1375 11555 1455 11560
rect 1775 11730 1855 11735
rect 1775 11670 1785 11730
rect 1845 11670 1855 11730
rect 1775 11620 1855 11670
rect 1775 11560 1785 11620
rect 1845 11560 1855 11620
rect 1775 11555 1855 11560
rect 2175 11730 2255 11735
rect 2175 11670 2185 11730
rect 2245 11670 2255 11730
rect 2175 11620 2255 11670
rect 2175 11560 2185 11620
rect 2245 11560 2255 11620
rect 2175 11555 2255 11560
rect 2575 11730 2655 11735
rect 2575 11670 2585 11730
rect 2645 11670 2655 11730
rect 2575 11620 2655 11670
rect 2575 11560 2585 11620
rect 2645 11560 2655 11620
rect 2575 11555 2655 11560
rect 2975 11730 3055 11735
rect 2975 11670 2985 11730
rect 3045 11670 3055 11730
rect 2975 11620 3055 11670
rect 2975 11560 2985 11620
rect 3045 11560 3055 11620
rect 2975 11555 3055 11560
rect 3375 11730 3455 11735
rect 3375 11670 3385 11730
rect 3445 11670 3455 11730
rect 3375 11620 3455 11670
rect 3375 11560 3385 11620
rect 3445 11560 3455 11620
rect 3375 11555 3455 11560
rect 3775 11730 3855 11735
rect 3775 11670 3785 11730
rect 3845 11670 3855 11730
rect 3775 11620 3855 11670
rect 3775 11560 3785 11620
rect 3845 11560 3855 11620
rect 3775 11555 3855 11560
rect 4175 11730 4255 11735
rect 4175 11670 4185 11730
rect 4245 11670 4255 11730
rect 4175 11620 4255 11670
rect 4175 11560 4185 11620
rect 4245 11560 4255 11620
rect 4175 11555 4255 11560
rect 4575 11730 4655 11735
rect 4575 11670 4585 11730
rect 4645 11670 4655 11730
rect 4575 11620 4655 11670
rect 4575 11560 4585 11620
rect 4645 11560 4655 11620
rect 4575 11555 4655 11560
rect 4975 11730 5055 11735
rect 4975 11670 4985 11730
rect 5045 11670 5055 11730
rect 4975 11620 5055 11670
rect 4975 11560 4985 11620
rect 5045 11560 5055 11620
rect 4975 11555 5055 11560
rect 5375 11730 5455 11735
rect 5375 11670 5385 11730
rect 5445 11670 5455 11730
rect 5375 11620 5455 11670
rect 5375 11560 5385 11620
rect 5445 11560 5455 11620
rect 5375 11555 5455 11560
rect 5775 11730 5855 11735
rect 5775 11670 5785 11730
rect 5845 11670 5855 11730
rect 5775 11620 5855 11670
rect 5775 11560 5785 11620
rect 5845 11560 5855 11620
rect 5775 11555 5855 11560
rect 6175 11730 6255 11735
rect 6175 11670 6185 11730
rect 6245 11670 6255 11730
rect 6175 11620 6255 11670
rect 6175 11560 6185 11620
rect 6245 11560 6255 11620
rect 6175 11555 6255 11560
rect 6575 11730 6655 11735
rect 6575 11670 6585 11730
rect 6645 11670 6655 11730
rect 6575 11620 6655 11670
rect 6575 11560 6585 11620
rect 6645 11560 6655 11620
rect 6575 11555 6655 11560
rect 6975 11730 7055 11735
rect 6975 11670 6985 11730
rect 7045 11670 7055 11730
rect 6975 11620 7055 11670
rect 6975 11560 6985 11620
rect 7045 11560 7055 11620
rect 6975 11555 7055 11560
rect 7375 11730 7455 11735
rect 7375 11670 7385 11730
rect 7445 11670 7455 11730
rect 7375 11620 7455 11670
rect 7375 11560 7385 11620
rect 7445 11560 7455 11620
rect 7375 11555 7455 11560
rect 7775 11730 7855 11735
rect 7775 11670 7785 11730
rect 7845 11670 7855 11730
rect 7775 11620 7855 11670
rect 7775 11560 7785 11620
rect 7845 11560 7855 11620
rect 7775 11555 7855 11560
rect 8175 11730 8255 11735
rect 8175 11670 8185 11730
rect 8245 11670 8255 11730
rect 8175 11620 8255 11670
rect 8175 11560 8185 11620
rect 8245 11560 8255 11620
rect 8175 11555 8255 11560
rect 8575 11730 8655 11735
rect 8575 11670 8585 11730
rect 8645 11670 8655 11730
rect 8575 11620 8655 11670
rect 8575 11560 8585 11620
rect 8645 11560 8655 11620
rect 8575 11555 8655 11560
rect 8975 11730 9055 11735
rect 8975 11670 8985 11730
rect 9045 11670 9055 11730
rect 8975 11620 9055 11670
rect 8975 11560 8985 11620
rect 9045 11560 9055 11620
rect 8975 11555 9055 11560
rect 9375 11730 9455 11735
rect 9375 11670 9385 11730
rect 9445 11670 9455 11730
rect 9375 11620 9455 11670
rect 9375 11560 9385 11620
rect 9445 11560 9455 11620
rect 9375 11555 9455 11560
rect 9775 11730 9855 11735
rect 9775 11670 9785 11730
rect 9845 11670 9855 11730
rect 9775 11620 9855 11670
rect 9775 11560 9785 11620
rect 9845 11560 9855 11620
rect 9775 11555 9855 11560
rect 10175 11730 10255 11735
rect 10175 11670 10185 11730
rect 10245 11670 10255 11730
rect 10175 11620 10255 11670
rect 10175 11560 10185 11620
rect 10245 11560 10255 11620
rect 10175 11555 10255 11560
rect 10575 11730 10655 11735
rect 10575 11670 10585 11730
rect 10645 11670 10655 11730
rect 10575 11620 10655 11670
rect 10575 11560 10585 11620
rect 10645 11560 10655 11620
rect 10575 11555 10655 11560
rect 10975 11730 11055 11735
rect 10975 11670 10985 11730
rect 11045 11670 11055 11730
rect 10975 11620 11055 11670
rect 10975 11560 10985 11620
rect 11045 11560 11055 11620
rect 10975 11555 11055 11560
rect 11375 11730 11455 11735
rect 11375 11670 11385 11730
rect 11445 11670 11455 11730
rect 11375 11620 11455 11670
rect 11375 11560 11385 11620
rect 11445 11560 11455 11620
rect 11375 11555 11455 11560
rect 11775 11730 11855 11735
rect 11775 11670 11785 11730
rect 11845 11670 11855 11730
rect 11775 11620 11855 11670
rect 11775 11560 11785 11620
rect 11845 11560 11855 11620
rect 11775 11555 11855 11560
rect 12175 11730 12255 11735
rect 12175 11670 12185 11730
rect 12245 11670 12255 11730
rect 12175 11620 12255 11670
rect 12175 11560 12185 11620
rect 12245 11560 12255 11620
rect 12175 11555 12255 11560
rect 12575 11730 12655 11735
rect 12575 11670 12585 11730
rect 12645 11670 12655 11730
rect 12575 11620 12655 11670
rect 12575 11560 12585 11620
rect 12645 11560 12655 11620
rect 12575 11555 12655 11560
rect 12975 11730 13055 11735
rect 12975 11670 12985 11730
rect 13045 11670 13055 11730
rect 12975 11620 13055 11670
rect 12975 11560 12985 11620
rect 13045 11560 13055 11620
rect 12975 11555 13055 11560
rect -215 11365 -155 11555
rect 185 11365 245 11555
rect 585 11365 645 11555
rect 985 11365 1045 11555
rect 1385 11365 1445 11555
rect 1785 11365 1845 11555
rect 2185 11365 2245 11555
rect 2585 11365 2645 11555
rect 2985 11365 3045 11555
rect 3385 11365 3445 11555
rect 3785 11365 3845 11555
rect 4185 11365 4245 11555
rect 4585 11365 4645 11555
rect 4985 11365 5045 11555
rect 5385 11365 5445 11555
rect 5785 11365 5845 11555
rect 6185 11365 6245 11555
rect 6585 11365 6645 11555
rect 6985 11365 7045 11555
rect 7385 11365 7445 11555
rect 7785 11365 7845 11555
rect 8185 11365 8245 11555
rect 8585 11365 8645 11555
rect 8985 11365 9045 11555
rect 9385 11365 9445 11555
rect 9785 11365 9845 11555
rect 10185 11365 10245 11555
rect 10585 11365 10645 11555
rect 10985 11365 11045 11555
rect 11385 11365 11445 11555
rect 11785 11365 11845 11555
rect 12185 11365 12245 11555
rect 12585 11365 12645 11555
rect 12985 11365 13045 11555
rect -225 11360 -145 11365
rect -225 11300 -215 11360
rect -155 11300 -145 11360
rect -225 11250 -145 11300
rect -225 11190 -215 11250
rect -155 11190 -145 11250
rect -225 11185 -145 11190
rect 175 11360 255 11365
rect 175 11300 185 11360
rect 245 11300 255 11360
rect 175 11250 255 11300
rect 175 11190 185 11250
rect 245 11190 255 11250
rect 175 11185 255 11190
rect 575 11360 655 11365
rect 575 11300 585 11360
rect 645 11300 655 11360
rect 575 11250 655 11300
rect 575 11190 585 11250
rect 645 11190 655 11250
rect 575 11185 655 11190
rect 975 11360 1055 11365
rect 975 11300 985 11360
rect 1045 11300 1055 11360
rect 975 11250 1055 11300
rect 975 11190 985 11250
rect 1045 11190 1055 11250
rect 975 11185 1055 11190
rect 1375 11360 1455 11365
rect 1375 11300 1385 11360
rect 1445 11300 1455 11360
rect 1375 11250 1455 11300
rect 1375 11190 1385 11250
rect 1445 11190 1455 11250
rect 1375 11185 1455 11190
rect 1775 11360 1855 11365
rect 1775 11300 1785 11360
rect 1845 11300 1855 11360
rect 1775 11250 1855 11300
rect 1775 11190 1785 11250
rect 1845 11190 1855 11250
rect 1775 11185 1855 11190
rect 2175 11360 2255 11365
rect 2175 11300 2185 11360
rect 2245 11300 2255 11360
rect 2175 11250 2255 11300
rect 2175 11190 2185 11250
rect 2245 11190 2255 11250
rect 2175 11185 2255 11190
rect 2575 11360 2655 11365
rect 2575 11300 2585 11360
rect 2645 11300 2655 11360
rect 2575 11250 2655 11300
rect 2575 11190 2585 11250
rect 2645 11190 2655 11250
rect 2575 11185 2655 11190
rect 2975 11360 3055 11365
rect 2975 11300 2985 11360
rect 3045 11300 3055 11360
rect 2975 11250 3055 11300
rect 2975 11190 2985 11250
rect 3045 11190 3055 11250
rect 2975 11185 3055 11190
rect 3375 11360 3455 11365
rect 3375 11300 3385 11360
rect 3445 11300 3455 11360
rect 3375 11250 3455 11300
rect 3375 11190 3385 11250
rect 3445 11190 3455 11250
rect 3375 11185 3455 11190
rect 3775 11360 3855 11365
rect 3775 11300 3785 11360
rect 3845 11300 3855 11360
rect 3775 11250 3855 11300
rect 3775 11190 3785 11250
rect 3845 11190 3855 11250
rect 3775 11185 3855 11190
rect 4175 11360 4255 11365
rect 4175 11300 4185 11360
rect 4245 11300 4255 11360
rect 4175 11250 4255 11300
rect 4175 11190 4185 11250
rect 4245 11190 4255 11250
rect 4175 11185 4255 11190
rect 4575 11360 4655 11365
rect 4575 11300 4585 11360
rect 4645 11300 4655 11360
rect 4575 11250 4655 11300
rect 4575 11190 4585 11250
rect 4645 11190 4655 11250
rect 4575 11185 4655 11190
rect 4975 11360 5055 11365
rect 4975 11300 4985 11360
rect 5045 11300 5055 11360
rect 4975 11250 5055 11300
rect 4975 11190 4985 11250
rect 5045 11190 5055 11250
rect 4975 11185 5055 11190
rect 5375 11360 5455 11365
rect 5375 11300 5385 11360
rect 5445 11300 5455 11360
rect 5375 11250 5455 11300
rect 5375 11190 5385 11250
rect 5445 11190 5455 11250
rect 5375 11185 5455 11190
rect 5775 11360 5855 11365
rect 5775 11300 5785 11360
rect 5845 11300 5855 11360
rect 5775 11250 5855 11300
rect 5775 11190 5785 11250
rect 5845 11190 5855 11250
rect 5775 11185 5855 11190
rect 6175 11360 6255 11365
rect 6175 11300 6185 11360
rect 6245 11300 6255 11360
rect 6175 11250 6255 11300
rect 6175 11190 6185 11250
rect 6245 11190 6255 11250
rect 6175 11185 6255 11190
rect 6575 11360 6655 11365
rect 6575 11300 6585 11360
rect 6645 11300 6655 11360
rect 6575 11250 6655 11300
rect 6575 11190 6585 11250
rect 6645 11190 6655 11250
rect 6575 11185 6655 11190
rect 6975 11360 7055 11365
rect 6975 11300 6985 11360
rect 7045 11300 7055 11360
rect 6975 11250 7055 11300
rect 6975 11190 6985 11250
rect 7045 11190 7055 11250
rect 6975 11185 7055 11190
rect 7375 11360 7455 11365
rect 7375 11300 7385 11360
rect 7445 11300 7455 11360
rect 7375 11250 7455 11300
rect 7375 11190 7385 11250
rect 7445 11190 7455 11250
rect 7375 11185 7455 11190
rect 7775 11360 7855 11365
rect 7775 11300 7785 11360
rect 7845 11300 7855 11360
rect 7775 11250 7855 11300
rect 7775 11190 7785 11250
rect 7845 11190 7855 11250
rect 7775 11185 7855 11190
rect 8175 11360 8255 11365
rect 8175 11300 8185 11360
rect 8245 11300 8255 11360
rect 8175 11250 8255 11300
rect 8175 11190 8185 11250
rect 8245 11190 8255 11250
rect 8175 11185 8255 11190
rect 8575 11360 8655 11365
rect 8575 11300 8585 11360
rect 8645 11300 8655 11360
rect 8575 11250 8655 11300
rect 8575 11190 8585 11250
rect 8645 11190 8655 11250
rect 8575 11185 8655 11190
rect 8975 11360 9055 11365
rect 8975 11300 8985 11360
rect 9045 11300 9055 11360
rect 8975 11250 9055 11300
rect 8975 11190 8985 11250
rect 9045 11190 9055 11250
rect 8975 11185 9055 11190
rect 9375 11360 9455 11365
rect 9375 11300 9385 11360
rect 9445 11300 9455 11360
rect 9375 11250 9455 11300
rect 9375 11190 9385 11250
rect 9445 11190 9455 11250
rect 9375 11185 9455 11190
rect 9775 11360 9855 11365
rect 9775 11300 9785 11360
rect 9845 11300 9855 11360
rect 9775 11250 9855 11300
rect 9775 11190 9785 11250
rect 9845 11190 9855 11250
rect 9775 11185 9855 11190
rect 10175 11360 10255 11365
rect 10175 11300 10185 11360
rect 10245 11300 10255 11360
rect 10175 11250 10255 11300
rect 10175 11190 10185 11250
rect 10245 11190 10255 11250
rect 10175 11185 10255 11190
rect 10575 11360 10655 11365
rect 10575 11300 10585 11360
rect 10645 11300 10655 11360
rect 10575 11250 10655 11300
rect 10575 11190 10585 11250
rect 10645 11190 10655 11250
rect 10575 11185 10655 11190
rect 10975 11360 11055 11365
rect 10975 11300 10985 11360
rect 11045 11300 11055 11360
rect 10975 11250 11055 11300
rect 10975 11190 10985 11250
rect 11045 11190 11055 11250
rect 10975 11185 11055 11190
rect 11375 11360 11455 11365
rect 11375 11300 11385 11360
rect 11445 11300 11455 11360
rect 11375 11250 11455 11300
rect 11375 11190 11385 11250
rect 11445 11190 11455 11250
rect 11375 11185 11455 11190
rect 11775 11360 11855 11365
rect 11775 11300 11785 11360
rect 11845 11300 11855 11360
rect 11775 11250 11855 11300
rect 11775 11190 11785 11250
rect 11845 11190 11855 11250
rect 11775 11185 11855 11190
rect 12175 11360 12255 11365
rect 12175 11300 12185 11360
rect 12245 11300 12255 11360
rect 12175 11250 12255 11300
rect 12175 11190 12185 11250
rect 12245 11190 12255 11250
rect 12175 11185 12255 11190
rect 12575 11360 12655 11365
rect 12575 11300 12585 11360
rect 12645 11300 12655 11360
rect 12575 11250 12655 11300
rect 12575 11190 12585 11250
rect 12645 11190 12655 11250
rect 12575 11185 12655 11190
rect 12975 11360 13055 11365
rect 12975 11300 12985 11360
rect 13045 11300 13055 11360
rect 12975 11250 13055 11300
rect 12975 11190 12985 11250
rect 13045 11190 13055 11250
rect 12975 11185 13055 11190
rect -215 10995 -155 11185
rect 185 10995 245 11185
rect 585 10995 645 11185
rect 985 10995 1045 11185
rect 1385 10995 1445 11185
rect 1785 10995 1845 11185
rect 2185 10995 2245 11185
rect 2585 10995 2645 11185
rect 2985 10995 3045 11185
rect 3385 10995 3445 11185
rect 3785 10995 3845 11185
rect 4185 10995 4245 11185
rect 4585 10995 4645 11185
rect 4985 10995 5045 11185
rect 5385 10995 5445 11185
rect 5785 10995 5845 11185
rect 6185 10995 6245 11185
rect 6585 10995 6645 11185
rect 6985 10995 7045 11185
rect 7385 10995 7445 11185
rect 7785 10995 7845 11185
rect 8185 10995 8245 11185
rect 8585 10995 8645 11185
rect 8985 10995 9045 11185
rect 9385 10995 9445 11185
rect 9785 10995 9845 11185
rect 10185 10995 10245 11185
rect 10585 10995 10645 11185
rect 10985 10995 11045 11185
rect 11385 10995 11445 11185
rect 11785 10995 11845 11185
rect 12185 10995 12245 11185
rect 12585 10995 12645 11185
rect 12985 10995 13045 11185
rect -225 10990 -145 10995
rect -225 10930 -215 10990
rect -155 10930 -145 10990
rect -225 10880 -145 10930
rect -225 10820 -215 10880
rect -155 10820 -145 10880
rect -225 10815 -145 10820
rect 175 10990 255 10995
rect 175 10930 185 10990
rect 245 10930 255 10990
rect 175 10880 255 10930
rect 175 10820 185 10880
rect 245 10820 255 10880
rect 175 10815 255 10820
rect 575 10990 655 10995
rect 575 10930 585 10990
rect 645 10930 655 10990
rect 575 10880 655 10930
rect 575 10820 585 10880
rect 645 10820 655 10880
rect 575 10815 655 10820
rect 975 10990 1055 10995
rect 975 10930 985 10990
rect 1045 10930 1055 10990
rect 975 10880 1055 10930
rect 975 10820 985 10880
rect 1045 10820 1055 10880
rect 975 10815 1055 10820
rect 1375 10990 1455 10995
rect 1375 10930 1385 10990
rect 1445 10930 1455 10990
rect 1375 10880 1455 10930
rect 1375 10820 1385 10880
rect 1445 10820 1455 10880
rect 1375 10815 1455 10820
rect 1775 10990 1855 10995
rect 1775 10930 1785 10990
rect 1845 10930 1855 10990
rect 1775 10880 1855 10930
rect 1775 10820 1785 10880
rect 1845 10820 1855 10880
rect 1775 10815 1855 10820
rect 2175 10990 2255 10995
rect 2175 10930 2185 10990
rect 2245 10930 2255 10990
rect 2175 10880 2255 10930
rect 2175 10820 2185 10880
rect 2245 10820 2255 10880
rect 2175 10815 2255 10820
rect 2575 10990 2655 10995
rect 2575 10930 2585 10990
rect 2645 10930 2655 10990
rect 2575 10880 2655 10930
rect 2575 10820 2585 10880
rect 2645 10820 2655 10880
rect 2575 10815 2655 10820
rect 2975 10990 3055 10995
rect 2975 10930 2985 10990
rect 3045 10930 3055 10990
rect 2975 10880 3055 10930
rect 2975 10820 2985 10880
rect 3045 10820 3055 10880
rect 2975 10815 3055 10820
rect 3375 10990 3455 10995
rect 3375 10930 3385 10990
rect 3445 10930 3455 10990
rect 3375 10880 3455 10930
rect 3375 10820 3385 10880
rect 3445 10820 3455 10880
rect 3375 10815 3455 10820
rect 3775 10990 3855 10995
rect 3775 10930 3785 10990
rect 3845 10930 3855 10990
rect 3775 10880 3855 10930
rect 3775 10820 3785 10880
rect 3845 10820 3855 10880
rect 3775 10815 3855 10820
rect 4175 10990 4255 10995
rect 4175 10930 4185 10990
rect 4245 10930 4255 10990
rect 4175 10880 4255 10930
rect 4175 10820 4185 10880
rect 4245 10820 4255 10880
rect 4175 10815 4255 10820
rect 4575 10990 4655 10995
rect 4575 10930 4585 10990
rect 4645 10930 4655 10990
rect 4575 10880 4655 10930
rect 4575 10820 4585 10880
rect 4645 10820 4655 10880
rect 4575 10815 4655 10820
rect 4975 10990 5055 10995
rect 4975 10930 4985 10990
rect 5045 10930 5055 10990
rect 4975 10880 5055 10930
rect 4975 10820 4985 10880
rect 5045 10820 5055 10880
rect 4975 10815 5055 10820
rect 5375 10990 5455 10995
rect 5375 10930 5385 10990
rect 5445 10930 5455 10990
rect 5375 10880 5455 10930
rect 5375 10820 5385 10880
rect 5445 10820 5455 10880
rect 5375 10815 5455 10820
rect 5775 10990 5855 10995
rect 5775 10930 5785 10990
rect 5845 10930 5855 10990
rect 5775 10880 5855 10930
rect 5775 10820 5785 10880
rect 5845 10820 5855 10880
rect 5775 10815 5855 10820
rect 6175 10990 6255 10995
rect 6175 10930 6185 10990
rect 6245 10930 6255 10990
rect 6175 10880 6255 10930
rect 6175 10820 6185 10880
rect 6245 10820 6255 10880
rect 6175 10815 6255 10820
rect 6575 10990 6655 10995
rect 6575 10930 6585 10990
rect 6645 10930 6655 10990
rect 6575 10880 6655 10930
rect 6575 10820 6585 10880
rect 6645 10820 6655 10880
rect 6575 10815 6655 10820
rect 6975 10990 7055 10995
rect 6975 10930 6985 10990
rect 7045 10930 7055 10990
rect 6975 10880 7055 10930
rect 6975 10820 6985 10880
rect 7045 10820 7055 10880
rect 6975 10815 7055 10820
rect 7375 10990 7455 10995
rect 7375 10930 7385 10990
rect 7445 10930 7455 10990
rect 7375 10880 7455 10930
rect 7375 10820 7385 10880
rect 7445 10820 7455 10880
rect 7375 10815 7455 10820
rect 7775 10990 7855 10995
rect 7775 10930 7785 10990
rect 7845 10930 7855 10990
rect 7775 10880 7855 10930
rect 7775 10820 7785 10880
rect 7845 10820 7855 10880
rect 7775 10815 7855 10820
rect 8175 10990 8255 10995
rect 8175 10930 8185 10990
rect 8245 10930 8255 10990
rect 8175 10880 8255 10930
rect 8175 10820 8185 10880
rect 8245 10820 8255 10880
rect 8175 10815 8255 10820
rect 8575 10990 8655 10995
rect 8575 10930 8585 10990
rect 8645 10930 8655 10990
rect 8575 10880 8655 10930
rect 8575 10820 8585 10880
rect 8645 10820 8655 10880
rect 8575 10815 8655 10820
rect 8975 10990 9055 10995
rect 8975 10930 8985 10990
rect 9045 10930 9055 10990
rect 8975 10880 9055 10930
rect 8975 10820 8985 10880
rect 9045 10820 9055 10880
rect 8975 10815 9055 10820
rect 9375 10990 9455 10995
rect 9375 10930 9385 10990
rect 9445 10930 9455 10990
rect 9375 10880 9455 10930
rect 9375 10820 9385 10880
rect 9445 10820 9455 10880
rect 9375 10815 9455 10820
rect 9775 10990 9855 10995
rect 9775 10930 9785 10990
rect 9845 10930 9855 10990
rect 9775 10880 9855 10930
rect 9775 10820 9785 10880
rect 9845 10820 9855 10880
rect 9775 10815 9855 10820
rect 10175 10990 10255 10995
rect 10175 10930 10185 10990
rect 10245 10930 10255 10990
rect 10175 10880 10255 10930
rect 10175 10820 10185 10880
rect 10245 10820 10255 10880
rect 10175 10815 10255 10820
rect 10575 10990 10655 10995
rect 10575 10930 10585 10990
rect 10645 10930 10655 10990
rect 10575 10880 10655 10930
rect 10575 10820 10585 10880
rect 10645 10820 10655 10880
rect 10575 10815 10655 10820
rect 10975 10990 11055 10995
rect 10975 10930 10985 10990
rect 11045 10930 11055 10990
rect 10975 10880 11055 10930
rect 10975 10820 10985 10880
rect 11045 10820 11055 10880
rect 10975 10815 11055 10820
rect 11375 10990 11455 10995
rect 11375 10930 11385 10990
rect 11445 10930 11455 10990
rect 11375 10880 11455 10930
rect 11375 10820 11385 10880
rect 11445 10820 11455 10880
rect 11375 10815 11455 10820
rect 11775 10990 11855 10995
rect 11775 10930 11785 10990
rect 11845 10930 11855 10990
rect 11775 10880 11855 10930
rect 11775 10820 11785 10880
rect 11845 10820 11855 10880
rect 11775 10815 11855 10820
rect 12175 10990 12255 10995
rect 12175 10930 12185 10990
rect 12245 10930 12255 10990
rect 12175 10880 12255 10930
rect 12175 10820 12185 10880
rect 12245 10820 12255 10880
rect 12175 10815 12255 10820
rect 12575 10990 12655 10995
rect 12575 10930 12585 10990
rect 12645 10930 12655 10990
rect 12575 10880 12655 10930
rect 12575 10820 12585 10880
rect 12645 10820 12655 10880
rect 12575 10815 12655 10820
rect 12975 10990 13055 10995
rect 12975 10930 12985 10990
rect 13045 10930 13055 10990
rect 12975 10880 13055 10930
rect 12975 10820 12985 10880
rect 13045 10820 13055 10880
rect 12975 10815 13055 10820
rect -215 10625 -155 10815
rect 185 10625 245 10815
rect 585 10625 645 10815
rect 985 10625 1045 10815
rect 1385 10625 1445 10815
rect 1785 10625 1845 10815
rect 2185 10625 2245 10815
rect 2585 10625 2645 10815
rect 2985 10625 3045 10815
rect 3385 10625 3445 10815
rect 3785 10625 3845 10815
rect 4185 10625 4245 10815
rect 4585 10625 4645 10815
rect 4985 10625 5045 10815
rect 5385 10625 5445 10815
rect 5785 10625 5845 10815
rect 6185 10625 6245 10815
rect 6585 10625 6645 10815
rect 6985 10625 7045 10815
rect 7385 10625 7445 10815
rect 7785 10625 7845 10815
rect 8185 10625 8245 10815
rect 8585 10625 8645 10815
rect 8985 10625 9045 10815
rect 9385 10625 9445 10815
rect 9785 10625 9845 10815
rect 10185 10625 10245 10815
rect 10585 10625 10645 10815
rect 10985 10625 11045 10815
rect 11385 10625 11445 10815
rect 11785 10625 11845 10815
rect 12185 10625 12245 10815
rect 12585 10625 12645 10815
rect 12985 10625 13045 10815
rect -225 10620 -145 10625
rect -225 10560 -215 10620
rect -155 10560 -145 10620
rect -225 10510 -145 10560
rect -225 10450 -215 10510
rect -155 10450 -145 10510
rect -225 10445 -145 10450
rect 175 10620 255 10625
rect 175 10560 185 10620
rect 245 10560 255 10620
rect 175 10510 255 10560
rect 175 10450 185 10510
rect 245 10450 255 10510
rect 175 10445 255 10450
rect 575 10620 655 10625
rect 575 10560 585 10620
rect 645 10560 655 10620
rect 575 10510 655 10560
rect 575 10450 585 10510
rect 645 10450 655 10510
rect 575 10445 655 10450
rect 975 10620 1055 10625
rect 975 10560 985 10620
rect 1045 10560 1055 10620
rect 975 10510 1055 10560
rect 975 10450 985 10510
rect 1045 10450 1055 10510
rect 975 10445 1055 10450
rect 1375 10620 1455 10625
rect 1375 10560 1385 10620
rect 1445 10560 1455 10620
rect 1375 10510 1455 10560
rect 1375 10450 1385 10510
rect 1445 10450 1455 10510
rect 1375 10445 1455 10450
rect 1775 10620 1855 10625
rect 1775 10560 1785 10620
rect 1845 10560 1855 10620
rect 1775 10510 1855 10560
rect 1775 10450 1785 10510
rect 1845 10450 1855 10510
rect 1775 10445 1855 10450
rect 2175 10620 2255 10625
rect 2175 10560 2185 10620
rect 2245 10560 2255 10620
rect 2175 10510 2255 10560
rect 2175 10450 2185 10510
rect 2245 10450 2255 10510
rect 2175 10445 2255 10450
rect 2575 10620 2655 10625
rect 2575 10560 2585 10620
rect 2645 10560 2655 10620
rect 2575 10510 2655 10560
rect 2575 10450 2585 10510
rect 2645 10450 2655 10510
rect 2575 10445 2655 10450
rect 2975 10620 3055 10625
rect 2975 10560 2985 10620
rect 3045 10560 3055 10620
rect 2975 10510 3055 10560
rect 2975 10450 2985 10510
rect 3045 10450 3055 10510
rect 2975 10445 3055 10450
rect 3375 10620 3455 10625
rect 3375 10560 3385 10620
rect 3445 10560 3455 10620
rect 3375 10510 3455 10560
rect 3375 10450 3385 10510
rect 3445 10450 3455 10510
rect 3375 10445 3455 10450
rect 3775 10620 3855 10625
rect 3775 10560 3785 10620
rect 3845 10560 3855 10620
rect 3775 10510 3855 10560
rect 3775 10450 3785 10510
rect 3845 10450 3855 10510
rect 3775 10445 3855 10450
rect 4175 10620 4255 10625
rect 4175 10560 4185 10620
rect 4245 10560 4255 10620
rect 4175 10510 4255 10560
rect 4175 10450 4185 10510
rect 4245 10450 4255 10510
rect 4175 10445 4255 10450
rect 4575 10620 4655 10625
rect 4575 10560 4585 10620
rect 4645 10560 4655 10620
rect 4575 10510 4655 10560
rect 4575 10450 4585 10510
rect 4645 10450 4655 10510
rect 4575 10445 4655 10450
rect 4975 10620 5055 10625
rect 4975 10560 4985 10620
rect 5045 10560 5055 10620
rect 4975 10510 5055 10560
rect 4975 10450 4985 10510
rect 5045 10450 5055 10510
rect 4975 10445 5055 10450
rect 5375 10620 5455 10625
rect 5375 10560 5385 10620
rect 5445 10560 5455 10620
rect 5375 10510 5455 10560
rect 5375 10450 5385 10510
rect 5445 10450 5455 10510
rect 5375 10445 5455 10450
rect 5775 10620 5855 10625
rect 5775 10560 5785 10620
rect 5845 10560 5855 10620
rect 5775 10510 5855 10560
rect 5775 10450 5785 10510
rect 5845 10450 5855 10510
rect 5775 10445 5855 10450
rect 6175 10620 6255 10625
rect 6175 10560 6185 10620
rect 6245 10560 6255 10620
rect 6175 10510 6255 10560
rect 6175 10450 6185 10510
rect 6245 10450 6255 10510
rect 6175 10445 6255 10450
rect 6575 10620 6655 10625
rect 6575 10560 6585 10620
rect 6645 10560 6655 10620
rect 6575 10510 6655 10560
rect 6575 10450 6585 10510
rect 6645 10450 6655 10510
rect 6575 10445 6655 10450
rect 6975 10620 7055 10625
rect 6975 10560 6985 10620
rect 7045 10560 7055 10620
rect 6975 10510 7055 10560
rect 6975 10450 6985 10510
rect 7045 10450 7055 10510
rect 6975 10445 7055 10450
rect 7375 10620 7455 10625
rect 7375 10560 7385 10620
rect 7445 10560 7455 10620
rect 7375 10510 7455 10560
rect 7375 10450 7385 10510
rect 7445 10450 7455 10510
rect 7375 10445 7455 10450
rect 7775 10620 7855 10625
rect 7775 10560 7785 10620
rect 7845 10560 7855 10620
rect 7775 10510 7855 10560
rect 7775 10450 7785 10510
rect 7845 10450 7855 10510
rect 7775 10445 7855 10450
rect 8175 10620 8255 10625
rect 8175 10560 8185 10620
rect 8245 10560 8255 10620
rect 8175 10510 8255 10560
rect 8175 10450 8185 10510
rect 8245 10450 8255 10510
rect 8175 10445 8255 10450
rect 8575 10620 8655 10625
rect 8575 10560 8585 10620
rect 8645 10560 8655 10620
rect 8575 10510 8655 10560
rect 8575 10450 8585 10510
rect 8645 10450 8655 10510
rect 8575 10445 8655 10450
rect 8975 10620 9055 10625
rect 8975 10560 8985 10620
rect 9045 10560 9055 10620
rect 8975 10510 9055 10560
rect 8975 10450 8985 10510
rect 9045 10450 9055 10510
rect 8975 10445 9055 10450
rect 9375 10620 9455 10625
rect 9375 10560 9385 10620
rect 9445 10560 9455 10620
rect 9375 10510 9455 10560
rect 9375 10450 9385 10510
rect 9445 10450 9455 10510
rect 9375 10445 9455 10450
rect 9775 10620 9855 10625
rect 9775 10560 9785 10620
rect 9845 10560 9855 10620
rect 9775 10510 9855 10560
rect 9775 10450 9785 10510
rect 9845 10450 9855 10510
rect 9775 10445 9855 10450
rect 10175 10620 10255 10625
rect 10175 10560 10185 10620
rect 10245 10560 10255 10620
rect 10175 10510 10255 10560
rect 10175 10450 10185 10510
rect 10245 10450 10255 10510
rect 10175 10445 10255 10450
rect 10575 10620 10655 10625
rect 10575 10560 10585 10620
rect 10645 10560 10655 10620
rect 10575 10510 10655 10560
rect 10575 10450 10585 10510
rect 10645 10450 10655 10510
rect 10575 10445 10655 10450
rect 10975 10620 11055 10625
rect 10975 10560 10985 10620
rect 11045 10560 11055 10620
rect 10975 10510 11055 10560
rect 10975 10450 10985 10510
rect 11045 10450 11055 10510
rect 10975 10445 11055 10450
rect 11375 10620 11455 10625
rect 11375 10560 11385 10620
rect 11445 10560 11455 10620
rect 11375 10510 11455 10560
rect 11375 10450 11385 10510
rect 11445 10450 11455 10510
rect 11375 10445 11455 10450
rect 11775 10620 11855 10625
rect 11775 10560 11785 10620
rect 11845 10560 11855 10620
rect 11775 10510 11855 10560
rect 11775 10450 11785 10510
rect 11845 10450 11855 10510
rect 11775 10445 11855 10450
rect 12175 10620 12255 10625
rect 12175 10560 12185 10620
rect 12245 10560 12255 10620
rect 12175 10510 12255 10560
rect 12175 10450 12185 10510
rect 12245 10450 12255 10510
rect 12175 10445 12255 10450
rect 12575 10620 12655 10625
rect 12575 10560 12585 10620
rect 12645 10560 12655 10620
rect 12575 10510 12655 10560
rect 12575 10450 12585 10510
rect 12645 10450 12655 10510
rect 12575 10445 12655 10450
rect 12975 10620 13055 10625
rect 12975 10560 12985 10620
rect 13045 10560 13055 10620
rect 12975 10510 13055 10560
rect 12975 10450 12985 10510
rect 13045 10450 13055 10510
rect 12975 10445 13055 10450
rect -215 10255 -155 10445
rect 185 10255 245 10445
rect 585 10255 645 10445
rect 985 10255 1045 10445
rect 1385 10255 1445 10445
rect 1785 10255 1845 10445
rect 2185 10255 2245 10445
rect 2585 10255 2645 10445
rect 2985 10255 3045 10445
rect 3385 10255 3445 10445
rect 3785 10255 3845 10445
rect 4185 10255 4245 10445
rect 4585 10255 4645 10445
rect 4985 10255 5045 10445
rect 5385 10255 5445 10445
rect 5785 10255 5845 10445
rect 6185 10255 6245 10445
rect 6585 10255 6645 10445
rect 6985 10255 7045 10445
rect 7385 10255 7445 10445
rect 7785 10255 7845 10445
rect 8185 10255 8245 10445
rect 8585 10255 8645 10445
rect 8985 10255 9045 10445
rect 9385 10255 9445 10445
rect 9785 10255 9845 10445
rect 10185 10255 10245 10445
rect 10585 10255 10645 10445
rect 10985 10255 11045 10445
rect 11385 10255 11445 10445
rect 11785 10255 11845 10445
rect 12185 10255 12245 10445
rect 12585 10255 12645 10445
rect 12985 10255 13045 10445
rect -225 10250 -145 10255
rect -225 10190 -215 10250
rect -155 10190 -145 10250
rect -225 10140 -145 10190
rect -225 10080 -215 10140
rect -155 10080 -145 10140
rect -225 10075 -145 10080
rect 175 10250 255 10255
rect 175 10190 185 10250
rect 245 10190 255 10250
rect 175 10140 255 10190
rect 175 10080 185 10140
rect 245 10080 255 10140
rect 175 10075 255 10080
rect 575 10250 655 10255
rect 575 10190 585 10250
rect 645 10190 655 10250
rect 575 10140 655 10190
rect 575 10080 585 10140
rect 645 10080 655 10140
rect 575 10075 655 10080
rect 975 10250 1055 10255
rect 975 10190 985 10250
rect 1045 10190 1055 10250
rect 975 10140 1055 10190
rect 975 10080 985 10140
rect 1045 10080 1055 10140
rect 975 10075 1055 10080
rect 1375 10250 1455 10255
rect 1375 10190 1385 10250
rect 1445 10190 1455 10250
rect 1375 10140 1455 10190
rect 1375 10080 1385 10140
rect 1445 10080 1455 10140
rect 1375 10075 1455 10080
rect 1775 10250 1855 10255
rect 1775 10190 1785 10250
rect 1845 10190 1855 10250
rect 1775 10140 1855 10190
rect 1775 10080 1785 10140
rect 1845 10080 1855 10140
rect 1775 10075 1855 10080
rect 2175 10250 2255 10255
rect 2175 10190 2185 10250
rect 2245 10190 2255 10250
rect 2175 10140 2255 10190
rect 2175 10080 2185 10140
rect 2245 10080 2255 10140
rect 2175 10075 2255 10080
rect 2575 10250 2655 10255
rect 2575 10190 2585 10250
rect 2645 10190 2655 10250
rect 2575 10140 2655 10190
rect 2575 10080 2585 10140
rect 2645 10080 2655 10140
rect 2575 10075 2655 10080
rect 2975 10250 3055 10255
rect 2975 10190 2985 10250
rect 3045 10190 3055 10250
rect 2975 10140 3055 10190
rect 2975 10080 2985 10140
rect 3045 10080 3055 10140
rect 2975 10075 3055 10080
rect 3375 10250 3455 10255
rect 3375 10190 3385 10250
rect 3445 10190 3455 10250
rect 3375 10140 3455 10190
rect 3375 10080 3385 10140
rect 3445 10080 3455 10140
rect 3375 10075 3455 10080
rect 3775 10250 3855 10255
rect 3775 10190 3785 10250
rect 3845 10190 3855 10250
rect 3775 10140 3855 10190
rect 3775 10080 3785 10140
rect 3845 10080 3855 10140
rect 3775 10075 3855 10080
rect 4175 10250 4255 10255
rect 4175 10190 4185 10250
rect 4245 10190 4255 10250
rect 4175 10140 4255 10190
rect 4175 10080 4185 10140
rect 4245 10080 4255 10140
rect 4175 10075 4255 10080
rect 4575 10250 4655 10255
rect 4575 10190 4585 10250
rect 4645 10190 4655 10250
rect 4575 10140 4655 10190
rect 4575 10080 4585 10140
rect 4645 10080 4655 10140
rect 4575 10075 4655 10080
rect 4975 10250 5055 10255
rect 4975 10190 4985 10250
rect 5045 10190 5055 10250
rect 4975 10140 5055 10190
rect 4975 10080 4985 10140
rect 5045 10080 5055 10140
rect 4975 10075 5055 10080
rect 5375 10250 5455 10255
rect 5375 10190 5385 10250
rect 5445 10190 5455 10250
rect 5375 10140 5455 10190
rect 5375 10080 5385 10140
rect 5445 10080 5455 10140
rect 5375 10075 5455 10080
rect 5775 10250 5855 10255
rect 5775 10190 5785 10250
rect 5845 10190 5855 10250
rect 5775 10140 5855 10190
rect 5775 10080 5785 10140
rect 5845 10080 5855 10140
rect 5775 10075 5855 10080
rect 6175 10250 6255 10255
rect 6175 10190 6185 10250
rect 6245 10190 6255 10250
rect 6175 10140 6255 10190
rect 6175 10080 6185 10140
rect 6245 10080 6255 10140
rect 6175 10075 6255 10080
rect 6575 10250 6655 10255
rect 6575 10190 6585 10250
rect 6645 10190 6655 10250
rect 6575 10140 6655 10190
rect 6575 10080 6585 10140
rect 6645 10080 6655 10140
rect 6575 10075 6655 10080
rect 6975 10250 7055 10255
rect 6975 10190 6985 10250
rect 7045 10190 7055 10250
rect 6975 10140 7055 10190
rect 6975 10080 6985 10140
rect 7045 10080 7055 10140
rect 6975 10075 7055 10080
rect 7375 10250 7455 10255
rect 7375 10190 7385 10250
rect 7445 10190 7455 10250
rect 7375 10140 7455 10190
rect 7375 10080 7385 10140
rect 7445 10080 7455 10140
rect 7375 10075 7455 10080
rect 7775 10250 7855 10255
rect 7775 10190 7785 10250
rect 7845 10190 7855 10250
rect 7775 10140 7855 10190
rect 7775 10080 7785 10140
rect 7845 10080 7855 10140
rect 7775 10075 7855 10080
rect 8175 10250 8255 10255
rect 8175 10190 8185 10250
rect 8245 10190 8255 10250
rect 8175 10140 8255 10190
rect 8175 10080 8185 10140
rect 8245 10080 8255 10140
rect 8175 10075 8255 10080
rect 8575 10250 8655 10255
rect 8575 10190 8585 10250
rect 8645 10190 8655 10250
rect 8575 10140 8655 10190
rect 8575 10080 8585 10140
rect 8645 10080 8655 10140
rect 8575 10075 8655 10080
rect 8975 10250 9055 10255
rect 8975 10190 8985 10250
rect 9045 10190 9055 10250
rect 8975 10140 9055 10190
rect 8975 10080 8985 10140
rect 9045 10080 9055 10140
rect 8975 10075 9055 10080
rect 9375 10250 9455 10255
rect 9375 10190 9385 10250
rect 9445 10190 9455 10250
rect 9375 10140 9455 10190
rect 9375 10080 9385 10140
rect 9445 10080 9455 10140
rect 9375 10075 9455 10080
rect 9775 10250 9855 10255
rect 9775 10190 9785 10250
rect 9845 10190 9855 10250
rect 9775 10140 9855 10190
rect 9775 10080 9785 10140
rect 9845 10080 9855 10140
rect 9775 10075 9855 10080
rect 10175 10250 10255 10255
rect 10175 10190 10185 10250
rect 10245 10190 10255 10250
rect 10175 10140 10255 10190
rect 10175 10080 10185 10140
rect 10245 10080 10255 10140
rect 10175 10075 10255 10080
rect 10575 10250 10655 10255
rect 10575 10190 10585 10250
rect 10645 10190 10655 10250
rect 10575 10140 10655 10190
rect 10575 10080 10585 10140
rect 10645 10080 10655 10140
rect 10575 10075 10655 10080
rect 10975 10250 11055 10255
rect 10975 10190 10985 10250
rect 11045 10190 11055 10250
rect 10975 10140 11055 10190
rect 10975 10080 10985 10140
rect 11045 10080 11055 10140
rect 10975 10075 11055 10080
rect 11375 10250 11455 10255
rect 11375 10190 11385 10250
rect 11445 10190 11455 10250
rect 11375 10140 11455 10190
rect 11375 10080 11385 10140
rect 11445 10080 11455 10140
rect 11375 10075 11455 10080
rect 11775 10250 11855 10255
rect 11775 10190 11785 10250
rect 11845 10190 11855 10250
rect 11775 10140 11855 10190
rect 11775 10080 11785 10140
rect 11845 10080 11855 10140
rect 11775 10075 11855 10080
rect 12175 10250 12255 10255
rect 12175 10190 12185 10250
rect 12245 10190 12255 10250
rect 12175 10140 12255 10190
rect 12175 10080 12185 10140
rect 12245 10080 12255 10140
rect 12175 10075 12255 10080
rect 12575 10250 12655 10255
rect 12575 10190 12585 10250
rect 12645 10190 12655 10250
rect 12575 10140 12655 10190
rect 12575 10080 12585 10140
rect 12645 10080 12655 10140
rect 12575 10075 12655 10080
rect 12975 10250 13055 10255
rect 12975 10190 12985 10250
rect 13045 10190 13055 10250
rect 12975 10140 13055 10190
rect 12975 10080 12985 10140
rect 13045 10080 13055 10140
rect 12975 10075 13055 10080
rect -215 9885 -155 10075
rect 185 9885 245 10075
rect 585 9885 645 10075
rect 985 9885 1045 10075
rect 1385 9885 1445 10075
rect 1785 9885 1845 10075
rect 2185 9885 2245 10075
rect 2585 9885 2645 10075
rect 2985 9885 3045 10075
rect 3385 9885 3445 10075
rect 3785 9885 3845 10075
rect 4185 9885 4245 10075
rect 4585 9885 4645 10075
rect 4985 9885 5045 10075
rect 5385 9885 5445 10075
rect 5785 9885 5845 10075
rect 6185 9885 6245 10075
rect 6585 9885 6645 10075
rect 6985 9885 7045 10075
rect 7385 9885 7445 10075
rect 7785 9885 7845 10075
rect 8185 9885 8245 10075
rect 8585 9885 8645 10075
rect 8985 9885 9045 10075
rect 9385 9885 9445 10075
rect 9785 9885 9845 10075
rect 10185 9885 10245 10075
rect 10585 9885 10645 10075
rect 10985 9885 11045 10075
rect 11385 9885 11445 10075
rect 11785 9885 11845 10075
rect 12185 9885 12245 10075
rect 12585 9885 12645 10075
rect 12985 9885 13045 10075
rect -225 9880 -145 9885
rect -225 9820 -215 9880
rect -155 9820 -145 9880
rect -225 9770 -145 9820
rect -225 9710 -215 9770
rect -155 9710 -145 9770
rect -225 9705 -145 9710
rect 175 9880 255 9885
rect 175 9820 185 9880
rect 245 9820 255 9880
rect 175 9770 255 9820
rect 175 9710 185 9770
rect 245 9710 255 9770
rect 175 9705 255 9710
rect 575 9880 655 9885
rect 575 9820 585 9880
rect 645 9820 655 9880
rect 575 9770 655 9820
rect 575 9710 585 9770
rect 645 9710 655 9770
rect 575 9705 655 9710
rect 975 9880 1055 9885
rect 975 9820 985 9880
rect 1045 9820 1055 9880
rect 975 9770 1055 9820
rect 975 9710 985 9770
rect 1045 9710 1055 9770
rect 975 9705 1055 9710
rect 1375 9880 1455 9885
rect 1375 9820 1385 9880
rect 1445 9820 1455 9880
rect 1375 9770 1455 9820
rect 1375 9710 1385 9770
rect 1445 9710 1455 9770
rect 1375 9705 1455 9710
rect 1775 9880 1855 9885
rect 1775 9820 1785 9880
rect 1845 9820 1855 9880
rect 1775 9770 1855 9820
rect 1775 9710 1785 9770
rect 1845 9710 1855 9770
rect 1775 9705 1855 9710
rect 2175 9880 2255 9885
rect 2175 9820 2185 9880
rect 2245 9820 2255 9880
rect 2175 9770 2255 9820
rect 2175 9710 2185 9770
rect 2245 9710 2255 9770
rect 2175 9705 2255 9710
rect 2575 9880 2655 9885
rect 2575 9820 2585 9880
rect 2645 9820 2655 9880
rect 2575 9770 2655 9820
rect 2575 9710 2585 9770
rect 2645 9710 2655 9770
rect 2575 9705 2655 9710
rect 2975 9880 3055 9885
rect 2975 9820 2985 9880
rect 3045 9820 3055 9880
rect 2975 9770 3055 9820
rect 2975 9710 2985 9770
rect 3045 9710 3055 9770
rect 2975 9705 3055 9710
rect 3375 9880 3455 9885
rect 3375 9820 3385 9880
rect 3445 9820 3455 9880
rect 3375 9770 3455 9820
rect 3375 9710 3385 9770
rect 3445 9710 3455 9770
rect 3375 9705 3455 9710
rect 3775 9880 3855 9885
rect 3775 9820 3785 9880
rect 3845 9820 3855 9880
rect 3775 9770 3855 9820
rect 3775 9710 3785 9770
rect 3845 9710 3855 9770
rect 3775 9705 3855 9710
rect 4175 9880 4255 9885
rect 4175 9820 4185 9880
rect 4245 9820 4255 9880
rect 4175 9770 4255 9820
rect 4175 9710 4185 9770
rect 4245 9710 4255 9770
rect 4175 9705 4255 9710
rect 4575 9880 4655 9885
rect 4575 9820 4585 9880
rect 4645 9820 4655 9880
rect 4575 9770 4655 9820
rect 4575 9710 4585 9770
rect 4645 9710 4655 9770
rect 4575 9705 4655 9710
rect 4975 9880 5055 9885
rect 4975 9820 4985 9880
rect 5045 9820 5055 9880
rect 4975 9770 5055 9820
rect 4975 9710 4985 9770
rect 5045 9710 5055 9770
rect 4975 9705 5055 9710
rect 5375 9880 5455 9885
rect 5375 9820 5385 9880
rect 5445 9820 5455 9880
rect 5375 9770 5455 9820
rect 5375 9710 5385 9770
rect 5445 9710 5455 9770
rect 5375 9705 5455 9710
rect 5775 9880 5855 9885
rect 5775 9820 5785 9880
rect 5845 9820 5855 9880
rect 5775 9770 5855 9820
rect 5775 9710 5785 9770
rect 5845 9710 5855 9770
rect 5775 9705 5855 9710
rect 6175 9880 6255 9885
rect 6175 9820 6185 9880
rect 6245 9820 6255 9880
rect 6175 9770 6255 9820
rect 6175 9710 6185 9770
rect 6245 9710 6255 9770
rect 6175 9705 6255 9710
rect 6575 9880 6655 9885
rect 6575 9820 6585 9880
rect 6645 9820 6655 9880
rect 6575 9770 6655 9820
rect 6575 9710 6585 9770
rect 6645 9710 6655 9770
rect 6575 9705 6655 9710
rect 6975 9880 7055 9885
rect 6975 9820 6985 9880
rect 7045 9820 7055 9880
rect 6975 9770 7055 9820
rect 6975 9710 6985 9770
rect 7045 9710 7055 9770
rect 6975 9705 7055 9710
rect 7375 9880 7455 9885
rect 7375 9820 7385 9880
rect 7445 9820 7455 9880
rect 7375 9770 7455 9820
rect 7375 9710 7385 9770
rect 7445 9710 7455 9770
rect 7375 9705 7455 9710
rect 7775 9880 7855 9885
rect 7775 9820 7785 9880
rect 7845 9820 7855 9880
rect 7775 9770 7855 9820
rect 7775 9710 7785 9770
rect 7845 9710 7855 9770
rect 7775 9705 7855 9710
rect 8175 9880 8255 9885
rect 8175 9820 8185 9880
rect 8245 9820 8255 9880
rect 8175 9770 8255 9820
rect 8175 9710 8185 9770
rect 8245 9710 8255 9770
rect 8175 9705 8255 9710
rect 8575 9880 8655 9885
rect 8575 9820 8585 9880
rect 8645 9820 8655 9880
rect 8575 9770 8655 9820
rect 8575 9710 8585 9770
rect 8645 9710 8655 9770
rect 8575 9705 8655 9710
rect 8975 9880 9055 9885
rect 8975 9820 8985 9880
rect 9045 9820 9055 9880
rect 8975 9770 9055 9820
rect 8975 9710 8985 9770
rect 9045 9710 9055 9770
rect 8975 9705 9055 9710
rect 9375 9880 9455 9885
rect 9375 9820 9385 9880
rect 9445 9820 9455 9880
rect 9375 9770 9455 9820
rect 9375 9710 9385 9770
rect 9445 9710 9455 9770
rect 9375 9705 9455 9710
rect 9775 9880 9855 9885
rect 9775 9820 9785 9880
rect 9845 9820 9855 9880
rect 9775 9770 9855 9820
rect 9775 9710 9785 9770
rect 9845 9710 9855 9770
rect 9775 9705 9855 9710
rect 10175 9880 10255 9885
rect 10175 9820 10185 9880
rect 10245 9820 10255 9880
rect 10175 9770 10255 9820
rect 10175 9710 10185 9770
rect 10245 9710 10255 9770
rect 10175 9705 10255 9710
rect 10575 9880 10655 9885
rect 10575 9820 10585 9880
rect 10645 9820 10655 9880
rect 10575 9770 10655 9820
rect 10575 9710 10585 9770
rect 10645 9710 10655 9770
rect 10575 9705 10655 9710
rect 10975 9880 11055 9885
rect 10975 9820 10985 9880
rect 11045 9820 11055 9880
rect 10975 9770 11055 9820
rect 10975 9710 10985 9770
rect 11045 9710 11055 9770
rect 10975 9705 11055 9710
rect 11375 9880 11455 9885
rect 11375 9820 11385 9880
rect 11445 9820 11455 9880
rect 11375 9770 11455 9820
rect 11375 9710 11385 9770
rect 11445 9710 11455 9770
rect 11375 9705 11455 9710
rect 11775 9880 11855 9885
rect 11775 9820 11785 9880
rect 11845 9820 11855 9880
rect 11775 9770 11855 9820
rect 11775 9710 11785 9770
rect 11845 9710 11855 9770
rect 11775 9705 11855 9710
rect 12175 9880 12255 9885
rect 12175 9820 12185 9880
rect 12245 9820 12255 9880
rect 12175 9770 12255 9820
rect 12175 9710 12185 9770
rect 12245 9710 12255 9770
rect 12175 9705 12255 9710
rect 12575 9880 12655 9885
rect 12575 9820 12585 9880
rect 12645 9820 12655 9880
rect 12575 9770 12655 9820
rect 12575 9710 12585 9770
rect 12645 9710 12655 9770
rect 12575 9705 12655 9710
rect 12975 9880 13055 9885
rect 12975 9820 12985 9880
rect 13045 9820 13055 9880
rect 12975 9770 13055 9820
rect 12975 9710 12985 9770
rect 13045 9710 13055 9770
rect 12975 9705 13055 9710
rect -215 9515 -155 9705
rect 185 9515 245 9705
rect 585 9515 645 9705
rect 985 9515 1045 9705
rect 1385 9515 1445 9705
rect 1785 9515 1845 9705
rect 2185 9515 2245 9705
rect 2585 9515 2645 9705
rect 2985 9515 3045 9705
rect 3385 9515 3445 9705
rect 3785 9515 3845 9705
rect 4185 9515 4245 9705
rect 4585 9515 4645 9705
rect 4985 9515 5045 9705
rect 5385 9515 5445 9705
rect 5785 9515 5845 9705
rect 6185 9515 6245 9705
rect 6585 9515 6645 9705
rect 6985 9515 7045 9705
rect 7385 9515 7445 9705
rect 7785 9515 7845 9705
rect 8185 9515 8245 9705
rect 8585 9515 8645 9705
rect 8985 9515 9045 9705
rect 9385 9515 9445 9705
rect 9785 9515 9845 9705
rect 10185 9515 10245 9705
rect 10585 9515 10645 9705
rect 10985 9515 11045 9705
rect 11385 9515 11445 9705
rect 11785 9515 11845 9705
rect 12185 9515 12245 9705
rect 12585 9515 12645 9705
rect 12985 9515 13045 9705
rect -225 9510 -145 9515
rect -225 9450 -215 9510
rect -155 9450 -145 9510
rect -225 9400 -145 9450
rect -225 9340 -215 9400
rect -155 9340 -145 9400
rect -225 9335 -145 9340
rect 175 9510 255 9515
rect 175 9450 185 9510
rect 245 9450 255 9510
rect 175 9400 255 9450
rect 175 9340 185 9400
rect 245 9340 255 9400
rect 175 9335 255 9340
rect 575 9510 655 9515
rect 575 9450 585 9510
rect 645 9450 655 9510
rect 575 9400 655 9450
rect 575 9340 585 9400
rect 645 9340 655 9400
rect 575 9335 655 9340
rect 975 9510 1055 9515
rect 975 9450 985 9510
rect 1045 9450 1055 9510
rect 975 9400 1055 9450
rect 975 9340 985 9400
rect 1045 9340 1055 9400
rect 975 9335 1055 9340
rect 1375 9510 1455 9515
rect 1375 9450 1385 9510
rect 1445 9450 1455 9510
rect 1375 9400 1455 9450
rect 1375 9340 1385 9400
rect 1445 9340 1455 9400
rect 1375 9335 1455 9340
rect 1775 9510 1855 9515
rect 1775 9450 1785 9510
rect 1845 9450 1855 9510
rect 1775 9400 1855 9450
rect 1775 9340 1785 9400
rect 1845 9340 1855 9400
rect 1775 9335 1855 9340
rect 2175 9510 2255 9515
rect 2175 9450 2185 9510
rect 2245 9450 2255 9510
rect 2175 9400 2255 9450
rect 2175 9340 2185 9400
rect 2245 9340 2255 9400
rect 2175 9335 2255 9340
rect 2575 9510 2655 9515
rect 2575 9450 2585 9510
rect 2645 9450 2655 9510
rect 2575 9400 2655 9450
rect 2575 9340 2585 9400
rect 2645 9340 2655 9400
rect 2575 9335 2655 9340
rect 2975 9510 3055 9515
rect 2975 9450 2985 9510
rect 3045 9450 3055 9510
rect 2975 9400 3055 9450
rect 2975 9340 2985 9400
rect 3045 9340 3055 9400
rect 2975 9335 3055 9340
rect 3375 9510 3455 9515
rect 3375 9450 3385 9510
rect 3445 9450 3455 9510
rect 3375 9400 3455 9450
rect 3375 9340 3385 9400
rect 3445 9340 3455 9400
rect 3375 9335 3455 9340
rect 3775 9510 3855 9515
rect 3775 9450 3785 9510
rect 3845 9450 3855 9510
rect 3775 9400 3855 9450
rect 3775 9340 3785 9400
rect 3845 9340 3855 9400
rect 3775 9335 3855 9340
rect 4175 9510 4255 9515
rect 4175 9450 4185 9510
rect 4245 9450 4255 9510
rect 4175 9400 4255 9450
rect 4175 9340 4185 9400
rect 4245 9340 4255 9400
rect 4175 9335 4255 9340
rect 4575 9510 4655 9515
rect 4575 9450 4585 9510
rect 4645 9450 4655 9510
rect 4575 9400 4655 9450
rect 4575 9340 4585 9400
rect 4645 9340 4655 9400
rect 4575 9335 4655 9340
rect 4975 9510 5055 9515
rect 4975 9450 4985 9510
rect 5045 9450 5055 9510
rect 4975 9400 5055 9450
rect 4975 9340 4985 9400
rect 5045 9340 5055 9400
rect 4975 9335 5055 9340
rect 5375 9510 5455 9515
rect 5375 9450 5385 9510
rect 5445 9450 5455 9510
rect 5375 9400 5455 9450
rect 5375 9340 5385 9400
rect 5445 9340 5455 9400
rect 5375 9335 5455 9340
rect 5775 9510 5855 9515
rect 5775 9450 5785 9510
rect 5845 9450 5855 9510
rect 5775 9400 5855 9450
rect 5775 9340 5785 9400
rect 5845 9340 5855 9400
rect 5775 9335 5855 9340
rect 6175 9510 6255 9515
rect 6175 9450 6185 9510
rect 6245 9450 6255 9510
rect 6175 9400 6255 9450
rect 6175 9340 6185 9400
rect 6245 9340 6255 9400
rect 6175 9335 6255 9340
rect 6575 9510 6655 9515
rect 6575 9450 6585 9510
rect 6645 9450 6655 9510
rect 6575 9400 6655 9450
rect 6575 9340 6585 9400
rect 6645 9340 6655 9400
rect 6575 9335 6655 9340
rect 6975 9510 7055 9515
rect 6975 9450 6985 9510
rect 7045 9450 7055 9510
rect 6975 9400 7055 9450
rect 6975 9340 6985 9400
rect 7045 9340 7055 9400
rect 6975 9335 7055 9340
rect 7375 9510 7455 9515
rect 7375 9450 7385 9510
rect 7445 9450 7455 9510
rect 7375 9400 7455 9450
rect 7375 9340 7385 9400
rect 7445 9340 7455 9400
rect 7375 9335 7455 9340
rect 7775 9510 7855 9515
rect 7775 9450 7785 9510
rect 7845 9450 7855 9510
rect 7775 9400 7855 9450
rect 7775 9340 7785 9400
rect 7845 9340 7855 9400
rect 7775 9335 7855 9340
rect 8175 9510 8255 9515
rect 8175 9450 8185 9510
rect 8245 9450 8255 9510
rect 8175 9400 8255 9450
rect 8175 9340 8185 9400
rect 8245 9340 8255 9400
rect 8175 9335 8255 9340
rect 8575 9510 8655 9515
rect 8575 9450 8585 9510
rect 8645 9450 8655 9510
rect 8575 9400 8655 9450
rect 8575 9340 8585 9400
rect 8645 9340 8655 9400
rect 8575 9335 8655 9340
rect 8975 9510 9055 9515
rect 8975 9450 8985 9510
rect 9045 9450 9055 9510
rect 8975 9400 9055 9450
rect 8975 9340 8985 9400
rect 9045 9340 9055 9400
rect 8975 9335 9055 9340
rect 9375 9510 9455 9515
rect 9375 9450 9385 9510
rect 9445 9450 9455 9510
rect 9375 9400 9455 9450
rect 9375 9340 9385 9400
rect 9445 9340 9455 9400
rect 9375 9335 9455 9340
rect 9775 9510 9855 9515
rect 9775 9450 9785 9510
rect 9845 9450 9855 9510
rect 9775 9400 9855 9450
rect 9775 9340 9785 9400
rect 9845 9340 9855 9400
rect 9775 9335 9855 9340
rect 10175 9510 10255 9515
rect 10175 9450 10185 9510
rect 10245 9450 10255 9510
rect 10175 9400 10255 9450
rect 10175 9340 10185 9400
rect 10245 9340 10255 9400
rect 10175 9335 10255 9340
rect 10575 9510 10655 9515
rect 10575 9450 10585 9510
rect 10645 9450 10655 9510
rect 10575 9400 10655 9450
rect 10575 9340 10585 9400
rect 10645 9340 10655 9400
rect 10575 9335 10655 9340
rect 10975 9510 11055 9515
rect 10975 9450 10985 9510
rect 11045 9450 11055 9510
rect 10975 9400 11055 9450
rect 10975 9340 10985 9400
rect 11045 9340 11055 9400
rect 10975 9335 11055 9340
rect 11375 9510 11455 9515
rect 11375 9450 11385 9510
rect 11445 9450 11455 9510
rect 11375 9400 11455 9450
rect 11375 9340 11385 9400
rect 11445 9340 11455 9400
rect 11375 9335 11455 9340
rect 11775 9510 11855 9515
rect 11775 9450 11785 9510
rect 11845 9450 11855 9510
rect 11775 9400 11855 9450
rect 11775 9340 11785 9400
rect 11845 9340 11855 9400
rect 11775 9335 11855 9340
rect 12175 9510 12255 9515
rect 12175 9450 12185 9510
rect 12245 9450 12255 9510
rect 12175 9400 12255 9450
rect 12175 9340 12185 9400
rect 12245 9340 12255 9400
rect 12175 9335 12255 9340
rect 12575 9510 12655 9515
rect 12575 9450 12585 9510
rect 12645 9450 12655 9510
rect 12575 9400 12655 9450
rect 12575 9340 12585 9400
rect 12645 9340 12655 9400
rect 12575 9335 12655 9340
rect 12975 9510 13055 9515
rect 12975 9450 12985 9510
rect 13045 9450 13055 9510
rect 12975 9400 13055 9450
rect 12975 9340 12985 9400
rect 13045 9340 13055 9400
rect 12975 9335 13055 9340
rect -215 9145 -155 9335
rect 185 9145 245 9335
rect 585 9145 645 9335
rect 985 9145 1045 9335
rect 1385 9145 1445 9335
rect 1785 9145 1845 9335
rect 2185 9145 2245 9335
rect 2585 9145 2645 9335
rect 2985 9145 3045 9335
rect 3385 9145 3445 9335
rect 3785 9145 3845 9335
rect 4185 9145 4245 9335
rect 4585 9145 4645 9335
rect 4985 9145 5045 9335
rect 5385 9145 5445 9335
rect 5785 9145 5845 9335
rect 6185 9145 6245 9335
rect 6585 9145 6645 9335
rect 6985 9145 7045 9335
rect 7385 9145 7445 9335
rect 7785 9145 7845 9335
rect 8185 9145 8245 9335
rect 8585 9145 8645 9335
rect 8985 9145 9045 9335
rect 9385 9145 9445 9335
rect 9785 9145 9845 9335
rect 10185 9145 10245 9335
rect 10585 9145 10645 9335
rect 10985 9145 11045 9335
rect 11385 9145 11445 9335
rect 11785 9145 11845 9335
rect 12185 9145 12245 9335
rect 12585 9145 12645 9335
rect 12985 9145 13045 9335
rect -225 9140 -145 9145
rect -225 9080 -215 9140
rect -155 9080 -145 9140
rect -225 9030 -145 9080
rect -225 8970 -215 9030
rect -155 8970 -145 9030
rect -225 8965 -145 8970
rect 175 9140 255 9145
rect 175 9080 185 9140
rect 245 9080 255 9140
rect 175 9030 255 9080
rect 175 8970 185 9030
rect 245 8970 255 9030
rect 175 8965 255 8970
rect 575 9140 655 9145
rect 575 9080 585 9140
rect 645 9080 655 9140
rect 575 9030 655 9080
rect 575 8970 585 9030
rect 645 8970 655 9030
rect 575 8965 655 8970
rect 975 9140 1055 9145
rect 975 9080 985 9140
rect 1045 9080 1055 9140
rect 975 9030 1055 9080
rect 975 8970 985 9030
rect 1045 8970 1055 9030
rect 975 8965 1055 8970
rect 1375 9140 1455 9145
rect 1375 9080 1385 9140
rect 1445 9080 1455 9140
rect 1375 9030 1455 9080
rect 1375 8970 1385 9030
rect 1445 8970 1455 9030
rect 1375 8965 1455 8970
rect 1775 9140 1855 9145
rect 1775 9080 1785 9140
rect 1845 9080 1855 9140
rect 1775 9030 1855 9080
rect 1775 8970 1785 9030
rect 1845 8970 1855 9030
rect 1775 8965 1855 8970
rect 2175 9140 2255 9145
rect 2175 9080 2185 9140
rect 2245 9080 2255 9140
rect 2175 9030 2255 9080
rect 2175 8970 2185 9030
rect 2245 8970 2255 9030
rect 2175 8965 2255 8970
rect 2575 9140 2655 9145
rect 2575 9080 2585 9140
rect 2645 9080 2655 9140
rect 2575 9030 2655 9080
rect 2575 8970 2585 9030
rect 2645 8970 2655 9030
rect 2575 8965 2655 8970
rect 2975 9140 3055 9145
rect 2975 9080 2985 9140
rect 3045 9080 3055 9140
rect 2975 9030 3055 9080
rect 2975 8970 2985 9030
rect 3045 8970 3055 9030
rect 2975 8965 3055 8970
rect 3375 9140 3455 9145
rect 3375 9080 3385 9140
rect 3445 9080 3455 9140
rect 3375 9030 3455 9080
rect 3375 8970 3385 9030
rect 3445 8970 3455 9030
rect 3375 8965 3455 8970
rect 3775 9140 3855 9145
rect 3775 9080 3785 9140
rect 3845 9080 3855 9140
rect 3775 9030 3855 9080
rect 3775 8970 3785 9030
rect 3845 8970 3855 9030
rect 3775 8965 3855 8970
rect 4175 9140 4255 9145
rect 4175 9080 4185 9140
rect 4245 9080 4255 9140
rect 4175 9030 4255 9080
rect 4175 8970 4185 9030
rect 4245 8970 4255 9030
rect 4175 8965 4255 8970
rect 4575 9140 4655 9145
rect 4575 9080 4585 9140
rect 4645 9080 4655 9140
rect 4575 9030 4655 9080
rect 4575 8970 4585 9030
rect 4645 8970 4655 9030
rect 4575 8965 4655 8970
rect 4975 9140 5055 9145
rect 4975 9080 4985 9140
rect 5045 9080 5055 9140
rect 4975 9030 5055 9080
rect 4975 8970 4985 9030
rect 5045 8970 5055 9030
rect 4975 8965 5055 8970
rect 5375 9140 5455 9145
rect 5375 9080 5385 9140
rect 5445 9080 5455 9140
rect 5375 9030 5455 9080
rect 5375 8970 5385 9030
rect 5445 8970 5455 9030
rect 5375 8965 5455 8970
rect 5775 9140 5855 9145
rect 5775 9080 5785 9140
rect 5845 9080 5855 9140
rect 5775 9030 5855 9080
rect 5775 8970 5785 9030
rect 5845 8970 5855 9030
rect 5775 8965 5855 8970
rect 6175 9140 6255 9145
rect 6175 9080 6185 9140
rect 6245 9080 6255 9140
rect 6175 9030 6255 9080
rect 6175 8970 6185 9030
rect 6245 8970 6255 9030
rect 6175 8965 6255 8970
rect 6575 9140 6655 9145
rect 6575 9080 6585 9140
rect 6645 9080 6655 9140
rect 6575 9030 6655 9080
rect 6575 8970 6585 9030
rect 6645 8970 6655 9030
rect 6575 8965 6655 8970
rect 6975 9140 7055 9145
rect 6975 9080 6985 9140
rect 7045 9080 7055 9140
rect 6975 9030 7055 9080
rect 6975 8970 6985 9030
rect 7045 8970 7055 9030
rect 6975 8965 7055 8970
rect 7375 9140 7455 9145
rect 7375 9080 7385 9140
rect 7445 9080 7455 9140
rect 7375 9030 7455 9080
rect 7375 8970 7385 9030
rect 7445 8970 7455 9030
rect 7375 8965 7455 8970
rect 7775 9140 7855 9145
rect 7775 9080 7785 9140
rect 7845 9080 7855 9140
rect 7775 9030 7855 9080
rect 7775 8970 7785 9030
rect 7845 8970 7855 9030
rect 7775 8965 7855 8970
rect 8175 9140 8255 9145
rect 8175 9080 8185 9140
rect 8245 9080 8255 9140
rect 8175 9030 8255 9080
rect 8175 8970 8185 9030
rect 8245 8970 8255 9030
rect 8175 8965 8255 8970
rect 8575 9140 8655 9145
rect 8575 9080 8585 9140
rect 8645 9080 8655 9140
rect 8575 9030 8655 9080
rect 8575 8970 8585 9030
rect 8645 8970 8655 9030
rect 8575 8965 8655 8970
rect 8975 9140 9055 9145
rect 8975 9080 8985 9140
rect 9045 9080 9055 9140
rect 8975 9030 9055 9080
rect 8975 8970 8985 9030
rect 9045 8970 9055 9030
rect 8975 8965 9055 8970
rect 9375 9140 9455 9145
rect 9375 9080 9385 9140
rect 9445 9080 9455 9140
rect 9375 9030 9455 9080
rect 9375 8970 9385 9030
rect 9445 8970 9455 9030
rect 9375 8965 9455 8970
rect 9775 9140 9855 9145
rect 9775 9080 9785 9140
rect 9845 9080 9855 9140
rect 9775 9030 9855 9080
rect 9775 8970 9785 9030
rect 9845 8970 9855 9030
rect 9775 8965 9855 8970
rect 10175 9140 10255 9145
rect 10175 9080 10185 9140
rect 10245 9080 10255 9140
rect 10175 9030 10255 9080
rect 10175 8970 10185 9030
rect 10245 8970 10255 9030
rect 10175 8965 10255 8970
rect 10575 9140 10655 9145
rect 10575 9080 10585 9140
rect 10645 9080 10655 9140
rect 10575 9030 10655 9080
rect 10575 8970 10585 9030
rect 10645 8970 10655 9030
rect 10575 8965 10655 8970
rect 10975 9140 11055 9145
rect 10975 9080 10985 9140
rect 11045 9080 11055 9140
rect 10975 9030 11055 9080
rect 10975 8970 10985 9030
rect 11045 8970 11055 9030
rect 10975 8965 11055 8970
rect 11375 9140 11455 9145
rect 11375 9080 11385 9140
rect 11445 9080 11455 9140
rect 11375 9030 11455 9080
rect 11375 8970 11385 9030
rect 11445 8970 11455 9030
rect 11375 8965 11455 8970
rect 11775 9140 11855 9145
rect 11775 9080 11785 9140
rect 11845 9080 11855 9140
rect 11775 9030 11855 9080
rect 11775 8970 11785 9030
rect 11845 8970 11855 9030
rect 11775 8965 11855 8970
rect 12175 9140 12255 9145
rect 12175 9080 12185 9140
rect 12245 9080 12255 9140
rect 12175 9030 12255 9080
rect 12175 8970 12185 9030
rect 12245 8970 12255 9030
rect 12175 8965 12255 8970
rect 12575 9140 12655 9145
rect 12575 9080 12585 9140
rect 12645 9080 12655 9140
rect 12575 9030 12655 9080
rect 12575 8970 12585 9030
rect 12645 8970 12655 9030
rect 12575 8965 12655 8970
rect 12975 9140 13055 9145
rect 12975 9080 12985 9140
rect 13045 9080 13055 9140
rect 12975 9030 13055 9080
rect 12975 8970 12985 9030
rect 13045 8970 13055 9030
rect 12975 8965 13055 8970
rect -215 8775 -155 8965
rect 185 8775 245 8965
rect 585 8775 645 8965
rect 985 8775 1045 8965
rect 1385 8775 1445 8965
rect 1785 8775 1845 8965
rect 2185 8775 2245 8965
rect 2585 8775 2645 8965
rect 2985 8775 3045 8965
rect 3385 8775 3445 8965
rect 3785 8775 3845 8965
rect 4185 8775 4245 8965
rect 4585 8775 4645 8965
rect 4985 8775 5045 8965
rect 5385 8775 5445 8965
rect 5785 8775 5845 8965
rect 6185 8775 6245 8965
rect 6585 8775 6645 8965
rect 6985 8775 7045 8965
rect 7385 8775 7445 8965
rect 7785 8775 7845 8965
rect 8185 8775 8245 8965
rect 8585 8775 8645 8965
rect 8985 8775 9045 8965
rect 9385 8775 9445 8965
rect 9785 8775 9845 8965
rect 10185 8775 10245 8965
rect 10585 8775 10645 8965
rect 10985 8775 11045 8965
rect 11385 8775 11445 8965
rect 11785 8775 11845 8965
rect 12185 8775 12245 8965
rect 12585 8775 12645 8965
rect 12985 8775 13045 8965
rect -225 8770 -145 8775
rect -225 8710 -215 8770
rect -155 8710 -145 8770
rect -225 8660 -145 8710
rect -225 8600 -215 8660
rect -155 8600 -145 8660
rect -225 8595 -145 8600
rect 175 8770 255 8775
rect 175 8710 185 8770
rect 245 8710 255 8770
rect 175 8660 255 8710
rect 175 8600 185 8660
rect 245 8600 255 8660
rect 175 8595 255 8600
rect 575 8770 655 8775
rect 575 8710 585 8770
rect 645 8710 655 8770
rect 575 8660 655 8710
rect 575 8600 585 8660
rect 645 8600 655 8660
rect 575 8595 655 8600
rect 975 8770 1055 8775
rect 975 8710 985 8770
rect 1045 8710 1055 8770
rect 975 8660 1055 8710
rect 975 8600 985 8660
rect 1045 8600 1055 8660
rect 975 8595 1055 8600
rect 1375 8770 1455 8775
rect 1375 8710 1385 8770
rect 1445 8710 1455 8770
rect 1375 8660 1455 8710
rect 1375 8600 1385 8660
rect 1445 8600 1455 8660
rect 1375 8595 1455 8600
rect 1775 8770 1855 8775
rect 1775 8710 1785 8770
rect 1845 8710 1855 8770
rect 1775 8660 1855 8710
rect 1775 8600 1785 8660
rect 1845 8600 1855 8660
rect 1775 8595 1855 8600
rect 2175 8770 2255 8775
rect 2175 8710 2185 8770
rect 2245 8710 2255 8770
rect 2175 8660 2255 8710
rect 2175 8600 2185 8660
rect 2245 8600 2255 8660
rect 2175 8595 2255 8600
rect 2575 8770 2655 8775
rect 2575 8710 2585 8770
rect 2645 8710 2655 8770
rect 2575 8660 2655 8710
rect 2575 8600 2585 8660
rect 2645 8600 2655 8660
rect 2575 8595 2655 8600
rect 2975 8770 3055 8775
rect 2975 8710 2985 8770
rect 3045 8710 3055 8770
rect 2975 8660 3055 8710
rect 2975 8600 2985 8660
rect 3045 8600 3055 8660
rect 2975 8595 3055 8600
rect 3375 8770 3455 8775
rect 3375 8710 3385 8770
rect 3445 8710 3455 8770
rect 3375 8660 3455 8710
rect 3375 8600 3385 8660
rect 3445 8600 3455 8660
rect 3375 8595 3455 8600
rect 3775 8770 3855 8775
rect 3775 8710 3785 8770
rect 3845 8710 3855 8770
rect 3775 8660 3855 8710
rect 3775 8600 3785 8660
rect 3845 8600 3855 8660
rect 3775 8595 3855 8600
rect 4175 8770 4255 8775
rect 4175 8710 4185 8770
rect 4245 8710 4255 8770
rect 4175 8660 4255 8710
rect 4175 8600 4185 8660
rect 4245 8600 4255 8660
rect 4175 8595 4255 8600
rect 4575 8770 4655 8775
rect 4575 8710 4585 8770
rect 4645 8710 4655 8770
rect 4575 8660 4655 8710
rect 4575 8600 4585 8660
rect 4645 8600 4655 8660
rect 4575 8595 4655 8600
rect 4975 8770 5055 8775
rect 4975 8710 4985 8770
rect 5045 8710 5055 8770
rect 4975 8660 5055 8710
rect 4975 8600 4985 8660
rect 5045 8600 5055 8660
rect 4975 8595 5055 8600
rect 5375 8770 5455 8775
rect 5375 8710 5385 8770
rect 5445 8710 5455 8770
rect 5375 8660 5455 8710
rect 5375 8600 5385 8660
rect 5445 8600 5455 8660
rect 5375 8595 5455 8600
rect 5775 8770 5855 8775
rect 5775 8710 5785 8770
rect 5845 8710 5855 8770
rect 5775 8660 5855 8710
rect 5775 8600 5785 8660
rect 5845 8600 5855 8660
rect 5775 8595 5855 8600
rect 6175 8770 6255 8775
rect 6175 8710 6185 8770
rect 6245 8710 6255 8770
rect 6175 8660 6255 8710
rect 6175 8600 6185 8660
rect 6245 8600 6255 8660
rect 6175 8595 6255 8600
rect 6575 8770 6655 8775
rect 6575 8710 6585 8770
rect 6645 8710 6655 8770
rect 6575 8660 6655 8710
rect 6575 8600 6585 8660
rect 6645 8600 6655 8660
rect 6575 8595 6655 8600
rect 6975 8770 7055 8775
rect 6975 8710 6985 8770
rect 7045 8710 7055 8770
rect 6975 8660 7055 8710
rect 6975 8600 6985 8660
rect 7045 8600 7055 8660
rect 6975 8595 7055 8600
rect 7375 8770 7455 8775
rect 7375 8710 7385 8770
rect 7445 8710 7455 8770
rect 7375 8660 7455 8710
rect 7375 8600 7385 8660
rect 7445 8600 7455 8660
rect 7375 8595 7455 8600
rect 7775 8770 7855 8775
rect 7775 8710 7785 8770
rect 7845 8710 7855 8770
rect 7775 8660 7855 8710
rect 7775 8600 7785 8660
rect 7845 8600 7855 8660
rect 7775 8595 7855 8600
rect 8175 8770 8255 8775
rect 8175 8710 8185 8770
rect 8245 8710 8255 8770
rect 8175 8660 8255 8710
rect 8175 8600 8185 8660
rect 8245 8600 8255 8660
rect 8175 8595 8255 8600
rect 8575 8770 8655 8775
rect 8575 8710 8585 8770
rect 8645 8710 8655 8770
rect 8575 8660 8655 8710
rect 8575 8600 8585 8660
rect 8645 8600 8655 8660
rect 8575 8595 8655 8600
rect 8975 8770 9055 8775
rect 8975 8710 8985 8770
rect 9045 8710 9055 8770
rect 8975 8660 9055 8710
rect 8975 8600 8985 8660
rect 9045 8600 9055 8660
rect 8975 8595 9055 8600
rect 9375 8770 9455 8775
rect 9375 8710 9385 8770
rect 9445 8710 9455 8770
rect 9375 8660 9455 8710
rect 9375 8600 9385 8660
rect 9445 8600 9455 8660
rect 9375 8595 9455 8600
rect 9775 8770 9855 8775
rect 9775 8710 9785 8770
rect 9845 8710 9855 8770
rect 9775 8660 9855 8710
rect 9775 8600 9785 8660
rect 9845 8600 9855 8660
rect 9775 8595 9855 8600
rect 10175 8770 10255 8775
rect 10175 8710 10185 8770
rect 10245 8710 10255 8770
rect 10175 8660 10255 8710
rect 10175 8600 10185 8660
rect 10245 8600 10255 8660
rect 10175 8595 10255 8600
rect 10575 8770 10655 8775
rect 10575 8710 10585 8770
rect 10645 8710 10655 8770
rect 10575 8660 10655 8710
rect 10575 8600 10585 8660
rect 10645 8600 10655 8660
rect 10575 8595 10655 8600
rect 10975 8770 11055 8775
rect 10975 8710 10985 8770
rect 11045 8710 11055 8770
rect 10975 8660 11055 8710
rect 10975 8600 10985 8660
rect 11045 8600 11055 8660
rect 10975 8595 11055 8600
rect 11375 8770 11455 8775
rect 11375 8710 11385 8770
rect 11445 8710 11455 8770
rect 11375 8660 11455 8710
rect 11375 8600 11385 8660
rect 11445 8600 11455 8660
rect 11375 8595 11455 8600
rect 11775 8770 11855 8775
rect 11775 8710 11785 8770
rect 11845 8710 11855 8770
rect 11775 8660 11855 8710
rect 11775 8600 11785 8660
rect 11845 8600 11855 8660
rect 11775 8595 11855 8600
rect 12175 8770 12255 8775
rect 12175 8710 12185 8770
rect 12245 8710 12255 8770
rect 12175 8660 12255 8710
rect 12175 8600 12185 8660
rect 12245 8600 12255 8660
rect 12175 8595 12255 8600
rect 12575 8770 12655 8775
rect 12575 8710 12585 8770
rect 12645 8710 12655 8770
rect 12575 8660 12655 8710
rect 12575 8600 12585 8660
rect 12645 8600 12655 8660
rect 12575 8595 12655 8600
rect 12975 8770 13055 8775
rect 12975 8710 12985 8770
rect 13045 8710 13055 8770
rect 12975 8660 13055 8710
rect 12975 8600 12985 8660
rect 13045 8600 13055 8660
rect 12975 8595 13055 8600
rect -215 8405 -155 8595
rect 185 8405 245 8595
rect 585 8405 645 8595
rect 985 8405 1045 8595
rect 1385 8405 1445 8595
rect 1785 8405 1845 8595
rect 2185 8405 2245 8595
rect 2585 8405 2645 8595
rect 2985 8405 3045 8595
rect 3385 8405 3445 8595
rect 3785 8405 3845 8595
rect 4185 8405 4245 8595
rect 4585 8405 4645 8595
rect 4985 8405 5045 8595
rect 5385 8405 5445 8595
rect 5785 8405 5845 8595
rect 6185 8405 6245 8595
rect 6585 8405 6645 8595
rect 6985 8405 7045 8595
rect 7385 8405 7445 8595
rect 7785 8405 7845 8595
rect 8185 8405 8245 8595
rect 8585 8405 8645 8595
rect 8985 8405 9045 8595
rect 9385 8405 9445 8595
rect 9785 8405 9845 8595
rect 10185 8405 10245 8595
rect 10585 8405 10645 8595
rect 10985 8405 11045 8595
rect 11385 8405 11445 8595
rect 11785 8405 11845 8595
rect 12185 8405 12245 8595
rect 12585 8405 12645 8595
rect 12985 8405 13045 8595
rect -225 8400 -145 8405
rect -225 8340 -215 8400
rect -155 8340 -145 8400
rect -225 8290 -145 8340
rect -225 8230 -215 8290
rect -155 8230 -145 8290
rect -225 8225 -145 8230
rect 175 8400 255 8405
rect 175 8340 185 8400
rect 245 8340 255 8400
rect 175 8290 255 8340
rect 175 8230 185 8290
rect 245 8230 255 8290
rect 175 8225 255 8230
rect 575 8400 655 8405
rect 575 8340 585 8400
rect 645 8340 655 8400
rect 575 8290 655 8340
rect 575 8230 585 8290
rect 645 8230 655 8290
rect 575 8225 655 8230
rect 975 8400 1055 8405
rect 975 8340 985 8400
rect 1045 8340 1055 8400
rect 975 8290 1055 8340
rect 975 8230 985 8290
rect 1045 8230 1055 8290
rect 975 8225 1055 8230
rect 1375 8400 1455 8405
rect 1375 8340 1385 8400
rect 1445 8340 1455 8400
rect 1375 8290 1455 8340
rect 1375 8230 1385 8290
rect 1445 8230 1455 8290
rect 1375 8225 1455 8230
rect 1775 8400 1855 8405
rect 1775 8340 1785 8400
rect 1845 8340 1855 8400
rect 1775 8290 1855 8340
rect 1775 8230 1785 8290
rect 1845 8230 1855 8290
rect 1775 8225 1855 8230
rect 2175 8400 2255 8405
rect 2175 8340 2185 8400
rect 2245 8340 2255 8400
rect 2175 8290 2255 8340
rect 2175 8230 2185 8290
rect 2245 8230 2255 8290
rect 2175 8225 2255 8230
rect 2575 8400 2655 8405
rect 2575 8340 2585 8400
rect 2645 8340 2655 8400
rect 2575 8290 2655 8340
rect 2575 8230 2585 8290
rect 2645 8230 2655 8290
rect 2575 8225 2655 8230
rect 2975 8400 3055 8405
rect 2975 8340 2985 8400
rect 3045 8340 3055 8400
rect 2975 8290 3055 8340
rect 2975 8230 2985 8290
rect 3045 8230 3055 8290
rect 2975 8225 3055 8230
rect 3375 8400 3455 8405
rect 3375 8340 3385 8400
rect 3445 8340 3455 8400
rect 3375 8290 3455 8340
rect 3375 8230 3385 8290
rect 3445 8230 3455 8290
rect 3375 8225 3455 8230
rect 3775 8400 3855 8405
rect 3775 8340 3785 8400
rect 3845 8340 3855 8400
rect 3775 8290 3855 8340
rect 3775 8230 3785 8290
rect 3845 8230 3855 8290
rect 3775 8225 3855 8230
rect 4175 8400 4255 8405
rect 4175 8340 4185 8400
rect 4245 8340 4255 8400
rect 4175 8290 4255 8340
rect 4175 8230 4185 8290
rect 4245 8230 4255 8290
rect 4175 8225 4255 8230
rect 4575 8400 4655 8405
rect 4575 8340 4585 8400
rect 4645 8340 4655 8400
rect 4575 8290 4655 8340
rect 4575 8230 4585 8290
rect 4645 8230 4655 8290
rect 4575 8225 4655 8230
rect 4975 8400 5055 8405
rect 4975 8340 4985 8400
rect 5045 8340 5055 8400
rect 4975 8290 5055 8340
rect 4975 8230 4985 8290
rect 5045 8230 5055 8290
rect 4975 8225 5055 8230
rect 5375 8400 5455 8405
rect 5375 8340 5385 8400
rect 5445 8340 5455 8400
rect 5375 8290 5455 8340
rect 5375 8230 5385 8290
rect 5445 8230 5455 8290
rect 5375 8225 5455 8230
rect 5775 8400 5855 8405
rect 5775 8340 5785 8400
rect 5845 8340 5855 8400
rect 5775 8290 5855 8340
rect 5775 8230 5785 8290
rect 5845 8230 5855 8290
rect 5775 8225 5855 8230
rect 6175 8400 6255 8405
rect 6175 8340 6185 8400
rect 6245 8340 6255 8400
rect 6175 8290 6255 8340
rect 6175 8230 6185 8290
rect 6245 8230 6255 8290
rect 6175 8225 6255 8230
rect 6575 8400 6655 8405
rect 6575 8340 6585 8400
rect 6645 8340 6655 8400
rect 6575 8290 6655 8340
rect 6575 8230 6585 8290
rect 6645 8230 6655 8290
rect 6575 8225 6655 8230
rect 6975 8400 7055 8405
rect 6975 8340 6985 8400
rect 7045 8340 7055 8400
rect 6975 8290 7055 8340
rect 6975 8230 6985 8290
rect 7045 8230 7055 8290
rect 6975 8225 7055 8230
rect 7375 8400 7455 8405
rect 7375 8340 7385 8400
rect 7445 8340 7455 8400
rect 7375 8290 7455 8340
rect 7375 8230 7385 8290
rect 7445 8230 7455 8290
rect 7375 8225 7455 8230
rect 7775 8400 7855 8405
rect 7775 8340 7785 8400
rect 7845 8340 7855 8400
rect 7775 8290 7855 8340
rect 7775 8230 7785 8290
rect 7845 8230 7855 8290
rect 7775 8225 7855 8230
rect 8175 8400 8255 8405
rect 8175 8340 8185 8400
rect 8245 8340 8255 8400
rect 8175 8290 8255 8340
rect 8175 8230 8185 8290
rect 8245 8230 8255 8290
rect 8175 8225 8255 8230
rect 8575 8400 8655 8405
rect 8575 8340 8585 8400
rect 8645 8340 8655 8400
rect 8575 8290 8655 8340
rect 8575 8230 8585 8290
rect 8645 8230 8655 8290
rect 8575 8225 8655 8230
rect 8975 8400 9055 8405
rect 8975 8340 8985 8400
rect 9045 8340 9055 8400
rect 8975 8290 9055 8340
rect 8975 8230 8985 8290
rect 9045 8230 9055 8290
rect 8975 8225 9055 8230
rect 9375 8400 9455 8405
rect 9375 8340 9385 8400
rect 9445 8340 9455 8400
rect 9375 8290 9455 8340
rect 9375 8230 9385 8290
rect 9445 8230 9455 8290
rect 9375 8225 9455 8230
rect 9775 8400 9855 8405
rect 9775 8340 9785 8400
rect 9845 8340 9855 8400
rect 9775 8290 9855 8340
rect 9775 8230 9785 8290
rect 9845 8230 9855 8290
rect 9775 8225 9855 8230
rect 10175 8400 10255 8405
rect 10175 8340 10185 8400
rect 10245 8340 10255 8400
rect 10175 8290 10255 8340
rect 10175 8230 10185 8290
rect 10245 8230 10255 8290
rect 10175 8225 10255 8230
rect 10575 8400 10655 8405
rect 10575 8340 10585 8400
rect 10645 8340 10655 8400
rect 10575 8290 10655 8340
rect 10575 8230 10585 8290
rect 10645 8230 10655 8290
rect 10575 8225 10655 8230
rect 10975 8400 11055 8405
rect 10975 8340 10985 8400
rect 11045 8340 11055 8400
rect 10975 8290 11055 8340
rect 10975 8230 10985 8290
rect 11045 8230 11055 8290
rect 10975 8225 11055 8230
rect 11375 8400 11455 8405
rect 11375 8340 11385 8400
rect 11445 8340 11455 8400
rect 11375 8290 11455 8340
rect 11375 8230 11385 8290
rect 11445 8230 11455 8290
rect 11375 8225 11455 8230
rect 11775 8400 11855 8405
rect 11775 8340 11785 8400
rect 11845 8340 11855 8400
rect 11775 8290 11855 8340
rect 11775 8230 11785 8290
rect 11845 8230 11855 8290
rect 11775 8225 11855 8230
rect 12175 8400 12255 8405
rect 12175 8340 12185 8400
rect 12245 8340 12255 8400
rect 12175 8290 12255 8340
rect 12175 8230 12185 8290
rect 12245 8230 12255 8290
rect 12175 8225 12255 8230
rect 12575 8400 12655 8405
rect 12575 8340 12585 8400
rect 12645 8340 12655 8400
rect 12575 8290 12655 8340
rect 12575 8230 12585 8290
rect 12645 8230 12655 8290
rect 12575 8225 12655 8230
rect 12975 8400 13055 8405
rect 12975 8340 12985 8400
rect 13045 8340 13055 8400
rect 12975 8290 13055 8340
rect 12975 8230 12985 8290
rect 13045 8230 13055 8290
rect 12975 8225 13055 8230
rect -215 8035 -155 8225
rect 185 8035 245 8225
rect 585 8035 645 8225
rect 985 8035 1045 8225
rect 1385 8035 1445 8225
rect 1785 8035 1845 8225
rect 2185 8035 2245 8225
rect 2585 8035 2645 8225
rect 2985 8035 3045 8225
rect 3385 8035 3445 8225
rect 3785 8035 3845 8225
rect 4185 8035 4245 8225
rect 4585 8035 4645 8225
rect 4985 8035 5045 8225
rect 5385 8035 5445 8225
rect 5785 8035 5845 8225
rect 6185 8035 6245 8225
rect 6585 8035 6645 8225
rect 6985 8035 7045 8225
rect 7385 8035 7445 8225
rect 7785 8035 7845 8225
rect 8185 8035 8245 8225
rect 8585 8035 8645 8225
rect 8985 8035 9045 8225
rect 9385 8035 9445 8225
rect 9785 8035 9845 8225
rect 10185 8035 10245 8225
rect 10585 8035 10645 8225
rect 10985 8035 11045 8225
rect 11385 8035 11445 8225
rect 11785 8035 11845 8225
rect 12185 8035 12245 8225
rect 12585 8035 12645 8225
rect 12985 8035 13045 8225
rect -225 8030 -145 8035
rect -225 7970 -215 8030
rect -155 7970 -145 8030
rect -225 7920 -145 7970
rect -225 7860 -215 7920
rect -155 7860 -145 7920
rect -225 7855 -145 7860
rect 175 8030 255 8035
rect 175 7970 185 8030
rect 245 7970 255 8030
rect 175 7920 255 7970
rect 175 7860 185 7920
rect 245 7860 255 7920
rect 175 7855 255 7860
rect 575 8030 655 8035
rect 575 7970 585 8030
rect 645 7970 655 8030
rect 575 7920 655 7970
rect 575 7860 585 7920
rect 645 7860 655 7920
rect 575 7855 655 7860
rect 975 8030 1055 8035
rect 975 7970 985 8030
rect 1045 7970 1055 8030
rect 975 7920 1055 7970
rect 975 7860 985 7920
rect 1045 7860 1055 7920
rect 975 7855 1055 7860
rect 1375 8030 1455 8035
rect 1375 7970 1385 8030
rect 1445 7970 1455 8030
rect 1375 7920 1455 7970
rect 1375 7860 1385 7920
rect 1445 7860 1455 7920
rect 1375 7855 1455 7860
rect 1775 8030 1855 8035
rect 1775 7970 1785 8030
rect 1845 7970 1855 8030
rect 1775 7920 1855 7970
rect 1775 7860 1785 7920
rect 1845 7860 1855 7920
rect 1775 7855 1855 7860
rect 2175 8030 2255 8035
rect 2175 7970 2185 8030
rect 2245 7970 2255 8030
rect 2175 7920 2255 7970
rect 2175 7860 2185 7920
rect 2245 7860 2255 7920
rect 2175 7855 2255 7860
rect 2575 8030 2655 8035
rect 2575 7970 2585 8030
rect 2645 7970 2655 8030
rect 2575 7920 2655 7970
rect 2575 7860 2585 7920
rect 2645 7860 2655 7920
rect 2575 7855 2655 7860
rect 2975 8030 3055 8035
rect 2975 7970 2985 8030
rect 3045 7970 3055 8030
rect 2975 7920 3055 7970
rect 2975 7860 2985 7920
rect 3045 7860 3055 7920
rect 2975 7855 3055 7860
rect 3375 8030 3455 8035
rect 3375 7970 3385 8030
rect 3445 7970 3455 8030
rect 3375 7920 3455 7970
rect 3375 7860 3385 7920
rect 3445 7860 3455 7920
rect 3375 7855 3455 7860
rect 3775 8030 3855 8035
rect 3775 7970 3785 8030
rect 3845 7970 3855 8030
rect 3775 7920 3855 7970
rect 3775 7860 3785 7920
rect 3845 7860 3855 7920
rect 3775 7855 3855 7860
rect 4175 8030 4255 8035
rect 4175 7970 4185 8030
rect 4245 7970 4255 8030
rect 4175 7920 4255 7970
rect 4175 7860 4185 7920
rect 4245 7860 4255 7920
rect 4175 7855 4255 7860
rect 4575 8030 4655 8035
rect 4575 7970 4585 8030
rect 4645 7970 4655 8030
rect 4575 7920 4655 7970
rect 4575 7860 4585 7920
rect 4645 7860 4655 7920
rect 4575 7855 4655 7860
rect 4975 8030 5055 8035
rect 4975 7970 4985 8030
rect 5045 7970 5055 8030
rect 4975 7920 5055 7970
rect 4975 7860 4985 7920
rect 5045 7860 5055 7920
rect 4975 7855 5055 7860
rect 5375 8030 5455 8035
rect 5375 7970 5385 8030
rect 5445 7970 5455 8030
rect 5375 7920 5455 7970
rect 5375 7860 5385 7920
rect 5445 7860 5455 7920
rect 5375 7855 5455 7860
rect 5775 8030 5855 8035
rect 5775 7970 5785 8030
rect 5845 7970 5855 8030
rect 5775 7920 5855 7970
rect 5775 7860 5785 7920
rect 5845 7860 5855 7920
rect 5775 7855 5855 7860
rect 6175 8030 6255 8035
rect 6175 7970 6185 8030
rect 6245 7970 6255 8030
rect 6175 7920 6255 7970
rect 6175 7860 6185 7920
rect 6245 7860 6255 7920
rect 6175 7855 6255 7860
rect 6575 8030 6655 8035
rect 6575 7970 6585 8030
rect 6645 7970 6655 8030
rect 6575 7920 6655 7970
rect 6575 7860 6585 7920
rect 6645 7860 6655 7920
rect 6575 7855 6655 7860
rect 6975 8030 7055 8035
rect 6975 7970 6985 8030
rect 7045 7970 7055 8030
rect 6975 7920 7055 7970
rect 6975 7860 6985 7920
rect 7045 7860 7055 7920
rect 6975 7855 7055 7860
rect 7375 8030 7455 8035
rect 7375 7970 7385 8030
rect 7445 7970 7455 8030
rect 7375 7920 7455 7970
rect 7375 7860 7385 7920
rect 7445 7860 7455 7920
rect 7375 7855 7455 7860
rect 7775 8030 7855 8035
rect 7775 7970 7785 8030
rect 7845 7970 7855 8030
rect 7775 7920 7855 7970
rect 7775 7860 7785 7920
rect 7845 7860 7855 7920
rect 7775 7855 7855 7860
rect 8175 8030 8255 8035
rect 8175 7970 8185 8030
rect 8245 7970 8255 8030
rect 8175 7920 8255 7970
rect 8175 7860 8185 7920
rect 8245 7860 8255 7920
rect 8175 7855 8255 7860
rect 8575 8030 8655 8035
rect 8575 7970 8585 8030
rect 8645 7970 8655 8030
rect 8575 7920 8655 7970
rect 8575 7860 8585 7920
rect 8645 7860 8655 7920
rect 8575 7855 8655 7860
rect 8975 8030 9055 8035
rect 8975 7970 8985 8030
rect 9045 7970 9055 8030
rect 8975 7920 9055 7970
rect 8975 7860 8985 7920
rect 9045 7860 9055 7920
rect 8975 7855 9055 7860
rect 9375 8030 9455 8035
rect 9375 7970 9385 8030
rect 9445 7970 9455 8030
rect 9375 7920 9455 7970
rect 9375 7860 9385 7920
rect 9445 7860 9455 7920
rect 9375 7855 9455 7860
rect 9775 8030 9855 8035
rect 9775 7970 9785 8030
rect 9845 7970 9855 8030
rect 9775 7920 9855 7970
rect 9775 7860 9785 7920
rect 9845 7860 9855 7920
rect 9775 7855 9855 7860
rect 10175 8030 10255 8035
rect 10175 7970 10185 8030
rect 10245 7970 10255 8030
rect 10175 7920 10255 7970
rect 10175 7860 10185 7920
rect 10245 7860 10255 7920
rect 10175 7855 10255 7860
rect 10575 8030 10655 8035
rect 10575 7970 10585 8030
rect 10645 7970 10655 8030
rect 10575 7920 10655 7970
rect 10575 7860 10585 7920
rect 10645 7860 10655 7920
rect 10575 7855 10655 7860
rect 10975 8030 11055 8035
rect 10975 7970 10985 8030
rect 11045 7970 11055 8030
rect 10975 7920 11055 7970
rect 10975 7860 10985 7920
rect 11045 7860 11055 7920
rect 10975 7855 11055 7860
rect 11375 8030 11455 8035
rect 11375 7970 11385 8030
rect 11445 7970 11455 8030
rect 11375 7920 11455 7970
rect 11375 7860 11385 7920
rect 11445 7860 11455 7920
rect 11375 7855 11455 7860
rect 11775 8030 11855 8035
rect 11775 7970 11785 8030
rect 11845 7970 11855 8030
rect 11775 7920 11855 7970
rect 11775 7860 11785 7920
rect 11845 7860 11855 7920
rect 11775 7855 11855 7860
rect 12175 8030 12255 8035
rect 12175 7970 12185 8030
rect 12245 7970 12255 8030
rect 12175 7920 12255 7970
rect 12175 7860 12185 7920
rect 12245 7860 12255 7920
rect 12175 7855 12255 7860
rect 12575 8030 12655 8035
rect 12575 7970 12585 8030
rect 12645 7970 12655 8030
rect 12575 7920 12655 7970
rect 12575 7860 12585 7920
rect 12645 7860 12655 7920
rect 12575 7855 12655 7860
rect 12975 8030 13055 8035
rect 12975 7970 12985 8030
rect 13045 7970 13055 8030
rect 12975 7920 13055 7970
rect 12975 7860 12985 7920
rect 13045 7860 13055 7920
rect 12975 7855 13055 7860
rect -215 7665 -155 7855
rect 185 7665 245 7855
rect 585 7665 645 7855
rect 985 7665 1045 7855
rect 1385 7665 1445 7855
rect 1785 7665 1845 7855
rect 2185 7665 2245 7855
rect 2585 7665 2645 7855
rect 2985 7665 3045 7855
rect 3385 7665 3445 7855
rect 3785 7665 3845 7855
rect 4185 7665 4245 7855
rect 4585 7665 4645 7855
rect 4985 7665 5045 7855
rect 5385 7665 5445 7855
rect 5785 7665 5845 7855
rect 6185 7665 6245 7855
rect 6585 7665 6645 7855
rect 6985 7665 7045 7855
rect 7385 7665 7445 7855
rect 7785 7665 7845 7855
rect 8185 7665 8245 7855
rect 8585 7665 8645 7855
rect 8985 7665 9045 7855
rect 9385 7665 9445 7855
rect 9785 7665 9845 7855
rect 10185 7665 10245 7855
rect 10585 7665 10645 7855
rect 10985 7665 11045 7855
rect 11385 7665 11445 7855
rect 11785 7665 11845 7855
rect 12185 7665 12245 7855
rect 12585 7665 12645 7855
rect 12985 7665 13045 7855
rect -225 7660 -145 7665
rect -225 7600 -215 7660
rect -155 7600 -145 7660
rect -225 7550 -145 7600
rect -225 7490 -215 7550
rect -155 7490 -145 7550
rect -225 7485 -145 7490
rect 175 7660 255 7665
rect 175 7600 185 7660
rect 245 7600 255 7660
rect 175 7550 255 7600
rect 175 7490 185 7550
rect 245 7490 255 7550
rect 175 7485 255 7490
rect 575 7660 655 7665
rect 575 7600 585 7660
rect 645 7600 655 7660
rect 575 7550 655 7600
rect 575 7490 585 7550
rect 645 7490 655 7550
rect 575 7485 655 7490
rect 975 7660 1055 7665
rect 975 7600 985 7660
rect 1045 7600 1055 7660
rect 975 7550 1055 7600
rect 975 7490 985 7550
rect 1045 7490 1055 7550
rect 975 7485 1055 7490
rect 1375 7660 1455 7665
rect 1375 7600 1385 7660
rect 1445 7600 1455 7660
rect 1375 7550 1455 7600
rect 1375 7490 1385 7550
rect 1445 7490 1455 7550
rect 1375 7485 1455 7490
rect 1775 7660 1855 7665
rect 1775 7600 1785 7660
rect 1845 7600 1855 7660
rect 1775 7550 1855 7600
rect 1775 7490 1785 7550
rect 1845 7490 1855 7550
rect 1775 7485 1855 7490
rect 2175 7660 2255 7665
rect 2175 7600 2185 7660
rect 2245 7600 2255 7660
rect 2175 7550 2255 7600
rect 2175 7490 2185 7550
rect 2245 7490 2255 7550
rect 2175 7485 2255 7490
rect 2575 7660 2655 7665
rect 2575 7600 2585 7660
rect 2645 7600 2655 7660
rect 2575 7550 2655 7600
rect 2575 7490 2585 7550
rect 2645 7490 2655 7550
rect 2575 7485 2655 7490
rect 2975 7660 3055 7665
rect 2975 7600 2985 7660
rect 3045 7600 3055 7660
rect 2975 7550 3055 7600
rect 2975 7490 2985 7550
rect 3045 7490 3055 7550
rect 2975 7485 3055 7490
rect 3375 7660 3455 7665
rect 3375 7600 3385 7660
rect 3445 7600 3455 7660
rect 3375 7550 3455 7600
rect 3375 7490 3385 7550
rect 3445 7490 3455 7550
rect 3375 7485 3455 7490
rect 3775 7660 3855 7665
rect 3775 7600 3785 7660
rect 3845 7600 3855 7660
rect 3775 7550 3855 7600
rect 3775 7490 3785 7550
rect 3845 7490 3855 7550
rect 3775 7485 3855 7490
rect 4175 7660 4255 7665
rect 4175 7600 4185 7660
rect 4245 7600 4255 7660
rect 4175 7550 4255 7600
rect 4175 7490 4185 7550
rect 4245 7490 4255 7550
rect 4175 7485 4255 7490
rect 4575 7660 4655 7665
rect 4575 7600 4585 7660
rect 4645 7600 4655 7660
rect 4575 7550 4655 7600
rect 4575 7490 4585 7550
rect 4645 7490 4655 7550
rect 4575 7485 4655 7490
rect 4975 7660 5055 7665
rect 4975 7600 4985 7660
rect 5045 7600 5055 7660
rect 4975 7550 5055 7600
rect 4975 7490 4985 7550
rect 5045 7490 5055 7550
rect 4975 7485 5055 7490
rect 5375 7660 5455 7665
rect 5375 7600 5385 7660
rect 5445 7600 5455 7660
rect 5375 7550 5455 7600
rect 5375 7490 5385 7550
rect 5445 7490 5455 7550
rect 5375 7485 5455 7490
rect 5775 7660 5855 7665
rect 5775 7600 5785 7660
rect 5845 7600 5855 7660
rect 5775 7550 5855 7600
rect 5775 7490 5785 7550
rect 5845 7490 5855 7550
rect 5775 7485 5855 7490
rect 6175 7660 6255 7665
rect 6175 7600 6185 7660
rect 6245 7600 6255 7660
rect 6175 7550 6255 7600
rect 6175 7490 6185 7550
rect 6245 7490 6255 7550
rect 6175 7485 6255 7490
rect 6575 7660 6655 7665
rect 6575 7600 6585 7660
rect 6645 7600 6655 7660
rect 6575 7550 6655 7600
rect 6575 7490 6585 7550
rect 6645 7490 6655 7550
rect 6575 7485 6655 7490
rect 6975 7660 7055 7665
rect 6975 7600 6985 7660
rect 7045 7600 7055 7660
rect 6975 7550 7055 7600
rect 6975 7490 6985 7550
rect 7045 7490 7055 7550
rect 6975 7485 7055 7490
rect 7375 7660 7455 7665
rect 7375 7600 7385 7660
rect 7445 7600 7455 7660
rect 7375 7550 7455 7600
rect 7375 7490 7385 7550
rect 7445 7490 7455 7550
rect 7375 7485 7455 7490
rect 7775 7660 7855 7665
rect 7775 7600 7785 7660
rect 7845 7600 7855 7660
rect 7775 7550 7855 7600
rect 7775 7490 7785 7550
rect 7845 7490 7855 7550
rect 7775 7485 7855 7490
rect 8175 7660 8255 7665
rect 8175 7600 8185 7660
rect 8245 7600 8255 7660
rect 8175 7550 8255 7600
rect 8175 7490 8185 7550
rect 8245 7490 8255 7550
rect 8175 7485 8255 7490
rect 8575 7660 8655 7665
rect 8575 7600 8585 7660
rect 8645 7600 8655 7660
rect 8575 7550 8655 7600
rect 8575 7490 8585 7550
rect 8645 7490 8655 7550
rect 8575 7485 8655 7490
rect 8975 7660 9055 7665
rect 8975 7600 8985 7660
rect 9045 7600 9055 7660
rect 8975 7550 9055 7600
rect 8975 7490 8985 7550
rect 9045 7490 9055 7550
rect 8975 7485 9055 7490
rect 9375 7660 9455 7665
rect 9375 7600 9385 7660
rect 9445 7600 9455 7660
rect 9375 7550 9455 7600
rect 9375 7490 9385 7550
rect 9445 7490 9455 7550
rect 9375 7485 9455 7490
rect 9775 7660 9855 7665
rect 9775 7600 9785 7660
rect 9845 7600 9855 7660
rect 9775 7550 9855 7600
rect 9775 7490 9785 7550
rect 9845 7490 9855 7550
rect 9775 7485 9855 7490
rect 10175 7660 10255 7665
rect 10175 7600 10185 7660
rect 10245 7600 10255 7660
rect 10175 7550 10255 7600
rect 10175 7490 10185 7550
rect 10245 7490 10255 7550
rect 10175 7485 10255 7490
rect 10575 7660 10655 7665
rect 10575 7600 10585 7660
rect 10645 7600 10655 7660
rect 10575 7550 10655 7600
rect 10575 7490 10585 7550
rect 10645 7490 10655 7550
rect 10575 7485 10655 7490
rect 10975 7660 11055 7665
rect 10975 7600 10985 7660
rect 11045 7600 11055 7660
rect 10975 7550 11055 7600
rect 10975 7490 10985 7550
rect 11045 7490 11055 7550
rect 10975 7485 11055 7490
rect 11375 7660 11455 7665
rect 11375 7600 11385 7660
rect 11445 7600 11455 7660
rect 11375 7550 11455 7600
rect 11375 7490 11385 7550
rect 11445 7490 11455 7550
rect 11375 7485 11455 7490
rect 11775 7660 11855 7665
rect 11775 7600 11785 7660
rect 11845 7600 11855 7660
rect 11775 7550 11855 7600
rect 11775 7490 11785 7550
rect 11845 7490 11855 7550
rect 11775 7485 11855 7490
rect 12175 7660 12255 7665
rect 12175 7600 12185 7660
rect 12245 7600 12255 7660
rect 12175 7550 12255 7600
rect 12175 7490 12185 7550
rect 12245 7490 12255 7550
rect 12175 7485 12255 7490
rect 12575 7660 12655 7665
rect 12575 7600 12585 7660
rect 12645 7600 12655 7660
rect 12575 7550 12655 7600
rect 12575 7490 12585 7550
rect 12645 7490 12655 7550
rect 12575 7485 12655 7490
rect 12975 7660 13055 7665
rect 12975 7600 12985 7660
rect 13045 7600 13055 7660
rect 12975 7550 13055 7600
rect 12975 7490 12985 7550
rect 13045 7490 13055 7550
rect 12975 7485 13055 7490
rect -215 7295 -155 7485
rect 185 7295 245 7485
rect 585 7295 645 7485
rect 985 7295 1045 7485
rect 1385 7295 1445 7485
rect 1785 7295 1845 7485
rect 2185 7295 2245 7485
rect 2585 7295 2645 7485
rect 2985 7295 3045 7485
rect 3385 7295 3445 7485
rect 3785 7295 3845 7485
rect 4185 7295 4245 7485
rect 4585 7295 4645 7485
rect 4985 7295 5045 7485
rect 5385 7295 5445 7485
rect 5785 7295 5845 7485
rect 6185 7295 6245 7485
rect 6585 7295 6645 7485
rect 6985 7295 7045 7485
rect 7385 7295 7445 7485
rect 7785 7295 7845 7485
rect 8185 7295 8245 7485
rect 8585 7295 8645 7485
rect 8985 7295 9045 7485
rect 9385 7295 9445 7485
rect 9785 7295 9845 7485
rect 10185 7295 10245 7485
rect 10585 7295 10645 7485
rect 10985 7295 11045 7485
rect 11385 7295 11445 7485
rect 11785 7295 11845 7485
rect 12185 7295 12245 7485
rect 12585 7295 12645 7485
rect 12985 7295 13045 7485
rect -225 7290 -145 7295
rect -225 7230 -215 7290
rect -155 7230 -145 7290
rect -225 7180 -145 7230
rect -225 7120 -215 7180
rect -155 7120 -145 7180
rect -225 7115 -145 7120
rect 175 7290 255 7295
rect 175 7230 185 7290
rect 245 7230 255 7290
rect 175 7180 255 7230
rect 175 7120 185 7180
rect 245 7120 255 7180
rect 175 7115 255 7120
rect 575 7290 655 7295
rect 575 7230 585 7290
rect 645 7230 655 7290
rect 575 7180 655 7230
rect 575 7120 585 7180
rect 645 7120 655 7180
rect 575 7115 655 7120
rect 975 7290 1055 7295
rect 975 7230 985 7290
rect 1045 7230 1055 7290
rect 975 7180 1055 7230
rect 975 7120 985 7180
rect 1045 7120 1055 7180
rect 975 7115 1055 7120
rect 1375 7290 1455 7295
rect 1375 7230 1385 7290
rect 1445 7230 1455 7290
rect 1375 7180 1455 7230
rect 1375 7120 1385 7180
rect 1445 7120 1455 7180
rect 1375 7115 1455 7120
rect 1775 7290 1855 7295
rect 1775 7230 1785 7290
rect 1845 7230 1855 7290
rect 1775 7180 1855 7230
rect 1775 7120 1785 7180
rect 1845 7120 1855 7180
rect 1775 7115 1855 7120
rect 2175 7290 2255 7295
rect 2175 7230 2185 7290
rect 2245 7230 2255 7290
rect 2175 7180 2255 7230
rect 2175 7120 2185 7180
rect 2245 7120 2255 7180
rect 2175 7115 2255 7120
rect 2575 7290 2655 7295
rect 2575 7230 2585 7290
rect 2645 7230 2655 7290
rect 2575 7180 2655 7230
rect 2575 7120 2585 7180
rect 2645 7120 2655 7180
rect 2575 7115 2655 7120
rect 2975 7290 3055 7295
rect 2975 7230 2985 7290
rect 3045 7230 3055 7290
rect 2975 7180 3055 7230
rect 2975 7120 2985 7180
rect 3045 7120 3055 7180
rect 2975 7115 3055 7120
rect 3375 7290 3455 7295
rect 3375 7230 3385 7290
rect 3445 7230 3455 7290
rect 3375 7180 3455 7230
rect 3375 7120 3385 7180
rect 3445 7120 3455 7180
rect 3375 7115 3455 7120
rect 3775 7290 3855 7295
rect 3775 7230 3785 7290
rect 3845 7230 3855 7290
rect 3775 7180 3855 7230
rect 3775 7120 3785 7180
rect 3845 7120 3855 7180
rect 3775 7115 3855 7120
rect 4175 7290 4255 7295
rect 4175 7230 4185 7290
rect 4245 7230 4255 7290
rect 4175 7180 4255 7230
rect 4175 7120 4185 7180
rect 4245 7120 4255 7180
rect 4175 7115 4255 7120
rect 4575 7290 4655 7295
rect 4575 7230 4585 7290
rect 4645 7230 4655 7290
rect 4575 7180 4655 7230
rect 4575 7120 4585 7180
rect 4645 7120 4655 7180
rect 4575 7115 4655 7120
rect 4975 7290 5055 7295
rect 4975 7230 4985 7290
rect 5045 7230 5055 7290
rect 4975 7180 5055 7230
rect 4975 7120 4985 7180
rect 5045 7120 5055 7180
rect 4975 7115 5055 7120
rect 5375 7290 5455 7295
rect 5375 7230 5385 7290
rect 5445 7230 5455 7290
rect 5375 7180 5455 7230
rect 5375 7120 5385 7180
rect 5445 7120 5455 7180
rect 5375 7115 5455 7120
rect 5775 7290 5855 7295
rect 5775 7230 5785 7290
rect 5845 7230 5855 7290
rect 5775 7180 5855 7230
rect 5775 7120 5785 7180
rect 5845 7120 5855 7180
rect 5775 7115 5855 7120
rect 6175 7290 6255 7295
rect 6175 7230 6185 7290
rect 6245 7230 6255 7290
rect 6175 7180 6255 7230
rect 6175 7120 6185 7180
rect 6245 7120 6255 7180
rect 6175 7115 6255 7120
rect 6575 7290 6655 7295
rect 6575 7230 6585 7290
rect 6645 7230 6655 7290
rect 6575 7180 6655 7230
rect 6575 7120 6585 7180
rect 6645 7120 6655 7180
rect 6575 7115 6655 7120
rect 6975 7290 7055 7295
rect 6975 7230 6985 7290
rect 7045 7230 7055 7290
rect 6975 7180 7055 7230
rect 6975 7120 6985 7180
rect 7045 7120 7055 7180
rect 6975 7115 7055 7120
rect 7375 7290 7455 7295
rect 7375 7230 7385 7290
rect 7445 7230 7455 7290
rect 7375 7180 7455 7230
rect 7375 7120 7385 7180
rect 7445 7120 7455 7180
rect 7375 7115 7455 7120
rect 7775 7290 7855 7295
rect 7775 7230 7785 7290
rect 7845 7230 7855 7290
rect 7775 7180 7855 7230
rect 7775 7120 7785 7180
rect 7845 7120 7855 7180
rect 7775 7115 7855 7120
rect 8175 7290 8255 7295
rect 8175 7230 8185 7290
rect 8245 7230 8255 7290
rect 8175 7180 8255 7230
rect 8175 7120 8185 7180
rect 8245 7120 8255 7180
rect 8175 7115 8255 7120
rect 8575 7290 8655 7295
rect 8575 7230 8585 7290
rect 8645 7230 8655 7290
rect 8575 7180 8655 7230
rect 8575 7120 8585 7180
rect 8645 7120 8655 7180
rect 8575 7115 8655 7120
rect 8975 7290 9055 7295
rect 8975 7230 8985 7290
rect 9045 7230 9055 7290
rect 8975 7180 9055 7230
rect 8975 7120 8985 7180
rect 9045 7120 9055 7180
rect 8975 7115 9055 7120
rect 9375 7290 9455 7295
rect 9375 7230 9385 7290
rect 9445 7230 9455 7290
rect 9375 7180 9455 7230
rect 9375 7120 9385 7180
rect 9445 7120 9455 7180
rect 9375 7115 9455 7120
rect 9775 7290 9855 7295
rect 9775 7230 9785 7290
rect 9845 7230 9855 7290
rect 9775 7180 9855 7230
rect 9775 7120 9785 7180
rect 9845 7120 9855 7180
rect 9775 7115 9855 7120
rect 10175 7290 10255 7295
rect 10175 7230 10185 7290
rect 10245 7230 10255 7290
rect 10175 7180 10255 7230
rect 10175 7120 10185 7180
rect 10245 7120 10255 7180
rect 10175 7115 10255 7120
rect 10575 7290 10655 7295
rect 10575 7230 10585 7290
rect 10645 7230 10655 7290
rect 10575 7180 10655 7230
rect 10575 7120 10585 7180
rect 10645 7120 10655 7180
rect 10575 7115 10655 7120
rect 10975 7290 11055 7295
rect 10975 7230 10985 7290
rect 11045 7230 11055 7290
rect 10975 7180 11055 7230
rect 10975 7120 10985 7180
rect 11045 7120 11055 7180
rect 10975 7115 11055 7120
rect 11375 7290 11455 7295
rect 11375 7230 11385 7290
rect 11445 7230 11455 7290
rect 11375 7180 11455 7230
rect 11375 7120 11385 7180
rect 11445 7120 11455 7180
rect 11375 7115 11455 7120
rect 11775 7290 11855 7295
rect 11775 7230 11785 7290
rect 11845 7230 11855 7290
rect 11775 7180 11855 7230
rect 11775 7120 11785 7180
rect 11845 7120 11855 7180
rect 11775 7115 11855 7120
rect 12175 7290 12255 7295
rect 12175 7230 12185 7290
rect 12245 7230 12255 7290
rect 12175 7180 12255 7230
rect 12175 7120 12185 7180
rect 12245 7120 12255 7180
rect 12175 7115 12255 7120
rect 12575 7290 12655 7295
rect 12575 7230 12585 7290
rect 12645 7230 12655 7290
rect 12575 7180 12655 7230
rect 12575 7120 12585 7180
rect 12645 7120 12655 7180
rect 12575 7115 12655 7120
rect 12975 7290 13055 7295
rect 12975 7230 12985 7290
rect 13045 7230 13055 7290
rect 12975 7180 13055 7230
rect 12975 7120 12985 7180
rect 13045 7120 13055 7180
rect 12975 7115 13055 7120
rect -215 6925 -155 7115
rect 185 6925 245 7115
rect 585 6925 645 7115
rect 985 6925 1045 7115
rect 1385 6925 1445 7115
rect 1785 6925 1845 7115
rect 2185 6925 2245 7115
rect 2585 6925 2645 7115
rect 2985 6925 3045 7115
rect 3385 6925 3445 7115
rect 3785 6925 3845 7115
rect 4185 6925 4245 7115
rect 4585 6925 4645 7115
rect 4985 6925 5045 7115
rect 5385 6925 5445 7115
rect 5785 6925 5845 7115
rect 6185 6925 6245 7115
rect 6585 6925 6645 7115
rect 6985 6925 7045 7115
rect 7385 6925 7445 7115
rect 7785 6925 7845 7115
rect 8185 6925 8245 7115
rect 8585 6925 8645 7115
rect 8985 6925 9045 7115
rect 9385 6925 9445 7115
rect 9785 6925 9845 7115
rect 10185 6925 10245 7115
rect 10585 6925 10645 7115
rect 10985 6925 11045 7115
rect 11385 6925 11445 7115
rect 11785 6925 11845 7115
rect 12185 6925 12245 7115
rect 12585 6925 12645 7115
rect 12985 6925 13045 7115
rect -225 6920 -145 6925
rect -225 6860 -215 6920
rect -155 6860 -145 6920
rect -225 6810 -145 6860
rect -225 6750 -215 6810
rect -155 6750 -145 6810
rect -225 6745 -145 6750
rect 175 6920 255 6925
rect 175 6860 185 6920
rect 245 6860 255 6920
rect 175 6810 255 6860
rect 175 6750 185 6810
rect 245 6750 255 6810
rect 175 6745 255 6750
rect 575 6920 655 6925
rect 575 6860 585 6920
rect 645 6860 655 6920
rect 575 6810 655 6860
rect 575 6750 585 6810
rect 645 6750 655 6810
rect 575 6745 655 6750
rect 975 6920 1055 6925
rect 975 6860 985 6920
rect 1045 6860 1055 6920
rect 975 6810 1055 6860
rect 975 6750 985 6810
rect 1045 6750 1055 6810
rect 975 6745 1055 6750
rect 1375 6920 1455 6925
rect 1375 6860 1385 6920
rect 1445 6860 1455 6920
rect 1375 6810 1455 6860
rect 1375 6750 1385 6810
rect 1445 6750 1455 6810
rect 1375 6745 1455 6750
rect 1775 6920 1855 6925
rect 1775 6860 1785 6920
rect 1845 6860 1855 6920
rect 1775 6810 1855 6860
rect 1775 6750 1785 6810
rect 1845 6750 1855 6810
rect 1775 6745 1855 6750
rect 2175 6920 2255 6925
rect 2175 6860 2185 6920
rect 2245 6860 2255 6920
rect 2175 6810 2255 6860
rect 2175 6750 2185 6810
rect 2245 6750 2255 6810
rect 2175 6745 2255 6750
rect 2575 6920 2655 6925
rect 2575 6860 2585 6920
rect 2645 6860 2655 6920
rect 2575 6810 2655 6860
rect 2575 6750 2585 6810
rect 2645 6750 2655 6810
rect 2575 6745 2655 6750
rect 2975 6920 3055 6925
rect 2975 6860 2985 6920
rect 3045 6860 3055 6920
rect 2975 6810 3055 6860
rect 2975 6750 2985 6810
rect 3045 6750 3055 6810
rect 2975 6745 3055 6750
rect 3375 6920 3455 6925
rect 3375 6860 3385 6920
rect 3445 6860 3455 6920
rect 3375 6810 3455 6860
rect 3375 6750 3385 6810
rect 3445 6750 3455 6810
rect 3375 6745 3455 6750
rect 3775 6920 3855 6925
rect 3775 6860 3785 6920
rect 3845 6860 3855 6920
rect 3775 6810 3855 6860
rect 3775 6750 3785 6810
rect 3845 6750 3855 6810
rect 3775 6745 3855 6750
rect 4175 6920 4255 6925
rect 4175 6860 4185 6920
rect 4245 6860 4255 6920
rect 4175 6810 4255 6860
rect 4175 6750 4185 6810
rect 4245 6750 4255 6810
rect 4175 6745 4255 6750
rect 4575 6920 4655 6925
rect 4575 6860 4585 6920
rect 4645 6860 4655 6920
rect 4575 6810 4655 6860
rect 4575 6750 4585 6810
rect 4645 6750 4655 6810
rect 4575 6745 4655 6750
rect 4975 6920 5055 6925
rect 4975 6860 4985 6920
rect 5045 6860 5055 6920
rect 4975 6810 5055 6860
rect 4975 6750 4985 6810
rect 5045 6750 5055 6810
rect 4975 6745 5055 6750
rect 5375 6920 5455 6925
rect 5375 6860 5385 6920
rect 5445 6860 5455 6920
rect 5375 6810 5455 6860
rect 5375 6750 5385 6810
rect 5445 6750 5455 6810
rect 5375 6745 5455 6750
rect 5775 6920 5855 6925
rect 5775 6860 5785 6920
rect 5845 6860 5855 6920
rect 5775 6810 5855 6860
rect 5775 6750 5785 6810
rect 5845 6750 5855 6810
rect 5775 6745 5855 6750
rect 6175 6920 6255 6925
rect 6175 6860 6185 6920
rect 6245 6860 6255 6920
rect 6175 6810 6255 6860
rect 6175 6750 6185 6810
rect 6245 6750 6255 6810
rect 6175 6745 6255 6750
rect 6575 6920 6655 6925
rect 6575 6860 6585 6920
rect 6645 6860 6655 6920
rect 6575 6810 6655 6860
rect 6575 6750 6585 6810
rect 6645 6750 6655 6810
rect 6575 6745 6655 6750
rect 6975 6920 7055 6925
rect 6975 6860 6985 6920
rect 7045 6860 7055 6920
rect 6975 6810 7055 6860
rect 6975 6750 6985 6810
rect 7045 6750 7055 6810
rect 6975 6745 7055 6750
rect 7375 6920 7455 6925
rect 7375 6860 7385 6920
rect 7445 6860 7455 6920
rect 7375 6810 7455 6860
rect 7375 6750 7385 6810
rect 7445 6750 7455 6810
rect 7375 6745 7455 6750
rect 7775 6920 7855 6925
rect 7775 6860 7785 6920
rect 7845 6860 7855 6920
rect 7775 6810 7855 6860
rect 7775 6750 7785 6810
rect 7845 6750 7855 6810
rect 7775 6745 7855 6750
rect 8175 6920 8255 6925
rect 8175 6860 8185 6920
rect 8245 6860 8255 6920
rect 8175 6810 8255 6860
rect 8175 6750 8185 6810
rect 8245 6750 8255 6810
rect 8175 6745 8255 6750
rect 8575 6920 8655 6925
rect 8575 6860 8585 6920
rect 8645 6860 8655 6920
rect 8575 6810 8655 6860
rect 8575 6750 8585 6810
rect 8645 6750 8655 6810
rect 8575 6745 8655 6750
rect 8975 6920 9055 6925
rect 8975 6860 8985 6920
rect 9045 6860 9055 6920
rect 8975 6810 9055 6860
rect 8975 6750 8985 6810
rect 9045 6750 9055 6810
rect 8975 6745 9055 6750
rect 9375 6920 9455 6925
rect 9375 6860 9385 6920
rect 9445 6860 9455 6920
rect 9375 6810 9455 6860
rect 9375 6750 9385 6810
rect 9445 6750 9455 6810
rect 9375 6745 9455 6750
rect 9775 6920 9855 6925
rect 9775 6860 9785 6920
rect 9845 6860 9855 6920
rect 9775 6810 9855 6860
rect 9775 6750 9785 6810
rect 9845 6750 9855 6810
rect 9775 6745 9855 6750
rect 10175 6920 10255 6925
rect 10175 6860 10185 6920
rect 10245 6860 10255 6920
rect 10175 6810 10255 6860
rect 10175 6750 10185 6810
rect 10245 6750 10255 6810
rect 10175 6745 10255 6750
rect 10575 6920 10655 6925
rect 10575 6860 10585 6920
rect 10645 6860 10655 6920
rect 10575 6810 10655 6860
rect 10575 6750 10585 6810
rect 10645 6750 10655 6810
rect 10575 6745 10655 6750
rect 10975 6920 11055 6925
rect 10975 6860 10985 6920
rect 11045 6860 11055 6920
rect 10975 6810 11055 6860
rect 10975 6750 10985 6810
rect 11045 6750 11055 6810
rect 10975 6745 11055 6750
rect 11375 6920 11455 6925
rect 11375 6860 11385 6920
rect 11445 6860 11455 6920
rect 11375 6810 11455 6860
rect 11375 6750 11385 6810
rect 11445 6750 11455 6810
rect 11375 6745 11455 6750
rect 11775 6920 11855 6925
rect 11775 6860 11785 6920
rect 11845 6860 11855 6920
rect 11775 6810 11855 6860
rect 11775 6750 11785 6810
rect 11845 6750 11855 6810
rect 11775 6745 11855 6750
rect 12175 6920 12255 6925
rect 12175 6860 12185 6920
rect 12245 6860 12255 6920
rect 12175 6810 12255 6860
rect 12175 6750 12185 6810
rect 12245 6750 12255 6810
rect 12175 6745 12255 6750
rect 12575 6920 12655 6925
rect 12575 6860 12585 6920
rect 12645 6860 12655 6920
rect 12575 6810 12655 6860
rect 12575 6750 12585 6810
rect 12645 6750 12655 6810
rect 12575 6745 12655 6750
rect 12975 6920 13055 6925
rect 12975 6860 12985 6920
rect 13045 6860 13055 6920
rect 12975 6810 13055 6860
rect 12975 6750 12985 6810
rect 13045 6750 13055 6810
rect 12975 6745 13055 6750
rect -215 6555 -155 6745
rect 185 6555 245 6745
rect 585 6555 645 6745
rect 985 6555 1045 6745
rect 1385 6555 1445 6745
rect 1785 6555 1845 6745
rect 2185 6555 2245 6745
rect 2585 6555 2645 6745
rect 2985 6555 3045 6745
rect 3385 6555 3445 6745
rect 3785 6555 3845 6745
rect 4185 6555 4245 6745
rect 4585 6555 4645 6745
rect 4985 6555 5045 6745
rect 5385 6555 5445 6745
rect 5785 6555 5845 6745
rect 6185 6555 6245 6745
rect 6585 6555 6645 6745
rect 6985 6555 7045 6745
rect 7385 6555 7445 6745
rect 7785 6555 7845 6745
rect 8185 6555 8245 6745
rect 8585 6555 8645 6745
rect 8985 6555 9045 6745
rect 9385 6555 9445 6745
rect 9785 6555 9845 6745
rect 10185 6555 10245 6745
rect 10585 6555 10645 6745
rect 10985 6555 11045 6745
rect 11385 6555 11445 6745
rect 11785 6555 11845 6745
rect 12185 6555 12245 6745
rect 12585 6555 12645 6745
rect 12985 6555 13045 6745
rect -225 6550 -145 6555
rect -225 6490 -215 6550
rect -155 6490 -145 6550
rect -225 6440 -145 6490
rect -225 6380 -215 6440
rect -155 6380 -145 6440
rect -225 6375 -145 6380
rect 175 6550 255 6555
rect 175 6490 185 6550
rect 245 6490 255 6550
rect 175 6440 255 6490
rect 175 6380 185 6440
rect 245 6380 255 6440
rect 175 6375 255 6380
rect 575 6550 655 6555
rect 575 6490 585 6550
rect 645 6490 655 6550
rect 575 6440 655 6490
rect 575 6380 585 6440
rect 645 6380 655 6440
rect 575 6375 655 6380
rect 975 6550 1055 6555
rect 975 6490 985 6550
rect 1045 6490 1055 6550
rect 975 6440 1055 6490
rect 975 6380 985 6440
rect 1045 6380 1055 6440
rect 975 6375 1055 6380
rect 1375 6550 1455 6555
rect 1375 6490 1385 6550
rect 1445 6490 1455 6550
rect 1375 6440 1455 6490
rect 1375 6380 1385 6440
rect 1445 6380 1455 6440
rect 1375 6375 1455 6380
rect 1775 6550 1855 6555
rect 1775 6490 1785 6550
rect 1845 6490 1855 6550
rect 1775 6440 1855 6490
rect 1775 6380 1785 6440
rect 1845 6380 1855 6440
rect 1775 6375 1855 6380
rect 2175 6550 2255 6555
rect 2175 6490 2185 6550
rect 2245 6490 2255 6550
rect 2175 6440 2255 6490
rect 2175 6380 2185 6440
rect 2245 6380 2255 6440
rect 2175 6375 2255 6380
rect 2575 6550 2655 6555
rect 2575 6490 2585 6550
rect 2645 6490 2655 6550
rect 2575 6440 2655 6490
rect 2575 6380 2585 6440
rect 2645 6380 2655 6440
rect 2575 6375 2655 6380
rect 2975 6550 3055 6555
rect 2975 6490 2985 6550
rect 3045 6490 3055 6550
rect 2975 6440 3055 6490
rect 2975 6380 2985 6440
rect 3045 6380 3055 6440
rect 2975 6375 3055 6380
rect 3375 6550 3455 6555
rect 3375 6490 3385 6550
rect 3445 6490 3455 6550
rect 3375 6440 3455 6490
rect 3375 6380 3385 6440
rect 3445 6380 3455 6440
rect 3375 6375 3455 6380
rect 3775 6550 3855 6555
rect 3775 6490 3785 6550
rect 3845 6490 3855 6550
rect 3775 6440 3855 6490
rect 3775 6380 3785 6440
rect 3845 6380 3855 6440
rect 3775 6375 3855 6380
rect 4175 6550 4255 6555
rect 4175 6490 4185 6550
rect 4245 6490 4255 6550
rect 4175 6440 4255 6490
rect 4175 6380 4185 6440
rect 4245 6380 4255 6440
rect 4175 6375 4255 6380
rect 4575 6550 4655 6555
rect 4575 6490 4585 6550
rect 4645 6490 4655 6550
rect 4575 6440 4655 6490
rect 4575 6380 4585 6440
rect 4645 6380 4655 6440
rect 4575 6375 4655 6380
rect 4975 6550 5055 6555
rect 4975 6490 4985 6550
rect 5045 6490 5055 6550
rect 4975 6440 5055 6490
rect 4975 6380 4985 6440
rect 5045 6380 5055 6440
rect 4975 6375 5055 6380
rect 5375 6550 5455 6555
rect 5375 6490 5385 6550
rect 5445 6490 5455 6550
rect 5375 6440 5455 6490
rect 5375 6380 5385 6440
rect 5445 6380 5455 6440
rect 5375 6375 5455 6380
rect 5775 6550 5855 6555
rect 5775 6490 5785 6550
rect 5845 6490 5855 6550
rect 5775 6440 5855 6490
rect 5775 6380 5785 6440
rect 5845 6380 5855 6440
rect 5775 6375 5855 6380
rect 6175 6550 6255 6555
rect 6175 6490 6185 6550
rect 6245 6490 6255 6550
rect 6175 6440 6255 6490
rect 6175 6380 6185 6440
rect 6245 6380 6255 6440
rect 6175 6375 6255 6380
rect 6575 6550 6655 6555
rect 6575 6490 6585 6550
rect 6645 6490 6655 6550
rect 6575 6440 6655 6490
rect 6575 6380 6585 6440
rect 6645 6380 6655 6440
rect 6575 6375 6655 6380
rect 6975 6550 7055 6555
rect 6975 6490 6985 6550
rect 7045 6490 7055 6550
rect 6975 6440 7055 6490
rect 6975 6380 6985 6440
rect 7045 6380 7055 6440
rect 6975 6375 7055 6380
rect 7375 6550 7455 6555
rect 7375 6490 7385 6550
rect 7445 6490 7455 6550
rect 7375 6440 7455 6490
rect 7375 6380 7385 6440
rect 7445 6380 7455 6440
rect 7375 6375 7455 6380
rect 7775 6550 7855 6555
rect 7775 6490 7785 6550
rect 7845 6490 7855 6550
rect 7775 6440 7855 6490
rect 7775 6380 7785 6440
rect 7845 6380 7855 6440
rect 7775 6375 7855 6380
rect 8175 6550 8255 6555
rect 8175 6490 8185 6550
rect 8245 6490 8255 6550
rect 8175 6440 8255 6490
rect 8175 6380 8185 6440
rect 8245 6380 8255 6440
rect 8175 6375 8255 6380
rect 8575 6550 8655 6555
rect 8575 6490 8585 6550
rect 8645 6490 8655 6550
rect 8575 6440 8655 6490
rect 8575 6380 8585 6440
rect 8645 6380 8655 6440
rect 8575 6375 8655 6380
rect 8975 6550 9055 6555
rect 8975 6490 8985 6550
rect 9045 6490 9055 6550
rect 8975 6440 9055 6490
rect 8975 6380 8985 6440
rect 9045 6380 9055 6440
rect 8975 6375 9055 6380
rect 9375 6550 9455 6555
rect 9375 6490 9385 6550
rect 9445 6490 9455 6550
rect 9375 6440 9455 6490
rect 9375 6380 9385 6440
rect 9445 6380 9455 6440
rect 9375 6375 9455 6380
rect 9775 6550 9855 6555
rect 9775 6490 9785 6550
rect 9845 6490 9855 6550
rect 9775 6440 9855 6490
rect 9775 6380 9785 6440
rect 9845 6380 9855 6440
rect 9775 6375 9855 6380
rect 10175 6550 10255 6555
rect 10175 6490 10185 6550
rect 10245 6490 10255 6550
rect 10175 6440 10255 6490
rect 10175 6380 10185 6440
rect 10245 6380 10255 6440
rect 10175 6375 10255 6380
rect 10575 6550 10655 6555
rect 10575 6490 10585 6550
rect 10645 6490 10655 6550
rect 10575 6440 10655 6490
rect 10575 6380 10585 6440
rect 10645 6380 10655 6440
rect 10575 6375 10655 6380
rect 10975 6550 11055 6555
rect 10975 6490 10985 6550
rect 11045 6490 11055 6550
rect 10975 6440 11055 6490
rect 10975 6380 10985 6440
rect 11045 6380 11055 6440
rect 10975 6375 11055 6380
rect 11375 6550 11455 6555
rect 11375 6490 11385 6550
rect 11445 6490 11455 6550
rect 11375 6440 11455 6490
rect 11375 6380 11385 6440
rect 11445 6380 11455 6440
rect 11375 6375 11455 6380
rect 11775 6550 11855 6555
rect 11775 6490 11785 6550
rect 11845 6490 11855 6550
rect 11775 6440 11855 6490
rect 11775 6380 11785 6440
rect 11845 6380 11855 6440
rect 11775 6375 11855 6380
rect 12175 6550 12255 6555
rect 12175 6490 12185 6550
rect 12245 6490 12255 6550
rect 12175 6440 12255 6490
rect 12175 6380 12185 6440
rect 12245 6380 12255 6440
rect 12175 6375 12255 6380
rect 12575 6550 12655 6555
rect 12575 6490 12585 6550
rect 12645 6490 12655 6550
rect 12575 6440 12655 6490
rect 12575 6380 12585 6440
rect 12645 6380 12655 6440
rect 12575 6375 12655 6380
rect 12975 6550 13055 6555
rect 12975 6490 12985 6550
rect 13045 6490 13055 6550
rect 12975 6440 13055 6490
rect 12975 6380 12985 6440
rect 13045 6380 13055 6440
rect 12975 6375 13055 6380
rect -215 6185 -155 6375
rect 185 6185 245 6375
rect 585 6185 645 6375
rect 985 6185 1045 6375
rect 1385 6185 1445 6375
rect 1785 6185 1845 6375
rect 2185 6185 2245 6375
rect 2585 6185 2645 6375
rect 2985 6185 3045 6375
rect 3385 6185 3445 6375
rect 3785 6185 3845 6375
rect 4185 6185 4245 6375
rect 4585 6185 4645 6375
rect 4985 6185 5045 6375
rect 5385 6185 5445 6375
rect 5785 6185 5845 6375
rect 6185 6185 6245 6375
rect 6585 6185 6645 6375
rect 6985 6185 7045 6375
rect 7385 6185 7445 6375
rect 7785 6185 7845 6375
rect 8185 6185 8245 6375
rect 8585 6185 8645 6375
rect 8985 6185 9045 6375
rect 9385 6185 9445 6375
rect 9785 6185 9845 6375
rect 10185 6185 10245 6375
rect 10585 6185 10645 6375
rect 10985 6185 11045 6375
rect 11385 6185 11445 6375
rect 11785 6185 11845 6375
rect 12185 6185 12245 6375
rect 12585 6185 12645 6375
rect 12985 6185 13045 6375
rect -225 6180 -145 6185
rect -225 6120 -215 6180
rect -155 6120 -145 6180
rect -225 6070 -145 6120
rect -225 6010 -215 6070
rect -155 6010 -145 6070
rect -225 6005 -145 6010
rect 175 6180 255 6185
rect 175 6120 185 6180
rect 245 6120 255 6180
rect 175 6070 255 6120
rect 175 6010 185 6070
rect 245 6010 255 6070
rect 175 6005 255 6010
rect 575 6180 655 6185
rect 575 6120 585 6180
rect 645 6120 655 6180
rect 575 6070 655 6120
rect 575 6010 585 6070
rect 645 6010 655 6070
rect 575 6005 655 6010
rect 975 6180 1055 6185
rect 975 6120 985 6180
rect 1045 6120 1055 6180
rect 975 6070 1055 6120
rect 975 6010 985 6070
rect 1045 6010 1055 6070
rect 975 6005 1055 6010
rect 1375 6180 1455 6185
rect 1375 6120 1385 6180
rect 1445 6120 1455 6180
rect 1375 6070 1455 6120
rect 1375 6010 1385 6070
rect 1445 6010 1455 6070
rect 1375 6005 1455 6010
rect 1775 6180 1855 6185
rect 1775 6120 1785 6180
rect 1845 6120 1855 6180
rect 1775 6070 1855 6120
rect 1775 6010 1785 6070
rect 1845 6010 1855 6070
rect 1775 6005 1855 6010
rect 2175 6180 2255 6185
rect 2175 6120 2185 6180
rect 2245 6120 2255 6180
rect 2175 6070 2255 6120
rect 2175 6010 2185 6070
rect 2245 6010 2255 6070
rect 2175 6005 2255 6010
rect 2575 6180 2655 6185
rect 2575 6120 2585 6180
rect 2645 6120 2655 6180
rect 2575 6070 2655 6120
rect 2575 6010 2585 6070
rect 2645 6010 2655 6070
rect 2575 6005 2655 6010
rect 2975 6180 3055 6185
rect 2975 6120 2985 6180
rect 3045 6120 3055 6180
rect 2975 6070 3055 6120
rect 2975 6010 2985 6070
rect 3045 6010 3055 6070
rect 2975 6005 3055 6010
rect 3375 6180 3455 6185
rect 3375 6120 3385 6180
rect 3445 6120 3455 6180
rect 3375 6070 3455 6120
rect 3375 6010 3385 6070
rect 3445 6010 3455 6070
rect 3375 6005 3455 6010
rect 3775 6180 3855 6185
rect 3775 6120 3785 6180
rect 3845 6120 3855 6180
rect 3775 6070 3855 6120
rect 3775 6010 3785 6070
rect 3845 6010 3855 6070
rect 3775 6005 3855 6010
rect 4175 6180 4255 6185
rect 4175 6120 4185 6180
rect 4245 6120 4255 6180
rect 4175 6070 4255 6120
rect 4175 6010 4185 6070
rect 4245 6010 4255 6070
rect 4175 6005 4255 6010
rect 4575 6180 4655 6185
rect 4575 6120 4585 6180
rect 4645 6120 4655 6180
rect 4575 6070 4655 6120
rect 4575 6010 4585 6070
rect 4645 6010 4655 6070
rect 4575 6005 4655 6010
rect 4975 6180 5055 6185
rect 4975 6120 4985 6180
rect 5045 6120 5055 6180
rect 4975 6070 5055 6120
rect 4975 6010 4985 6070
rect 5045 6010 5055 6070
rect 4975 6005 5055 6010
rect 5375 6180 5455 6185
rect 5375 6120 5385 6180
rect 5445 6120 5455 6180
rect 5375 6070 5455 6120
rect 5375 6010 5385 6070
rect 5445 6010 5455 6070
rect 5375 6005 5455 6010
rect 5775 6180 5855 6185
rect 5775 6120 5785 6180
rect 5845 6120 5855 6180
rect 5775 6070 5855 6120
rect 5775 6010 5785 6070
rect 5845 6010 5855 6070
rect 5775 6005 5855 6010
rect 6175 6180 6255 6185
rect 6175 6120 6185 6180
rect 6245 6120 6255 6180
rect 6175 6070 6255 6120
rect 6175 6010 6185 6070
rect 6245 6010 6255 6070
rect 6175 6005 6255 6010
rect 6575 6180 6655 6185
rect 6575 6120 6585 6180
rect 6645 6120 6655 6180
rect 6575 6070 6655 6120
rect 6575 6010 6585 6070
rect 6645 6010 6655 6070
rect 6575 6005 6655 6010
rect 6975 6180 7055 6185
rect 6975 6120 6985 6180
rect 7045 6120 7055 6180
rect 6975 6070 7055 6120
rect 6975 6010 6985 6070
rect 7045 6010 7055 6070
rect 6975 6005 7055 6010
rect 7375 6180 7455 6185
rect 7375 6120 7385 6180
rect 7445 6120 7455 6180
rect 7375 6070 7455 6120
rect 7375 6010 7385 6070
rect 7445 6010 7455 6070
rect 7375 6005 7455 6010
rect 7775 6180 7855 6185
rect 7775 6120 7785 6180
rect 7845 6120 7855 6180
rect 7775 6070 7855 6120
rect 7775 6010 7785 6070
rect 7845 6010 7855 6070
rect 7775 6005 7855 6010
rect 8175 6180 8255 6185
rect 8175 6120 8185 6180
rect 8245 6120 8255 6180
rect 8175 6070 8255 6120
rect 8175 6010 8185 6070
rect 8245 6010 8255 6070
rect 8175 6005 8255 6010
rect 8575 6180 8655 6185
rect 8575 6120 8585 6180
rect 8645 6120 8655 6180
rect 8575 6070 8655 6120
rect 8575 6010 8585 6070
rect 8645 6010 8655 6070
rect 8575 6005 8655 6010
rect 8975 6180 9055 6185
rect 8975 6120 8985 6180
rect 9045 6120 9055 6180
rect 8975 6070 9055 6120
rect 8975 6010 8985 6070
rect 9045 6010 9055 6070
rect 8975 6005 9055 6010
rect 9375 6180 9455 6185
rect 9375 6120 9385 6180
rect 9445 6120 9455 6180
rect 9375 6070 9455 6120
rect 9375 6010 9385 6070
rect 9445 6010 9455 6070
rect 9375 6005 9455 6010
rect 9775 6180 9855 6185
rect 9775 6120 9785 6180
rect 9845 6120 9855 6180
rect 9775 6070 9855 6120
rect 9775 6010 9785 6070
rect 9845 6010 9855 6070
rect 9775 6005 9855 6010
rect 10175 6180 10255 6185
rect 10175 6120 10185 6180
rect 10245 6120 10255 6180
rect 10175 6070 10255 6120
rect 10175 6010 10185 6070
rect 10245 6010 10255 6070
rect 10175 6005 10255 6010
rect 10575 6180 10655 6185
rect 10575 6120 10585 6180
rect 10645 6120 10655 6180
rect 10575 6070 10655 6120
rect 10575 6010 10585 6070
rect 10645 6010 10655 6070
rect 10575 6005 10655 6010
rect 10975 6180 11055 6185
rect 10975 6120 10985 6180
rect 11045 6120 11055 6180
rect 10975 6070 11055 6120
rect 10975 6010 10985 6070
rect 11045 6010 11055 6070
rect 10975 6005 11055 6010
rect 11375 6180 11455 6185
rect 11375 6120 11385 6180
rect 11445 6120 11455 6180
rect 11375 6070 11455 6120
rect 11375 6010 11385 6070
rect 11445 6010 11455 6070
rect 11375 6005 11455 6010
rect 11775 6180 11855 6185
rect 11775 6120 11785 6180
rect 11845 6120 11855 6180
rect 11775 6070 11855 6120
rect 11775 6010 11785 6070
rect 11845 6010 11855 6070
rect 11775 6005 11855 6010
rect 12175 6180 12255 6185
rect 12175 6120 12185 6180
rect 12245 6120 12255 6180
rect 12175 6070 12255 6120
rect 12175 6010 12185 6070
rect 12245 6010 12255 6070
rect 12175 6005 12255 6010
rect 12575 6180 12655 6185
rect 12575 6120 12585 6180
rect 12645 6120 12655 6180
rect 12575 6070 12655 6120
rect 12575 6010 12585 6070
rect 12645 6010 12655 6070
rect 12575 6005 12655 6010
rect 12975 6180 13055 6185
rect 12975 6120 12985 6180
rect 13045 6120 13055 6180
rect 12975 6070 13055 6120
rect 12975 6010 12985 6070
rect 13045 6010 13055 6070
rect 12975 6005 13055 6010
rect -215 5815 -155 6005
rect 185 5815 245 6005
rect 585 5815 645 6005
rect 985 5815 1045 6005
rect 1385 5815 1445 6005
rect 1785 5815 1845 6005
rect 2185 5815 2245 6005
rect 2585 5815 2645 6005
rect 2985 5815 3045 6005
rect 3385 5815 3445 6005
rect 3785 5815 3845 6005
rect 4185 5815 4245 6005
rect 4585 5815 4645 6005
rect 4985 5815 5045 6005
rect 5385 5815 5445 6005
rect 5785 5815 5845 6005
rect 6185 5815 6245 6005
rect 6585 5815 6645 6005
rect 6985 5815 7045 6005
rect 7385 5815 7445 6005
rect 7785 5815 7845 6005
rect 8185 5815 8245 6005
rect 8585 5815 8645 6005
rect 8985 5815 9045 6005
rect 9385 5815 9445 6005
rect 9785 5815 9845 6005
rect 10185 5815 10245 6005
rect 10585 5815 10645 6005
rect 10985 5815 11045 6005
rect 11385 5815 11445 6005
rect 11785 5815 11845 6005
rect 12185 5815 12245 6005
rect 12585 5815 12645 6005
rect 12985 5815 13045 6005
rect -225 5810 -145 5815
rect -225 5750 -215 5810
rect -155 5750 -145 5810
rect -225 5700 -145 5750
rect -225 5640 -215 5700
rect -155 5640 -145 5700
rect -225 5635 -145 5640
rect 175 5810 255 5815
rect 175 5750 185 5810
rect 245 5750 255 5810
rect 175 5700 255 5750
rect 175 5640 185 5700
rect 245 5640 255 5700
rect 175 5635 255 5640
rect 575 5810 655 5815
rect 575 5750 585 5810
rect 645 5750 655 5810
rect 575 5700 655 5750
rect 575 5640 585 5700
rect 645 5640 655 5700
rect 575 5635 655 5640
rect 975 5810 1055 5815
rect 975 5750 985 5810
rect 1045 5750 1055 5810
rect 975 5700 1055 5750
rect 975 5640 985 5700
rect 1045 5640 1055 5700
rect 975 5635 1055 5640
rect 1375 5810 1455 5815
rect 1375 5750 1385 5810
rect 1445 5750 1455 5810
rect 1375 5700 1455 5750
rect 1375 5640 1385 5700
rect 1445 5640 1455 5700
rect 1375 5635 1455 5640
rect 1775 5810 1855 5815
rect 1775 5750 1785 5810
rect 1845 5750 1855 5810
rect 1775 5700 1855 5750
rect 1775 5640 1785 5700
rect 1845 5640 1855 5700
rect 1775 5635 1855 5640
rect 2175 5810 2255 5815
rect 2175 5750 2185 5810
rect 2245 5750 2255 5810
rect 2175 5700 2255 5750
rect 2175 5640 2185 5700
rect 2245 5640 2255 5700
rect 2175 5635 2255 5640
rect 2575 5810 2655 5815
rect 2575 5750 2585 5810
rect 2645 5750 2655 5810
rect 2575 5700 2655 5750
rect 2575 5640 2585 5700
rect 2645 5640 2655 5700
rect 2575 5635 2655 5640
rect 2975 5810 3055 5815
rect 2975 5750 2985 5810
rect 3045 5750 3055 5810
rect 2975 5700 3055 5750
rect 2975 5640 2985 5700
rect 3045 5640 3055 5700
rect 2975 5635 3055 5640
rect 3375 5810 3455 5815
rect 3375 5750 3385 5810
rect 3445 5750 3455 5810
rect 3375 5700 3455 5750
rect 3375 5640 3385 5700
rect 3445 5640 3455 5700
rect 3375 5635 3455 5640
rect 3775 5810 3855 5815
rect 3775 5750 3785 5810
rect 3845 5750 3855 5810
rect 3775 5700 3855 5750
rect 3775 5640 3785 5700
rect 3845 5640 3855 5700
rect 3775 5635 3855 5640
rect 4175 5810 4255 5815
rect 4175 5750 4185 5810
rect 4245 5750 4255 5810
rect 4175 5700 4255 5750
rect 4175 5640 4185 5700
rect 4245 5640 4255 5700
rect 4175 5635 4255 5640
rect 4575 5810 4655 5815
rect 4575 5750 4585 5810
rect 4645 5750 4655 5810
rect 4575 5700 4655 5750
rect 4575 5640 4585 5700
rect 4645 5640 4655 5700
rect 4575 5635 4655 5640
rect 4975 5810 5055 5815
rect 4975 5750 4985 5810
rect 5045 5750 5055 5810
rect 4975 5700 5055 5750
rect 4975 5640 4985 5700
rect 5045 5640 5055 5700
rect 4975 5635 5055 5640
rect 5375 5810 5455 5815
rect 5375 5750 5385 5810
rect 5445 5750 5455 5810
rect 5375 5700 5455 5750
rect 5375 5640 5385 5700
rect 5445 5640 5455 5700
rect 5375 5635 5455 5640
rect 5775 5810 5855 5815
rect 5775 5750 5785 5810
rect 5845 5750 5855 5810
rect 5775 5700 5855 5750
rect 5775 5640 5785 5700
rect 5845 5640 5855 5700
rect 5775 5635 5855 5640
rect 6175 5810 6255 5815
rect 6175 5750 6185 5810
rect 6245 5750 6255 5810
rect 6175 5700 6255 5750
rect 6175 5640 6185 5700
rect 6245 5640 6255 5700
rect 6175 5635 6255 5640
rect 6575 5810 6655 5815
rect 6575 5750 6585 5810
rect 6645 5750 6655 5810
rect 6575 5700 6655 5750
rect 6575 5640 6585 5700
rect 6645 5640 6655 5700
rect 6575 5635 6655 5640
rect 6975 5810 7055 5815
rect 6975 5750 6985 5810
rect 7045 5750 7055 5810
rect 6975 5700 7055 5750
rect 6975 5640 6985 5700
rect 7045 5640 7055 5700
rect 6975 5635 7055 5640
rect 7375 5810 7455 5815
rect 7375 5750 7385 5810
rect 7445 5750 7455 5810
rect 7375 5700 7455 5750
rect 7375 5640 7385 5700
rect 7445 5640 7455 5700
rect 7375 5635 7455 5640
rect 7775 5810 7855 5815
rect 7775 5750 7785 5810
rect 7845 5750 7855 5810
rect 7775 5700 7855 5750
rect 7775 5640 7785 5700
rect 7845 5640 7855 5700
rect 7775 5635 7855 5640
rect 8175 5810 8255 5815
rect 8175 5750 8185 5810
rect 8245 5750 8255 5810
rect 8175 5700 8255 5750
rect 8175 5640 8185 5700
rect 8245 5640 8255 5700
rect 8175 5635 8255 5640
rect 8575 5810 8655 5815
rect 8575 5750 8585 5810
rect 8645 5750 8655 5810
rect 8575 5700 8655 5750
rect 8575 5640 8585 5700
rect 8645 5640 8655 5700
rect 8575 5635 8655 5640
rect 8975 5810 9055 5815
rect 8975 5750 8985 5810
rect 9045 5750 9055 5810
rect 8975 5700 9055 5750
rect 8975 5640 8985 5700
rect 9045 5640 9055 5700
rect 8975 5635 9055 5640
rect 9375 5810 9455 5815
rect 9375 5750 9385 5810
rect 9445 5750 9455 5810
rect 9375 5700 9455 5750
rect 9375 5640 9385 5700
rect 9445 5640 9455 5700
rect 9375 5635 9455 5640
rect 9775 5810 9855 5815
rect 9775 5750 9785 5810
rect 9845 5750 9855 5810
rect 9775 5700 9855 5750
rect 9775 5640 9785 5700
rect 9845 5640 9855 5700
rect 9775 5635 9855 5640
rect 10175 5810 10255 5815
rect 10175 5750 10185 5810
rect 10245 5750 10255 5810
rect 10175 5700 10255 5750
rect 10175 5640 10185 5700
rect 10245 5640 10255 5700
rect 10175 5635 10255 5640
rect 10575 5810 10655 5815
rect 10575 5750 10585 5810
rect 10645 5750 10655 5810
rect 10575 5700 10655 5750
rect 10575 5640 10585 5700
rect 10645 5640 10655 5700
rect 10575 5635 10655 5640
rect 10975 5810 11055 5815
rect 10975 5750 10985 5810
rect 11045 5750 11055 5810
rect 10975 5700 11055 5750
rect 10975 5640 10985 5700
rect 11045 5640 11055 5700
rect 10975 5635 11055 5640
rect 11375 5810 11455 5815
rect 11375 5750 11385 5810
rect 11445 5750 11455 5810
rect 11375 5700 11455 5750
rect 11375 5640 11385 5700
rect 11445 5640 11455 5700
rect 11375 5635 11455 5640
rect 11775 5810 11855 5815
rect 11775 5750 11785 5810
rect 11845 5750 11855 5810
rect 11775 5700 11855 5750
rect 11775 5640 11785 5700
rect 11845 5640 11855 5700
rect 11775 5635 11855 5640
rect 12175 5810 12255 5815
rect 12175 5750 12185 5810
rect 12245 5750 12255 5810
rect 12175 5700 12255 5750
rect 12175 5640 12185 5700
rect 12245 5640 12255 5700
rect 12175 5635 12255 5640
rect 12575 5810 12655 5815
rect 12575 5750 12585 5810
rect 12645 5750 12655 5810
rect 12575 5700 12655 5750
rect 12575 5640 12585 5700
rect 12645 5640 12655 5700
rect 12575 5635 12655 5640
rect 12975 5810 13055 5815
rect 12975 5750 12985 5810
rect 13045 5750 13055 5810
rect 12975 5700 13055 5750
rect 12975 5640 12985 5700
rect 13045 5640 13055 5700
rect 12975 5635 13055 5640
rect -215 5445 -155 5635
rect 185 5445 245 5635
rect 585 5445 645 5635
rect 985 5445 1045 5635
rect 1385 5445 1445 5635
rect 1785 5445 1845 5635
rect 2185 5445 2245 5635
rect 2585 5445 2645 5635
rect 2985 5445 3045 5635
rect 3385 5445 3445 5635
rect 3785 5445 3845 5635
rect 4185 5445 4245 5635
rect 4585 5445 4645 5635
rect 4985 5445 5045 5635
rect 5385 5445 5445 5635
rect 5785 5445 5845 5635
rect 6185 5445 6245 5635
rect 6585 5445 6645 5635
rect 6985 5445 7045 5635
rect 7385 5445 7445 5635
rect 7785 5445 7845 5635
rect 8185 5445 8245 5635
rect 8585 5445 8645 5635
rect 8985 5445 9045 5635
rect 9385 5445 9445 5635
rect 9785 5445 9845 5635
rect 10185 5445 10245 5635
rect 10585 5445 10645 5635
rect 10985 5445 11045 5635
rect 11385 5445 11445 5635
rect 11785 5445 11845 5635
rect 12185 5445 12245 5635
rect 12585 5445 12645 5635
rect 12985 5445 13045 5635
rect -225 5440 -145 5445
rect -225 5380 -215 5440
rect -155 5380 -145 5440
rect -225 5330 -145 5380
rect -225 5270 -215 5330
rect -155 5270 -145 5330
rect -225 5265 -145 5270
rect 175 5440 255 5445
rect 175 5380 185 5440
rect 245 5380 255 5440
rect 175 5330 255 5380
rect 175 5270 185 5330
rect 245 5270 255 5330
rect 175 5265 255 5270
rect 575 5440 655 5445
rect 575 5380 585 5440
rect 645 5380 655 5440
rect 575 5330 655 5380
rect 575 5270 585 5330
rect 645 5270 655 5330
rect 575 5265 655 5270
rect 975 5440 1055 5445
rect 975 5380 985 5440
rect 1045 5380 1055 5440
rect 975 5330 1055 5380
rect 975 5270 985 5330
rect 1045 5270 1055 5330
rect 975 5265 1055 5270
rect 1375 5440 1455 5445
rect 1375 5380 1385 5440
rect 1445 5380 1455 5440
rect 1375 5330 1455 5380
rect 1375 5270 1385 5330
rect 1445 5270 1455 5330
rect 1375 5265 1455 5270
rect 1775 5440 1855 5445
rect 1775 5380 1785 5440
rect 1845 5380 1855 5440
rect 1775 5330 1855 5380
rect 1775 5270 1785 5330
rect 1845 5270 1855 5330
rect 1775 5265 1855 5270
rect 2175 5440 2255 5445
rect 2175 5380 2185 5440
rect 2245 5380 2255 5440
rect 2175 5330 2255 5380
rect 2175 5270 2185 5330
rect 2245 5270 2255 5330
rect 2175 5265 2255 5270
rect 2575 5440 2655 5445
rect 2575 5380 2585 5440
rect 2645 5380 2655 5440
rect 2575 5330 2655 5380
rect 2575 5270 2585 5330
rect 2645 5270 2655 5330
rect 2575 5265 2655 5270
rect 2975 5440 3055 5445
rect 2975 5380 2985 5440
rect 3045 5380 3055 5440
rect 2975 5330 3055 5380
rect 2975 5270 2985 5330
rect 3045 5270 3055 5330
rect 2975 5265 3055 5270
rect 3375 5440 3455 5445
rect 3375 5380 3385 5440
rect 3445 5380 3455 5440
rect 3375 5330 3455 5380
rect 3375 5270 3385 5330
rect 3445 5270 3455 5330
rect 3375 5265 3455 5270
rect 3775 5440 3855 5445
rect 3775 5380 3785 5440
rect 3845 5380 3855 5440
rect 3775 5330 3855 5380
rect 3775 5270 3785 5330
rect 3845 5270 3855 5330
rect 3775 5265 3855 5270
rect 4175 5440 4255 5445
rect 4175 5380 4185 5440
rect 4245 5380 4255 5440
rect 4175 5330 4255 5380
rect 4175 5270 4185 5330
rect 4245 5270 4255 5330
rect 4175 5265 4255 5270
rect 4575 5440 4655 5445
rect 4575 5380 4585 5440
rect 4645 5380 4655 5440
rect 4575 5330 4655 5380
rect 4575 5270 4585 5330
rect 4645 5270 4655 5330
rect 4575 5265 4655 5270
rect 4975 5440 5055 5445
rect 4975 5380 4985 5440
rect 5045 5380 5055 5440
rect 4975 5330 5055 5380
rect 4975 5270 4985 5330
rect 5045 5270 5055 5330
rect 4975 5265 5055 5270
rect 5375 5440 5455 5445
rect 5375 5380 5385 5440
rect 5445 5380 5455 5440
rect 5375 5330 5455 5380
rect 5375 5270 5385 5330
rect 5445 5270 5455 5330
rect 5375 5265 5455 5270
rect 5775 5440 5855 5445
rect 5775 5380 5785 5440
rect 5845 5380 5855 5440
rect 5775 5330 5855 5380
rect 5775 5270 5785 5330
rect 5845 5270 5855 5330
rect 5775 5265 5855 5270
rect 6175 5440 6255 5445
rect 6175 5380 6185 5440
rect 6245 5380 6255 5440
rect 6175 5330 6255 5380
rect 6175 5270 6185 5330
rect 6245 5270 6255 5330
rect 6175 5265 6255 5270
rect 6575 5440 6655 5445
rect 6575 5380 6585 5440
rect 6645 5380 6655 5440
rect 6575 5330 6655 5380
rect 6575 5270 6585 5330
rect 6645 5270 6655 5330
rect 6575 5265 6655 5270
rect 6975 5440 7055 5445
rect 6975 5380 6985 5440
rect 7045 5380 7055 5440
rect 6975 5330 7055 5380
rect 6975 5270 6985 5330
rect 7045 5270 7055 5330
rect 6975 5265 7055 5270
rect 7375 5440 7455 5445
rect 7375 5380 7385 5440
rect 7445 5380 7455 5440
rect 7375 5330 7455 5380
rect 7375 5270 7385 5330
rect 7445 5270 7455 5330
rect 7375 5265 7455 5270
rect 7775 5440 7855 5445
rect 7775 5380 7785 5440
rect 7845 5380 7855 5440
rect 7775 5330 7855 5380
rect 7775 5270 7785 5330
rect 7845 5270 7855 5330
rect 7775 5265 7855 5270
rect 8175 5440 8255 5445
rect 8175 5380 8185 5440
rect 8245 5380 8255 5440
rect 8175 5330 8255 5380
rect 8175 5270 8185 5330
rect 8245 5270 8255 5330
rect 8175 5265 8255 5270
rect 8575 5440 8655 5445
rect 8575 5380 8585 5440
rect 8645 5380 8655 5440
rect 8575 5330 8655 5380
rect 8575 5270 8585 5330
rect 8645 5270 8655 5330
rect 8575 5265 8655 5270
rect 8975 5440 9055 5445
rect 8975 5380 8985 5440
rect 9045 5380 9055 5440
rect 8975 5330 9055 5380
rect 8975 5270 8985 5330
rect 9045 5270 9055 5330
rect 8975 5265 9055 5270
rect 9375 5440 9455 5445
rect 9375 5380 9385 5440
rect 9445 5380 9455 5440
rect 9375 5330 9455 5380
rect 9375 5270 9385 5330
rect 9445 5270 9455 5330
rect 9375 5265 9455 5270
rect 9775 5440 9855 5445
rect 9775 5380 9785 5440
rect 9845 5380 9855 5440
rect 9775 5330 9855 5380
rect 9775 5270 9785 5330
rect 9845 5270 9855 5330
rect 9775 5265 9855 5270
rect 10175 5440 10255 5445
rect 10175 5380 10185 5440
rect 10245 5380 10255 5440
rect 10175 5330 10255 5380
rect 10175 5270 10185 5330
rect 10245 5270 10255 5330
rect 10175 5265 10255 5270
rect 10575 5440 10655 5445
rect 10575 5380 10585 5440
rect 10645 5380 10655 5440
rect 10575 5330 10655 5380
rect 10575 5270 10585 5330
rect 10645 5270 10655 5330
rect 10575 5265 10655 5270
rect 10975 5440 11055 5445
rect 10975 5380 10985 5440
rect 11045 5380 11055 5440
rect 10975 5330 11055 5380
rect 10975 5270 10985 5330
rect 11045 5270 11055 5330
rect 10975 5265 11055 5270
rect 11375 5440 11455 5445
rect 11375 5380 11385 5440
rect 11445 5380 11455 5440
rect 11375 5330 11455 5380
rect 11375 5270 11385 5330
rect 11445 5270 11455 5330
rect 11375 5265 11455 5270
rect 11775 5440 11855 5445
rect 11775 5380 11785 5440
rect 11845 5380 11855 5440
rect 11775 5330 11855 5380
rect 11775 5270 11785 5330
rect 11845 5270 11855 5330
rect 11775 5265 11855 5270
rect 12175 5440 12255 5445
rect 12175 5380 12185 5440
rect 12245 5380 12255 5440
rect 12175 5330 12255 5380
rect 12175 5270 12185 5330
rect 12245 5270 12255 5330
rect 12175 5265 12255 5270
rect 12575 5440 12655 5445
rect 12575 5380 12585 5440
rect 12645 5380 12655 5440
rect 12575 5330 12655 5380
rect 12575 5270 12585 5330
rect 12645 5270 12655 5330
rect 12575 5265 12655 5270
rect 12975 5440 13055 5445
rect 12975 5380 12985 5440
rect 13045 5380 13055 5440
rect 12975 5330 13055 5380
rect 12975 5270 12985 5330
rect 13045 5270 13055 5330
rect 12975 5265 13055 5270
rect -215 5075 -155 5265
rect 185 5075 245 5265
rect 585 5075 645 5265
rect 985 5075 1045 5265
rect 1385 5075 1445 5265
rect 1785 5075 1845 5265
rect 2185 5075 2245 5265
rect 2585 5075 2645 5265
rect 2985 5075 3045 5265
rect 3385 5075 3445 5265
rect 3785 5075 3845 5265
rect 4185 5075 4245 5265
rect 4585 5075 4645 5265
rect 4985 5075 5045 5265
rect 5385 5075 5445 5265
rect 5785 5075 5845 5265
rect 6185 5075 6245 5265
rect 6585 5075 6645 5265
rect 6985 5075 7045 5265
rect 7385 5075 7445 5265
rect 7785 5075 7845 5265
rect 8185 5075 8245 5265
rect 8585 5075 8645 5265
rect 8985 5075 9045 5265
rect 9385 5075 9445 5265
rect 9785 5075 9845 5265
rect 10185 5075 10245 5265
rect 10585 5075 10645 5265
rect 10985 5075 11045 5265
rect 11385 5075 11445 5265
rect 11785 5075 11845 5265
rect 12185 5075 12245 5265
rect 12585 5075 12645 5265
rect 12985 5075 13045 5265
rect -225 5070 -145 5075
rect -225 5010 -215 5070
rect -155 5010 -145 5070
rect -225 4960 -145 5010
rect -225 4900 -215 4960
rect -155 4900 -145 4960
rect -225 4895 -145 4900
rect 175 5070 255 5075
rect 175 5010 185 5070
rect 245 5010 255 5070
rect 175 4960 255 5010
rect 175 4900 185 4960
rect 245 4900 255 4960
rect 175 4895 255 4900
rect 575 5070 655 5075
rect 575 5010 585 5070
rect 645 5010 655 5070
rect 575 4960 655 5010
rect 575 4900 585 4960
rect 645 4900 655 4960
rect 575 4895 655 4900
rect 975 5070 1055 5075
rect 975 5010 985 5070
rect 1045 5010 1055 5070
rect 975 4960 1055 5010
rect 975 4900 985 4960
rect 1045 4900 1055 4960
rect 975 4895 1055 4900
rect 1375 5070 1455 5075
rect 1375 5010 1385 5070
rect 1445 5010 1455 5070
rect 1375 4960 1455 5010
rect 1375 4900 1385 4960
rect 1445 4900 1455 4960
rect 1375 4895 1455 4900
rect 1775 5070 1855 5075
rect 1775 5010 1785 5070
rect 1845 5010 1855 5070
rect 1775 4960 1855 5010
rect 1775 4900 1785 4960
rect 1845 4900 1855 4960
rect 1775 4895 1855 4900
rect 2175 5070 2255 5075
rect 2175 5010 2185 5070
rect 2245 5010 2255 5070
rect 2175 4960 2255 5010
rect 2175 4900 2185 4960
rect 2245 4900 2255 4960
rect 2175 4895 2255 4900
rect 2575 5070 2655 5075
rect 2575 5010 2585 5070
rect 2645 5010 2655 5070
rect 2575 4960 2655 5010
rect 2575 4900 2585 4960
rect 2645 4900 2655 4960
rect 2575 4895 2655 4900
rect 2975 5070 3055 5075
rect 2975 5010 2985 5070
rect 3045 5010 3055 5070
rect 2975 4960 3055 5010
rect 2975 4900 2985 4960
rect 3045 4900 3055 4960
rect 2975 4895 3055 4900
rect 3375 5070 3455 5075
rect 3375 5010 3385 5070
rect 3445 5010 3455 5070
rect 3375 4960 3455 5010
rect 3375 4900 3385 4960
rect 3445 4900 3455 4960
rect 3375 4895 3455 4900
rect 3775 5070 3855 5075
rect 3775 5010 3785 5070
rect 3845 5010 3855 5070
rect 3775 4960 3855 5010
rect 3775 4900 3785 4960
rect 3845 4900 3855 4960
rect 3775 4895 3855 4900
rect 4175 5070 4255 5075
rect 4175 5010 4185 5070
rect 4245 5010 4255 5070
rect 4175 4960 4255 5010
rect 4175 4900 4185 4960
rect 4245 4900 4255 4960
rect 4175 4895 4255 4900
rect 4575 5070 4655 5075
rect 4575 5010 4585 5070
rect 4645 5010 4655 5070
rect 4575 4960 4655 5010
rect 4575 4900 4585 4960
rect 4645 4900 4655 4960
rect 4575 4895 4655 4900
rect 4975 5070 5055 5075
rect 4975 5010 4985 5070
rect 5045 5010 5055 5070
rect 4975 4960 5055 5010
rect 4975 4900 4985 4960
rect 5045 4900 5055 4960
rect 4975 4895 5055 4900
rect 5375 5070 5455 5075
rect 5375 5010 5385 5070
rect 5445 5010 5455 5070
rect 5375 4960 5455 5010
rect 5375 4900 5385 4960
rect 5445 4900 5455 4960
rect 5375 4895 5455 4900
rect 5775 5070 5855 5075
rect 5775 5010 5785 5070
rect 5845 5010 5855 5070
rect 5775 4960 5855 5010
rect 5775 4900 5785 4960
rect 5845 4900 5855 4960
rect 5775 4895 5855 4900
rect 6175 5070 6255 5075
rect 6175 5010 6185 5070
rect 6245 5010 6255 5070
rect 6175 4960 6255 5010
rect 6175 4900 6185 4960
rect 6245 4900 6255 4960
rect 6175 4895 6255 4900
rect 6575 5070 6655 5075
rect 6575 5010 6585 5070
rect 6645 5010 6655 5070
rect 6575 4960 6655 5010
rect 6575 4900 6585 4960
rect 6645 4900 6655 4960
rect 6575 4895 6655 4900
rect 6975 5070 7055 5075
rect 6975 5010 6985 5070
rect 7045 5010 7055 5070
rect 6975 4960 7055 5010
rect 6975 4900 6985 4960
rect 7045 4900 7055 4960
rect 6975 4895 7055 4900
rect 7375 5070 7455 5075
rect 7375 5010 7385 5070
rect 7445 5010 7455 5070
rect 7375 4960 7455 5010
rect 7375 4900 7385 4960
rect 7445 4900 7455 4960
rect 7375 4895 7455 4900
rect 7775 5070 7855 5075
rect 7775 5010 7785 5070
rect 7845 5010 7855 5070
rect 7775 4960 7855 5010
rect 7775 4900 7785 4960
rect 7845 4900 7855 4960
rect 7775 4895 7855 4900
rect 8175 5070 8255 5075
rect 8175 5010 8185 5070
rect 8245 5010 8255 5070
rect 8175 4960 8255 5010
rect 8175 4900 8185 4960
rect 8245 4900 8255 4960
rect 8175 4895 8255 4900
rect 8575 5070 8655 5075
rect 8575 5010 8585 5070
rect 8645 5010 8655 5070
rect 8575 4960 8655 5010
rect 8575 4900 8585 4960
rect 8645 4900 8655 4960
rect 8575 4895 8655 4900
rect 8975 5070 9055 5075
rect 8975 5010 8985 5070
rect 9045 5010 9055 5070
rect 8975 4960 9055 5010
rect 8975 4900 8985 4960
rect 9045 4900 9055 4960
rect 8975 4895 9055 4900
rect 9375 5070 9455 5075
rect 9375 5010 9385 5070
rect 9445 5010 9455 5070
rect 9375 4960 9455 5010
rect 9375 4900 9385 4960
rect 9445 4900 9455 4960
rect 9375 4895 9455 4900
rect 9775 5070 9855 5075
rect 9775 5010 9785 5070
rect 9845 5010 9855 5070
rect 9775 4960 9855 5010
rect 9775 4900 9785 4960
rect 9845 4900 9855 4960
rect 9775 4895 9855 4900
rect 10175 5070 10255 5075
rect 10175 5010 10185 5070
rect 10245 5010 10255 5070
rect 10175 4960 10255 5010
rect 10175 4900 10185 4960
rect 10245 4900 10255 4960
rect 10175 4895 10255 4900
rect 10575 5070 10655 5075
rect 10575 5010 10585 5070
rect 10645 5010 10655 5070
rect 10575 4960 10655 5010
rect 10575 4900 10585 4960
rect 10645 4900 10655 4960
rect 10575 4895 10655 4900
rect 10975 5070 11055 5075
rect 10975 5010 10985 5070
rect 11045 5010 11055 5070
rect 10975 4960 11055 5010
rect 10975 4900 10985 4960
rect 11045 4900 11055 4960
rect 10975 4895 11055 4900
rect 11375 5070 11455 5075
rect 11375 5010 11385 5070
rect 11445 5010 11455 5070
rect 11375 4960 11455 5010
rect 11375 4900 11385 4960
rect 11445 4900 11455 4960
rect 11375 4895 11455 4900
rect 11775 5070 11855 5075
rect 11775 5010 11785 5070
rect 11845 5010 11855 5070
rect 11775 4960 11855 5010
rect 11775 4900 11785 4960
rect 11845 4900 11855 4960
rect 11775 4895 11855 4900
rect 12175 5070 12255 5075
rect 12175 5010 12185 5070
rect 12245 5010 12255 5070
rect 12175 4960 12255 5010
rect 12175 4900 12185 4960
rect 12245 4900 12255 4960
rect 12175 4895 12255 4900
rect 12575 5070 12655 5075
rect 12575 5010 12585 5070
rect 12645 5010 12655 5070
rect 12575 4960 12655 5010
rect 12575 4900 12585 4960
rect 12645 4900 12655 4960
rect 12575 4895 12655 4900
rect 12975 5070 13055 5075
rect 12975 5010 12985 5070
rect 13045 5010 13055 5070
rect 12975 4960 13055 5010
rect 12975 4900 12985 4960
rect 13045 4900 13055 4960
rect 12975 4895 13055 4900
rect -215 4705 -155 4895
rect 185 4705 245 4895
rect 585 4705 645 4895
rect 985 4705 1045 4895
rect 1385 4705 1445 4895
rect 1785 4705 1845 4895
rect 2185 4705 2245 4895
rect 2585 4705 2645 4895
rect 2985 4705 3045 4895
rect 3385 4705 3445 4895
rect 3785 4705 3845 4895
rect 4185 4705 4245 4895
rect 4585 4705 4645 4895
rect 4985 4705 5045 4895
rect 5385 4705 5445 4895
rect 5785 4705 5845 4895
rect 6185 4705 6245 4895
rect 6585 4705 6645 4895
rect 6985 4705 7045 4895
rect 7385 4705 7445 4895
rect 7785 4705 7845 4895
rect 8185 4705 8245 4895
rect 8585 4705 8645 4895
rect 8985 4705 9045 4895
rect 9385 4705 9445 4895
rect 9785 4705 9845 4895
rect 10185 4705 10245 4895
rect 10585 4705 10645 4895
rect 10985 4705 11045 4895
rect 11385 4705 11445 4895
rect 11785 4705 11845 4895
rect 12185 4705 12245 4895
rect 12585 4705 12645 4895
rect 12985 4705 13045 4895
rect -225 4700 -145 4705
rect -225 4640 -215 4700
rect -155 4640 -145 4700
rect -225 4590 -145 4640
rect -225 4530 -215 4590
rect -155 4530 -145 4590
rect -225 4525 -145 4530
rect 175 4700 255 4705
rect 175 4640 185 4700
rect 245 4640 255 4700
rect 175 4590 255 4640
rect 175 4530 185 4590
rect 245 4530 255 4590
rect 175 4525 255 4530
rect 575 4700 655 4705
rect 575 4640 585 4700
rect 645 4640 655 4700
rect 575 4590 655 4640
rect 575 4530 585 4590
rect 645 4530 655 4590
rect 575 4525 655 4530
rect 975 4700 1055 4705
rect 975 4640 985 4700
rect 1045 4640 1055 4700
rect 975 4590 1055 4640
rect 975 4530 985 4590
rect 1045 4530 1055 4590
rect 975 4525 1055 4530
rect 1375 4700 1455 4705
rect 1375 4640 1385 4700
rect 1445 4640 1455 4700
rect 1375 4590 1455 4640
rect 1375 4530 1385 4590
rect 1445 4530 1455 4590
rect 1375 4525 1455 4530
rect 1775 4700 1855 4705
rect 1775 4640 1785 4700
rect 1845 4640 1855 4700
rect 1775 4590 1855 4640
rect 1775 4530 1785 4590
rect 1845 4530 1855 4590
rect 1775 4525 1855 4530
rect 2175 4700 2255 4705
rect 2175 4640 2185 4700
rect 2245 4640 2255 4700
rect 2175 4590 2255 4640
rect 2175 4530 2185 4590
rect 2245 4530 2255 4590
rect 2175 4525 2255 4530
rect 2575 4700 2655 4705
rect 2575 4640 2585 4700
rect 2645 4640 2655 4700
rect 2575 4590 2655 4640
rect 2575 4530 2585 4590
rect 2645 4530 2655 4590
rect 2575 4525 2655 4530
rect 2975 4700 3055 4705
rect 2975 4640 2985 4700
rect 3045 4640 3055 4700
rect 2975 4590 3055 4640
rect 2975 4530 2985 4590
rect 3045 4530 3055 4590
rect 2975 4525 3055 4530
rect 3375 4700 3455 4705
rect 3375 4640 3385 4700
rect 3445 4640 3455 4700
rect 3375 4590 3455 4640
rect 3375 4530 3385 4590
rect 3445 4530 3455 4590
rect 3375 4525 3455 4530
rect 3775 4700 3855 4705
rect 3775 4640 3785 4700
rect 3845 4640 3855 4700
rect 3775 4590 3855 4640
rect 3775 4530 3785 4590
rect 3845 4530 3855 4590
rect 3775 4525 3855 4530
rect 4175 4700 4255 4705
rect 4175 4640 4185 4700
rect 4245 4640 4255 4700
rect 4175 4590 4255 4640
rect 4175 4530 4185 4590
rect 4245 4530 4255 4590
rect 4175 4525 4255 4530
rect 4575 4700 4655 4705
rect 4575 4640 4585 4700
rect 4645 4640 4655 4700
rect 4575 4590 4655 4640
rect 4575 4530 4585 4590
rect 4645 4530 4655 4590
rect 4575 4525 4655 4530
rect 4975 4700 5055 4705
rect 4975 4640 4985 4700
rect 5045 4640 5055 4700
rect 4975 4590 5055 4640
rect 4975 4530 4985 4590
rect 5045 4530 5055 4590
rect 4975 4525 5055 4530
rect 5375 4700 5455 4705
rect 5375 4640 5385 4700
rect 5445 4640 5455 4700
rect 5375 4590 5455 4640
rect 5375 4530 5385 4590
rect 5445 4530 5455 4590
rect 5375 4525 5455 4530
rect 5775 4700 5855 4705
rect 5775 4640 5785 4700
rect 5845 4640 5855 4700
rect 5775 4590 5855 4640
rect 5775 4530 5785 4590
rect 5845 4530 5855 4590
rect 5775 4525 5855 4530
rect 6175 4700 6255 4705
rect 6175 4640 6185 4700
rect 6245 4640 6255 4700
rect 6175 4590 6255 4640
rect 6175 4530 6185 4590
rect 6245 4530 6255 4590
rect 6175 4525 6255 4530
rect 6575 4700 6655 4705
rect 6575 4640 6585 4700
rect 6645 4640 6655 4700
rect 6575 4590 6655 4640
rect 6575 4530 6585 4590
rect 6645 4530 6655 4590
rect 6575 4525 6655 4530
rect 6975 4700 7055 4705
rect 6975 4640 6985 4700
rect 7045 4640 7055 4700
rect 6975 4590 7055 4640
rect 6975 4530 6985 4590
rect 7045 4530 7055 4590
rect 6975 4525 7055 4530
rect 7375 4700 7455 4705
rect 7375 4640 7385 4700
rect 7445 4640 7455 4700
rect 7375 4590 7455 4640
rect 7375 4530 7385 4590
rect 7445 4530 7455 4590
rect 7375 4525 7455 4530
rect 7775 4700 7855 4705
rect 7775 4640 7785 4700
rect 7845 4640 7855 4700
rect 7775 4590 7855 4640
rect 7775 4530 7785 4590
rect 7845 4530 7855 4590
rect 7775 4525 7855 4530
rect 8175 4700 8255 4705
rect 8175 4640 8185 4700
rect 8245 4640 8255 4700
rect 8175 4590 8255 4640
rect 8175 4530 8185 4590
rect 8245 4530 8255 4590
rect 8175 4525 8255 4530
rect 8575 4700 8655 4705
rect 8575 4640 8585 4700
rect 8645 4640 8655 4700
rect 8575 4590 8655 4640
rect 8575 4530 8585 4590
rect 8645 4530 8655 4590
rect 8575 4525 8655 4530
rect 8975 4700 9055 4705
rect 8975 4640 8985 4700
rect 9045 4640 9055 4700
rect 8975 4590 9055 4640
rect 8975 4530 8985 4590
rect 9045 4530 9055 4590
rect 8975 4525 9055 4530
rect 9375 4700 9455 4705
rect 9375 4640 9385 4700
rect 9445 4640 9455 4700
rect 9375 4590 9455 4640
rect 9375 4530 9385 4590
rect 9445 4530 9455 4590
rect 9375 4525 9455 4530
rect 9775 4700 9855 4705
rect 9775 4640 9785 4700
rect 9845 4640 9855 4700
rect 9775 4590 9855 4640
rect 9775 4530 9785 4590
rect 9845 4530 9855 4590
rect 9775 4525 9855 4530
rect 10175 4700 10255 4705
rect 10175 4640 10185 4700
rect 10245 4640 10255 4700
rect 10175 4590 10255 4640
rect 10175 4530 10185 4590
rect 10245 4530 10255 4590
rect 10175 4525 10255 4530
rect 10575 4700 10655 4705
rect 10575 4640 10585 4700
rect 10645 4640 10655 4700
rect 10575 4590 10655 4640
rect 10575 4530 10585 4590
rect 10645 4530 10655 4590
rect 10575 4525 10655 4530
rect 10975 4700 11055 4705
rect 10975 4640 10985 4700
rect 11045 4640 11055 4700
rect 10975 4590 11055 4640
rect 10975 4530 10985 4590
rect 11045 4530 11055 4590
rect 10975 4525 11055 4530
rect 11375 4700 11455 4705
rect 11375 4640 11385 4700
rect 11445 4640 11455 4700
rect 11375 4590 11455 4640
rect 11375 4530 11385 4590
rect 11445 4530 11455 4590
rect 11375 4525 11455 4530
rect 11775 4700 11855 4705
rect 11775 4640 11785 4700
rect 11845 4640 11855 4700
rect 11775 4590 11855 4640
rect 11775 4530 11785 4590
rect 11845 4530 11855 4590
rect 11775 4525 11855 4530
rect 12175 4700 12255 4705
rect 12175 4640 12185 4700
rect 12245 4640 12255 4700
rect 12175 4590 12255 4640
rect 12175 4530 12185 4590
rect 12245 4530 12255 4590
rect 12175 4525 12255 4530
rect 12575 4700 12655 4705
rect 12575 4640 12585 4700
rect 12645 4640 12655 4700
rect 12575 4590 12655 4640
rect 12575 4530 12585 4590
rect 12645 4530 12655 4590
rect 12575 4525 12655 4530
rect 12975 4700 13055 4705
rect 12975 4640 12985 4700
rect 13045 4640 13055 4700
rect 12975 4590 13055 4640
rect 12975 4530 12985 4590
rect 13045 4530 13055 4590
rect 12975 4525 13055 4530
rect -215 4335 -155 4525
rect 185 4335 245 4525
rect 585 4335 645 4525
rect 985 4335 1045 4525
rect 1385 4335 1445 4525
rect 1785 4335 1845 4525
rect 2185 4335 2245 4525
rect 2585 4335 2645 4525
rect 2985 4335 3045 4525
rect 3385 4335 3445 4525
rect 3785 4335 3845 4525
rect 4185 4335 4245 4525
rect 4585 4335 4645 4525
rect 4985 4335 5045 4525
rect 5385 4335 5445 4525
rect 5785 4335 5845 4525
rect 6185 4335 6245 4525
rect 6585 4335 6645 4525
rect 6985 4335 7045 4525
rect 7385 4335 7445 4525
rect 7785 4335 7845 4525
rect 8185 4335 8245 4525
rect 8585 4335 8645 4525
rect 8985 4335 9045 4525
rect 9385 4335 9445 4525
rect 9785 4335 9845 4525
rect 10185 4335 10245 4525
rect 10585 4335 10645 4525
rect 10985 4335 11045 4525
rect 11385 4335 11445 4525
rect 11785 4335 11845 4525
rect 12185 4335 12245 4525
rect 12585 4335 12645 4525
rect 12985 4335 13045 4525
rect -225 4330 -145 4335
rect -225 4270 -215 4330
rect -155 4270 -145 4330
rect -225 4220 -145 4270
rect -225 4160 -215 4220
rect -155 4160 -145 4220
rect -225 4155 -145 4160
rect 175 4330 255 4335
rect 175 4270 185 4330
rect 245 4270 255 4330
rect 175 4220 255 4270
rect 175 4160 185 4220
rect 245 4160 255 4220
rect 175 4155 255 4160
rect 575 4330 655 4335
rect 575 4270 585 4330
rect 645 4270 655 4330
rect 575 4220 655 4270
rect 575 4160 585 4220
rect 645 4160 655 4220
rect 575 4155 655 4160
rect 975 4330 1055 4335
rect 975 4270 985 4330
rect 1045 4270 1055 4330
rect 975 4220 1055 4270
rect 975 4160 985 4220
rect 1045 4160 1055 4220
rect 975 4155 1055 4160
rect 1375 4330 1455 4335
rect 1375 4270 1385 4330
rect 1445 4270 1455 4330
rect 1375 4220 1455 4270
rect 1375 4160 1385 4220
rect 1445 4160 1455 4220
rect 1375 4155 1455 4160
rect 1775 4330 1855 4335
rect 1775 4270 1785 4330
rect 1845 4270 1855 4330
rect 1775 4220 1855 4270
rect 1775 4160 1785 4220
rect 1845 4160 1855 4220
rect 1775 4155 1855 4160
rect 2175 4330 2255 4335
rect 2175 4270 2185 4330
rect 2245 4270 2255 4330
rect 2175 4220 2255 4270
rect 2175 4160 2185 4220
rect 2245 4160 2255 4220
rect 2175 4155 2255 4160
rect 2575 4330 2655 4335
rect 2575 4270 2585 4330
rect 2645 4270 2655 4330
rect 2575 4220 2655 4270
rect 2575 4160 2585 4220
rect 2645 4160 2655 4220
rect 2575 4155 2655 4160
rect 2975 4330 3055 4335
rect 2975 4270 2985 4330
rect 3045 4270 3055 4330
rect 2975 4220 3055 4270
rect 2975 4160 2985 4220
rect 3045 4160 3055 4220
rect 2975 4155 3055 4160
rect 3375 4330 3455 4335
rect 3375 4270 3385 4330
rect 3445 4270 3455 4330
rect 3375 4220 3455 4270
rect 3375 4160 3385 4220
rect 3445 4160 3455 4220
rect 3375 4155 3455 4160
rect 3775 4330 3855 4335
rect 3775 4270 3785 4330
rect 3845 4270 3855 4330
rect 3775 4220 3855 4270
rect 3775 4160 3785 4220
rect 3845 4160 3855 4220
rect 3775 4155 3855 4160
rect 4175 4330 4255 4335
rect 4175 4270 4185 4330
rect 4245 4270 4255 4330
rect 4175 4220 4255 4270
rect 4175 4160 4185 4220
rect 4245 4160 4255 4220
rect 4175 4155 4255 4160
rect 4575 4330 4655 4335
rect 4575 4270 4585 4330
rect 4645 4270 4655 4330
rect 4575 4220 4655 4270
rect 4575 4160 4585 4220
rect 4645 4160 4655 4220
rect 4575 4155 4655 4160
rect 4975 4330 5055 4335
rect 4975 4270 4985 4330
rect 5045 4270 5055 4330
rect 4975 4220 5055 4270
rect 4975 4160 4985 4220
rect 5045 4160 5055 4220
rect 4975 4155 5055 4160
rect 5375 4330 5455 4335
rect 5375 4270 5385 4330
rect 5445 4270 5455 4330
rect 5375 4220 5455 4270
rect 5375 4160 5385 4220
rect 5445 4160 5455 4220
rect 5375 4155 5455 4160
rect 5775 4330 5855 4335
rect 5775 4270 5785 4330
rect 5845 4270 5855 4330
rect 5775 4220 5855 4270
rect 5775 4160 5785 4220
rect 5845 4160 5855 4220
rect 5775 4155 5855 4160
rect 6175 4330 6255 4335
rect 6175 4270 6185 4330
rect 6245 4270 6255 4330
rect 6175 4220 6255 4270
rect 6175 4160 6185 4220
rect 6245 4160 6255 4220
rect 6175 4155 6255 4160
rect 6575 4330 6655 4335
rect 6575 4270 6585 4330
rect 6645 4270 6655 4330
rect 6575 4220 6655 4270
rect 6575 4160 6585 4220
rect 6645 4160 6655 4220
rect 6575 4155 6655 4160
rect 6975 4330 7055 4335
rect 6975 4270 6985 4330
rect 7045 4270 7055 4330
rect 6975 4220 7055 4270
rect 6975 4160 6985 4220
rect 7045 4160 7055 4220
rect 6975 4155 7055 4160
rect 7375 4330 7455 4335
rect 7375 4270 7385 4330
rect 7445 4270 7455 4330
rect 7375 4220 7455 4270
rect 7375 4160 7385 4220
rect 7445 4160 7455 4220
rect 7375 4155 7455 4160
rect 7775 4330 7855 4335
rect 7775 4270 7785 4330
rect 7845 4270 7855 4330
rect 7775 4220 7855 4270
rect 7775 4160 7785 4220
rect 7845 4160 7855 4220
rect 7775 4155 7855 4160
rect 8175 4330 8255 4335
rect 8175 4270 8185 4330
rect 8245 4270 8255 4330
rect 8175 4220 8255 4270
rect 8175 4160 8185 4220
rect 8245 4160 8255 4220
rect 8175 4155 8255 4160
rect 8575 4330 8655 4335
rect 8575 4270 8585 4330
rect 8645 4270 8655 4330
rect 8575 4220 8655 4270
rect 8575 4160 8585 4220
rect 8645 4160 8655 4220
rect 8575 4155 8655 4160
rect 8975 4330 9055 4335
rect 8975 4270 8985 4330
rect 9045 4270 9055 4330
rect 8975 4220 9055 4270
rect 8975 4160 8985 4220
rect 9045 4160 9055 4220
rect 8975 4155 9055 4160
rect 9375 4330 9455 4335
rect 9375 4270 9385 4330
rect 9445 4270 9455 4330
rect 9375 4220 9455 4270
rect 9375 4160 9385 4220
rect 9445 4160 9455 4220
rect 9375 4155 9455 4160
rect 9775 4330 9855 4335
rect 9775 4270 9785 4330
rect 9845 4270 9855 4330
rect 9775 4220 9855 4270
rect 9775 4160 9785 4220
rect 9845 4160 9855 4220
rect 9775 4155 9855 4160
rect 10175 4330 10255 4335
rect 10175 4270 10185 4330
rect 10245 4270 10255 4330
rect 10175 4220 10255 4270
rect 10175 4160 10185 4220
rect 10245 4160 10255 4220
rect 10175 4155 10255 4160
rect 10575 4330 10655 4335
rect 10575 4270 10585 4330
rect 10645 4270 10655 4330
rect 10575 4220 10655 4270
rect 10575 4160 10585 4220
rect 10645 4160 10655 4220
rect 10575 4155 10655 4160
rect 10975 4330 11055 4335
rect 10975 4270 10985 4330
rect 11045 4270 11055 4330
rect 10975 4220 11055 4270
rect 10975 4160 10985 4220
rect 11045 4160 11055 4220
rect 10975 4155 11055 4160
rect 11375 4330 11455 4335
rect 11375 4270 11385 4330
rect 11445 4270 11455 4330
rect 11375 4220 11455 4270
rect 11375 4160 11385 4220
rect 11445 4160 11455 4220
rect 11375 4155 11455 4160
rect 11775 4330 11855 4335
rect 11775 4270 11785 4330
rect 11845 4270 11855 4330
rect 11775 4220 11855 4270
rect 11775 4160 11785 4220
rect 11845 4160 11855 4220
rect 11775 4155 11855 4160
rect 12175 4330 12255 4335
rect 12175 4270 12185 4330
rect 12245 4270 12255 4330
rect 12175 4220 12255 4270
rect 12175 4160 12185 4220
rect 12245 4160 12255 4220
rect 12175 4155 12255 4160
rect 12575 4330 12655 4335
rect 12575 4270 12585 4330
rect 12645 4270 12655 4330
rect 12575 4220 12655 4270
rect 12575 4160 12585 4220
rect 12645 4160 12655 4220
rect 12575 4155 12655 4160
rect 12975 4330 13055 4335
rect 12975 4270 12985 4330
rect 13045 4270 13055 4330
rect 12975 4220 13055 4270
rect 12975 4160 12985 4220
rect 13045 4160 13055 4220
rect 12975 4155 13055 4160
rect -215 3965 -155 4155
rect 185 3965 245 4155
rect 585 3965 645 4155
rect 985 3965 1045 4155
rect 1385 3965 1445 4155
rect 1785 3965 1845 4155
rect 2185 3965 2245 4155
rect 2585 3965 2645 4155
rect 2985 3965 3045 4155
rect 3385 3965 3445 4155
rect 3785 3965 3845 4155
rect 4185 3965 4245 4155
rect 4585 3965 4645 4155
rect 4985 3965 5045 4155
rect 5385 3965 5445 4155
rect 5785 3965 5845 4155
rect 6185 3965 6245 4155
rect 6585 3965 6645 4155
rect 6985 3965 7045 4155
rect 7385 3965 7445 4155
rect 7785 3965 7845 4155
rect 8185 3965 8245 4155
rect 8585 3965 8645 4155
rect 8985 3965 9045 4155
rect 9385 3965 9445 4155
rect 9785 3965 9845 4155
rect 10185 3965 10245 4155
rect 10585 3965 10645 4155
rect 10985 3965 11045 4155
rect 11385 3965 11445 4155
rect 11785 3965 11845 4155
rect 12185 3965 12245 4155
rect 12585 3965 12645 4155
rect 12985 3965 13045 4155
rect -225 3960 -145 3965
rect -225 3900 -215 3960
rect -155 3900 -145 3960
rect -225 3850 -145 3900
rect -225 3790 -215 3850
rect -155 3790 -145 3850
rect -225 3785 -145 3790
rect 175 3960 255 3965
rect 175 3900 185 3960
rect 245 3900 255 3960
rect 175 3850 255 3900
rect 175 3790 185 3850
rect 245 3790 255 3850
rect 175 3785 255 3790
rect 575 3960 655 3965
rect 575 3900 585 3960
rect 645 3900 655 3960
rect 575 3850 655 3900
rect 575 3790 585 3850
rect 645 3790 655 3850
rect 575 3785 655 3790
rect 975 3960 1055 3965
rect 975 3900 985 3960
rect 1045 3900 1055 3960
rect 975 3850 1055 3900
rect 975 3790 985 3850
rect 1045 3790 1055 3850
rect 975 3785 1055 3790
rect 1375 3960 1455 3965
rect 1375 3900 1385 3960
rect 1445 3900 1455 3960
rect 1375 3850 1455 3900
rect 1375 3790 1385 3850
rect 1445 3790 1455 3850
rect 1375 3785 1455 3790
rect 1775 3960 1855 3965
rect 1775 3900 1785 3960
rect 1845 3900 1855 3960
rect 1775 3850 1855 3900
rect 1775 3790 1785 3850
rect 1845 3790 1855 3850
rect 1775 3785 1855 3790
rect 2175 3960 2255 3965
rect 2175 3900 2185 3960
rect 2245 3900 2255 3960
rect 2175 3850 2255 3900
rect 2175 3790 2185 3850
rect 2245 3790 2255 3850
rect 2175 3785 2255 3790
rect 2575 3960 2655 3965
rect 2575 3900 2585 3960
rect 2645 3900 2655 3960
rect 2575 3850 2655 3900
rect 2575 3790 2585 3850
rect 2645 3790 2655 3850
rect 2575 3785 2655 3790
rect 2975 3960 3055 3965
rect 2975 3900 2985 3960
rect 3045 3900 3055 3960
rect 2975 3850 3055 3900
rect 2975 3790 2985 3850
rect 3045 3790 3055 3850
rect 2975 3785 3055 3790
rect 3375 3960 3455 3965
rect 3375 3900 3385 3960
rect 3445 3900 3455 3960
rect 3375 3850 3455 3900
rect 3375 3790 3385 3850
rect 3445 3790 3455 3850
rect 3375 3785 3455 3790
rect 3775 3960 3855 3965
rect 3775 3900 3785 3960
rect 3845 3900 3855 3960
rect 3775 3850 3855 3900
rect 3775 3790 3785 3850
rect 3845 3790 3855 3850
rect 3775 3785 3855 3790
rect 4175 3960 4255 3965
rect 4175 3900 4185 3960
rect 4245 3900 4255 3960
rect 4175 3850 4255 3900
rect 4175 3790 4185 3850
rect 4245 3790 4255 3850
rect 4175 3785 4255 3790
rect 4575 3960 4655 3965
rect 4575 3900 4585 3960
rect 4645 3900 4655 3960
rect 4575 3850 4655 3900
rect 4575 3790 4585 3850
rect 4645 3790 4655 3850
rect 4575 3785 4655 3790
rect 4975 3960 5055 3965
rect 4975 3900 4985 3960
rect 5045 3900 5055 3960
rect 4975 3850 5055 3900
rect 4975 3790 4985 3850
rect 5045 3790 5055 3850
rect 4975 3785 5055 3790
rect 5375 3960 5455 3965
rect 5375 3900 5385 3960
rect 5445 3900 5455 3960
rect 5375 3850 5455 3900
rect 5375 3790 5385 3850
rect 5445 3790 5455 3850
rect 5375 3785 5455 3790
rect 5775 3960 5855 3965
rect 5775 3900 5785 3960
rect 5845 3900 5855 3960
rect 5775 3850 5855 3900
rect 5775 3790 5785 3850
rect 5845 3790 5855 3850
rect 5775 3785 5855 3790
rect 6175 3960 6255 3965
rect 6175 3900 6185 3960
rect 6245 3900 6255 3960
rect 6175 3850 6255 3900
rect 6175 3790 6185 3850
rect 6245 3790 6255 3850
rect 6175 3785 6255 3790
rect 6575 3960 6655 3965
rect 6575 3900 6585 3960
rect 6645 3900 6655 3960
rect 6575 3850 6655 3900
rect 6575 3790 6585 3850
rect 6645 3790 6655 3850
rect 6575 3785 6655 3790
rect 6975 3960 7055 3965
rect 6975 3900 6985 3960
rect 7045 3900 7055 3960
rect 6975 3850 7055 3900
rect 6975 3790 6985 3850
rect 7045 3790 7055 3850
rect 6975 3785 7055 3790
rect 7375 3960 7455 3965
rect 7375 3900 7385 3960
rect 7445 3900 7455 3960
rect 7375 3850 7455 3900
rect 7375 3790 7385 3850
rect 7445 3790 7455 3850
rect 7375 3785 7455 3790
rect 7775 3960 7855 3965
rect 7775 3900 7785 3960
rect 7845 3900 7855 3960
rect 7775 3850 7855 3900
rect 7775 3790 7785 3850
rect 7845 3790 7855 3850
rect 7775 3785 7855 3790
rect 8175 3960 8255 3965
rect 8175 3900 8185 3960
rect 8245 3900 8255 3960
rect 8175 3850 8255 3900
rect 8175 3790 8185 3850
rect 8245 3790 8255 3850
rect 8175 3785 8255 3790
rect 8575 3960 8655 3965
rect 8575 3900 8585 3960
rect 8645 3900 8655 3960
rect 8575 3850 8655 3900
rect 8575 3790 8585 3850
rect 8645 3790 8655 3850
rect 8575 3785 8655 3790
rect 8975 3960 9055 3965
rect 8975 3900 8985 3960
rect 9045 3900 9055 3960
rect 8975 3850 9055 3900
rect 8975 3790 8985 3850
rect 9045 3790 9055 3850
rect 8975 3785 9055 3790
rect 9375 3960 9455 3965
rect 9375 3900 9385 3960
rect 9445 3900 9455 3960
rect 9375 3850 9455 3900
rect 9375 3790 9385 3850
rect 9445 3790 9455 3850
rect 9375 3785 9455 3790
rect 9775 3960 9855 3965
rect 9775 3900 9785 3960
rect 9845 3900 9855 3960
rect 9775 3850 9855 3900
rect 9775 3790 9785 3850
rect 9845 3790 9855 3850
rect 9775 3785 9855 3790
rect 10175 3960 10255 3965
rect 10175 3900 10185 3960
rect 10245 3900 10255 3960
rect 10175 3850 10255 3900
rect 10175 3790 10185 3850
rect 10245 3790 10255 3850
rect 10175 3785 10255 3790
rect 10575 3960 10655 3965
rect 10575 3900 10585 3960
rect 10645 3900 10655 3960
rect 10575 3850 10655 3900
rect 10575 3790 10585 3850
rect 10645 3790 10655 3850
rect 10575 3785 10655 3790
rect 10975 3960 11055 3965
rect 10975 3900 10985 3960
rect 11045 3900 11055 3960
rect 10975 3850 11055 3900
rect 10975 3790 10985 3850
rect 11045 3790 11055 3850
rect 10975 3785 11055 3790
rect 11375 3960 11455 3965
rect 11375 3900 11385 3960
rect 11445 3900 11455 3960
rect 11375 3850 11455 3900
rect 11375 3790 11385 3850
rect 11445 3790 11455 3850
rect 11375 3785 11455 3790
rect 11775 3960 11855 3965
rect 11775 3900 11785 3960
rect 11845 3900 11855 3960
rect 11775 3850 11855 3900
rect 11775 3790 11785 3850
rect 11845 3790 11855 3850
rect 11775 3785 11855 3790
rect 12175 3960 12255 3965
rect 12175 3900 12185 3960
rect 12245 3900 12255 3960
rect 12175 3850 12255 3900
rect 12175 3790 12185 3850
rect 12245 3790 12255 3850
rect 12175 3785 12255 3790
rect 12575 3960 12655 3965
rect 12575 3900 12585 3960
rect 12645 3900 12655 3960
rect 12575 3850 12655 3900
rect 12575 3790 12585 3850
rect 12645 3790 12655 3850
rect 12575 3785 12655 3790
rect 12975 3960 13055 3965
rect 12975 3900 12985 3960
rect 13045 3900 13055 3960
rect 12975 3850 13055 3900
rect 12975 3790 12985 3850
rect 13045 3790 13055 3850
rect 12975 3785 13055 3790
rect -215 3595 -155 3785
rect 185 3595 245 3785
rect 585 3595 645 3785
rect 985 3595 1045 3785
rect 1385 3595 1445 3785
rect 1785 3595 1845 3785
rect 2185 3595 2245 3785
rect 2585 3595 2645 3785
rect 2985 3595 3045 3785
rect 3385 3595 3445 3785
rect 3785 3595 3845 3785
rect 4185 3595 4245 3785
rect 4585 3595 4645 3785
rect 4985 3595 5045 3785
rect 5385 3595 5445 3785
rect 5785 3595 5845 3785
rect 6185 3595 6245 3785
rect 6585 3595 6645 3785
rect 6985 3595 7045 3785
rect 7385 3595 7445 3785
rect 7785 3595 7845 3785
rect 8185 3595 8245 3785
rect 8585 3595 8645 3785
rect 8985 3595 9045 3785
rect 9385 3595 9445 3785
rect 9785 3595 9845 3785
rect 10185 3595 10245 3785
rect 10585 3595 10645 3785
rect 10985 3595 11045 3785
rect 11385 3595 11445 3785
rect 11785 3595 11845 3785
rect 12185 3595 12245 3785
rect 12585 3595 12645 3785
rect 12985 3595 13045 3785
rect -225 3590 -145 3595
rect -225 3530 -215 3590
rect -155 3530 -145 3590
rect -225 3480 -145 3530
rect -225 3420 -215 3480
rect -155 3420 -145 3480
rect -225 3415 -145 3420
rect 175 3590 255 3595
rect 175 3530 185 3590
rect 245 3530 255 3590
rect 175 3480 255 3530
rect 175 3420 185 3480
rect 245 3420 255 3480
rect 175 3415 255 3420
rect 575 3590 655 3595
rect 575 3530 585 3590
rect 645 3530 655 3590
rect 575 3480 655 3530
rect 575 3420 585 3480
rect 645 3420 655 3480
rect 575 3415 655 3420
rect 975 3590 1055 3595
rect 975 3530 985 3590
rect 1045 3530 1055 3590
rect 975 3480 1055 3530
rect 975 3420 985 3480
rect 1045 3420 1055 3480
rect 975 3415 1055 3420
rect 1375 3590 1455 3595
rect 1375 3530 1385 3590
rect 1445 3530 1455 3590
rect 1375 3480 1455 3530
rect 1375 3420 1385 3480
rect 1445 3420 1455 3480
rect 1375 3415 1455 3420
rect 1775 3590 1855 3595
rect 1775 3530 1785 3590
rect 1845 3530 1855 3590
rect 1775 3480 1855 3530
rect 1775 3420 1785 3480
rect 1845 3420 1855 3480
rect 1775 3415 1855 3420
rect 2175 3590 2255 3595
rect 2175 3530 2185 3590
rect 2245 3530 2255 3590
rect 2175 3480 2255 3530
rect 2175 3420 2185 3480
rect 2245 3420 2255 3480
rect 2175 3415 2255 3420
rect 2575 3590 2655 3595
rect 2575 3530 2585 3590
rect 2645 3530 2655 3590
rect 2575 3480 2655 3530
rect 2575 3420 2585 3480
rect 2645 3420 2655 3480
rect 2575 3415 2655 3420
rect 2975 3590 3055 3595
rect 2975 3530 2985 3590
rect 3045 3530 3055 3590
rect 2975 3480 3055 3530
rect 2975 3420 2985 3480
rect 3045 3420 3055 3480
rect 2975 3415 3055 3420
rect 3375 3590 3455 3595
rect 3375 3530 3385 3590
rect 3445 3530 3455 3590
rect 3375 3480 3455 3530
rect 3375 3420 3385 3480
rect 3445 3420 3455 3480
rect 3375 3415 3455 3420
rect 3775 3590 3855 3595
rect 3775 3530 3785 3590
rect 3845 3530 3855 3590
rect 3775 3480 3855 3530
rect 3775 3420 3785 3480
rect 3845 3420 3855 3480
rect 3775 3415 3855 3420
rect 4175 3590 4255 3595
rect 4175 3530 4185 3590
rect 4245 3530 4255 3590
rect 4175 3480 4255 3530
rect 4175 3420 4185 3480
rect 4245 3420 4255 3480
rect 4175 3415 4255 3420
rect 4575 3590 4655 3595
rect 4575 3530 4585 3590
rect 4645 3530 4655 3590
rect 4575 3480 4655 3530
rect 4575 3420 4585 3480
rect 4645 3420 4655 3480
rect 4575 3415 4655 3420
rect 4975 3590 5055 3595
rect 4975 3530 4985 3590
rect 5045 3530 5055 3590
rect 4975 3480 5055 3530
rect 4975 3420 4985 3480
rect 5045 3420 5055 3480
rect 4975 3415 5055 3420
rect 5375 3590 5455 3595
rect 5375 3530 5385 3590
rect 5445 3530 5455 3590
rect 5375 3480 5455 3530
rect 5375 3420 5385 3480
rect 5445 3420 5455 3480
rect 5375 3415 5455 3420
rect 5775 3590 5855 3595
rect 5775 3530 5785 3590
rect 5845 3530 5855 3590
rect 5775 3480 5855 3530
rect 5775 3420 5785 3480
rect 5845 3420 5855 3480
rect 5775 3415 5855 3420
rect 6175 3590 6255 3595
rect 6175 3530 6185 3590
rect 6245 3530 6255 3590
rect 6175 3480 6255 3530
rect 6175 3420 6185 3480
rect 6245 3420 6255 3480
rect 6175 3415 6255 3420
rect 6575 3590 6655 3595
rect 6575 3530 6585 3590
rect 6645 3530 6655 3590
rect 6575 3480 6655 3530
rect 6575 3420 6585 3480
rect 6645 3420 6655 3480
rect 6575 3415 6655 3420
rect 6975 3590 7055 3595
rect 6975 3530 6985 3590
rect 7045 3530 7055 3590
rect 6975 3480 7055 3530
rect 6975 3420 6985 3480
rect 7045 3420 7055 3480
rect 6975 3415 7055 3420
rect 7375 3590 7455 3595
rect 7375 3530 7385 3590
rect 7445 3530 7455 3590
rect 7375 3480 7455 3530
rect 7375 3420 7385 3480
rect 7445 3420 7455 3480
rect 7375 3415 7455 3420
rect 7775 3590 7855 3595
rect 7775 3530 7785 3590
rect 7845 3530 7855 3590
rect 7775 3480 7855 3530
rect 7775 3420 7785 3480
rect 7845 3420 7855 3480
rect 7775 3415 7855 3420
rect 8175 3590 8255 3595
rect 8175 3530 8185 3590
rect 8245 3530 8255 3590
rect 8175 3480 8255 3530
rect 8175 3420 8185 3480
rect 8245 3420 8255 3480
rect 8175 3415 8255 3420
rect 8575 3590 8655 3595
rect 8575 3530 8585 3590
rect 8645 3530 8655 3590
rect 8575 3480 8655 3530
rect 8575 3420 8585 3480
rect 8645 3420 8655 3480
rect 8575 3415 8655 3420
rect 8975 3590 9055 3595
rect 8975 3530 8985 3590
rect 9045 3530 9055 3590
rect 8975 3480 9055 3530
rect 8975 3420 8985 3480
rect 9045 3420 9055 3480
rect 8975 3415 9055 3420
rect 9375 3590 9455 3595
rect 9375 3530 9385 3590
rect 9445 3530 9455 3590
rect 9375 3480 9455 3530
rect 9375 3420 9385 3480
rect 9445 3420 9455 3480
rect 9375 3415 9455 3420
rect 9775 3590 9855 3595
rect 9775 3530 9785 3590
rect 9845 3530 9855 3590
rect 9775 3480 9855 3530
rect 9775 3420 9785 3480
rect 9845 3420 9855 3480
rect 9775 3415 9855 3420
rect 10175 3590 10255 3595
rect 10175 3530 10185 3590
rect 10245 3530 10255 3590
rect 10175 3480 10255 3530
rect 10175 3420 10185 3480
rect 10245 3420 10255 3480
rect 10175 3415 10255 3420
rect 10575 3590 10655 3595
rect 10575 3530 10585 3590
rect 10645 3530 10655 3590
rect 10575 3480 10655 3530
rect 10575 3420 10585 3480
rect 10645 3420 10655 3480
rect 10575 3415 10655 3420
rect 10975 3590 11055 3595
rect 10975 3530 10985 3590
rect 11045 3530 11055 3590
rect 10975 3480 11055 3530
rect 10975 3420 10985 3480
rect 11045 3420 11055 3480
rect 10975 3415 11055 3420
rect 11375 3590 11455 3595
rect 11375 3530 11385 3590
rect 11445 3530 11455 3590
rect 11375 3480 11455 3530
rect 11375 3420 11385 3480
rect 11445 3420 11455 3480
rect 11375 3415 11455 3420
rect 11775 3590 11855 3595
rect 11775 3530 11785 3590
rect 11845 3530 11855 3590
rect 11775 3480 11855 3530
rect 11775 3420 11785 3480
rect 11845 3420 11855 3480
rect 11775 3415 11855 3420
rect 12175 3590 12255 3595
rect 12175 3530 12185 3590
rect 12245 3530 12255 3590
rect 12175 3480 12255 3530
rect 12175 3420 12185 3480
rect 12245 3420 12255 3480
rect 12175 3415 12255 3420
rect 12575 3590 12655 3595
rect 12575 3530 12585 3590
rect 12645 3530 12655 3590
rect 12575 3480 12655 3530
rect 12575 3420 12585 3480
rect 12645 3420 12655 3480
rect 12575 3415 12655 3420
rect 12975 3590 13055 3595
rect 12975 3530 12985 3590
rect 13045 3530 13055 3590
rect 12975 3480 13055 3530
rect 12975 3420 12985 3480
rect 13045 3420 13055 3480
rect 12975 3415 13055 3420
rect -215 3225 -155 3415
rect 185 3225 245 3415
rect 585 3225 645 3415
rect 985 3225 1045 3415
rect 1385 3225 1445 3415
rect 1785 3225 1845 3415
rect 2185 3225 2245 3415
rect 2585 3225 2645 3415
rect 2985 3225 3045 3415
rect 3385 3225 3445 3415
rect 3785 3225 3845 3415
rect 4185 3225 4245 3415
rect 4585 3225 4645 3415
rect 4985 3225 5045 3415
rect 5385 3225 5445 3415
rect 5785 3225 5845 3415
rect 6185 3225 6245 3415
rect 6585 3225 6645 3415
rect 6985 3225 7045 3415
rect 7385 3225 7445 3415
rect 7785 3225 7845 3415
rect 8185 3225 8245 3415
rect 8585 3225 8645 3415
rect 8985 3225 9045 3415
rect 9385 3225 9445 3415
rect 9785 3225 9845 3415
rect 10185 3225 10245 3415
rect 10585 3225 10645 3415
rect 10985 3225 11045 3415
rect 11385 3225 11445 3415
rect 11785 3225 11845 3415
rect 12185 3225 12245 3415
rect 12585 3225 12645 3415
rect 12985 3225 13045 3415
rect -225 3220 -145 3225
rect -225 3160 -215 3220
rect -155 3160 -145 3220
rect -225 3110 -145 3160
rect -225 3050 -215 3110
rect -155 3050 -145 3110
rect -225 3045 -145 3050
rect 175 3220 255 3225
rect 175 3160 185 3220
rect 245 3160 255 3220
rect 175 3110 255 3160
rect 175 3050 185 3110
rect 245 3050 255 3110
rect 175 3045 255 3050
rect 575 3220 655 3225
rect 575 3160 585 3220
rect 645 3160 655 3220
rect 575 3110 655 3160
rect 575 3050 585 3110
rect 645 3050 655 3110
rect 575 3045 655 3050
rect 975 3220 1055 3225
rect 975 3160 985 3220
rect 1045 3160 1055 3220
rect 975 3110 1055 3160
rect 975 3050 985 3110
rect 1045 3050 1055 3110
rect 975 3045 1055 3050
rect 1375 3220 1455 3225
rect 1375 3160 1385 3220
rect 1445 3160 1455 3220
rect 1375 3110 1455 3160
rect 1375 3050 1385 3110
rect 1445 3050 1455 3110
rect 1375 3045 1455 3050
rect 1775 3220 1855 3225
rect 1775 3160 1785 3220
rect 1845 3160 1855 3220
rect 1775 3110 1855 3160
rect 1775 3050 1785 3110
rect 1845 3050 1855 3110
rect 1775 3045 1855 3050
rect 2175 3220 2255 3225
rect 2175 3160 2185 3220
rect 2245 3160 2255 3220
rect 2175 3110 2255 3160
rect 2175 3050 2185 3110
rect 2245 3050 2255 3110
rect 2175 3045 2255 3050
rect 2575 3220 2655 3225
rect 2575 3160 2585 3220
rect 2645 3160 2655 3220
rect 2575 3110 2655 3160
rect 2575 3050 2585 3110
rect 2645 3050 2655 3110
rect 2575 3045 2655 3050
rect 2975 3220 3055 3225
rect 2975 3160 2985 3220
rect 3045 3160 3055 3220
rect 2975 3110 3055 3160
rect 2975 3050 2985 3110
rect 3045 3050 3055 3110
rect 2975 3045 3055 3050
rect 3375 3220 3455 3225
rect 3375 3160 3385 3220
rect 3445 3160 3455 3220
rect 3375 3110 3455 3160
rect 3375 3050 3385 3110
rect 3445 3050 3455 3110
rect 3375 3045 3455 3050
rect 3775 3220 3855 3225
rect 3775 3160 3785 3220
rect 3845 3160 3855 3220
rect 3775 3110 3855 3160
rect 3775 3050 3785 3110
rect 3845 3050 3855 3110
rect 3775 3045 3855 3050
rect 4175 3220 4255 3225
rect 4175 3160 4185 3220
rect 4245 3160 4255 3220
rect 4175 3110 4255 3160
rect 4175 3050 4185 3110
rect 4245 3050 4255 3110
rect 4175 3045 4255 3050
rect 4575 3220 4655 3225
rect 4575 3160 4585 3220
rect 4645 3160 4655 3220
rect 4575 3110 4655 3160
rect 4575 3050 4585 3110
rect 4645 3050 4655 3110
rect 4575 3045 4655 3050
rect 4975 3220 5055 3225
rect 4975 3160 4985 3220
rect 5045 3160 5055 3220
rect 4975 3110 5055 3160
rect 4975 3050 4985 3110
rect 5045 3050 5055 3110
rect 4975 3045 5055 3050
rect 5375 3220 5455 3225
rect 5375 3160 5385 3220
rect 5445 3160 5455 3220
rect 5375 3110 5455 3160
rect 5375 3050 5385 3110
rect 5445 3050 5455 3110
rect 5375 3045 5455 3050
rect 5775 3220 5855 3225
rect 5775 3160 5785 3220
rect 5845 3160 5855 3220
rect 5775 3110 5855 3160
rect 5775 3050 5785 3110
rect 5845 3050 5855 3110
rect 5775 3045 5855 3050
rect 6175 3220 6255 3225
rect 6175 3160 6185 3220
rect 6245 3160 6255 3220
rect 6175 3110 6255 3160
rect 6175 3050 6185 3110
rect 6245 3050 6255 3110
rect 6175 3045 6255 3050
rect 6575 3220 6655 3225
rect 6575 3160 6585 3220
rect 6645 3160 6655 3220
rect 6575 3110 6655 3160
rect 6575 3050 6585 3110
rect 6645 3050 6655 3110
rect 6575 3045 6655 3050
rect 6975 3220 7055 3225
rect 6975 3160 6985 3220
rect 7045 3160 7055 3220
rect 6975 3110 7055 3160
rect 6975 3050 6985 3110
rect 7045 3050 7055 3110
rect 6975 3045 7055 3050
rect 7375 3220 7455 3225
rect 7375 3160 7385 3220
rect 7445 3160 7455 3220
rect 7375 3110 7455 3160
rect 7375 3050 7385 3110
rect 7445 3050 7455 3110
rect 7375 3045 7455 3050
rect 7775 3220 7855 3225
rect 7775 3160 7785 3220
rect 7845 3160 7855 3220
rect 7775 3110 7855 3160
rect 7775 3050 7785 3110
rect 7845 3050 7855 3110
rect 7775 3045 7855 3050
rect 8175 3220 8255 3225
rect 8175 3160 8185 3220
rect 8245 3160 8255 3220
rect 8175 3110 8255 3160
rect 8175 3050 8185 3110
rect 8245 3050 8255 3110
rect 8175 3045 8255 3050
rect 8575 3220 8655 3225
rect 8575 3160 8585 3220
rect 8645 3160 8655 3220
rect 8575 3110 8655 3160
rect 8575 3050 8585 3110
rect 8645 3050 8655 3110
rect 8575 3045 8655 3050
rect 8975 3220 9055 3225
rect 8975 3160 8985 3220
rect 9045 3160 9055 3220
rect 8975 3110 9055 3160
rect 8975 3050 8985 3110
rect 9045 3050 9055 3110
rect 8975 3045 9055 3050
rect 9375 3220 9455 3225
rect 9375 3160 9385 3220
rect 9445 3160 9455 3220
rect 9375 3110 9455 3160
rect 9375 3050 9385 3110
rect 9445 3050 9455 3110
rect 9375 3045 9455 3050
rect 9775 3220 9855 3225
rect 9775 3160 9785 3220
rect 9845 3160 9855 3220
rect 9775 3110 9855 3160
rect 9775 3050 9785 3110
rect 9845 3050 9855 3110
rect 9775 3045 9855 3050
rect 10175 3220 10255 3225
rect 10175 3160 10185 3220
rect 10245 3160 10255 3220
rect 10175 3110 10255 3160
rect 10175 3050 10185 3110
rect 10245 3050 10255 3110
rect 10175 3045 10255 3050
rect 10575 3220 10655 3225
rect 10575 3160 10585 3220
rect 10645 3160 10655 3220
rect 10575 3110 10655 3160
rect 10575 3050 10585 3110
rect 10645 3050 10655 3110
rect 10575 3045 10655 3050
rect 10975 3220 11055 3225
rect 10975 3160 10985 3220
rect 11045 3160 11055 3220
rect 10975 3110 11055 3160
rect 10975 3050 10985 3110
rect 11045 3050 11055 3110
rect 10975 3045 11055 3050
rect 11375 3220 11455 3225
rect 11375 3160 11385 3220
rect 11445 3160 11455 3220
rect 11375 3110 11455 3160
rect 11375 3050 11385 3110
rect 11445 3050 11455 3110
rect 11375 3045 11455 3050
rect 11775 3220 11855 3225
rect 11775 3160 11785 3220
rect 11845 3160 11855 3220
rect 11775 3110 11855 3160
rect 11775 3050 11785 3110
rect 11845 3050 11855 3110
rect 11775 3045 11855 3050
rect 12175 3220 12255 3225
rect 12175 3160 12185 3220
rect 12245 3160 12255 3220
rect 12175 3110 12255 3160
rect 12175 3050 12185 3110
rect 12245 3050 12255 3110
rect 12175 3045 12255 3050
rect 12575 3220 12655 3225
rect 12575 3160 12585 3220
rect 12645 3160 12655 3220
rect 12575 3110 12655 3160
rect 12575 3050 12585 3110
rect 12645 3050 12655 3110
rect 12575 3045 12655 3050
rect 12975 3220 13055 3225
rect 12975 3160 12985 3220
rect 13045 3160 13055 3220
rect 12975 3110 13055 3160
rect 12975 3050 12985 3110
rect 13045 3050 13055 3110
rect 12975 3045 13055 3050
rect -215 2855 -155 3045
rect 185 2855 245 3045
rect 585 2855 645 3045
rect 985 2855 1045 3045
rect 1385 2855 1445 3045
rect 1785 2855 1845 3045
rect 2185 2855 2245 3045
rect 2585 2855 2645 3045
rect 2985 2855 3045 3045
rect 3385 2855 3445 3045
rect 3785 2855 3845 3045
rect 4185 2855 4245 3045
rect 4585 2855 4645 3045
rect 4985 2855 5045 3045
rect 5385 2855 5445 3045
rect 5785 2855 5845 3045
rect 6185 2855 6245 3045
rect 6585 2855 6645 3045
rect 6985 2855 7045 3045
rect 7385 2855 7445 3045
rect 7785 2855 7845 3045
rect 8185 2855 8245 3045
rect 8585 2855 8645 3045
rect 8985 2855 9045 3045
rect 9385 2855 9445 3045
rect 9785 2855 9845 3045
rect 10185 2855 10245 3045
rect 10585 2855 10645 3045
rect 10985 2855 11045 3045
rect 11385 2855 11445 3045
rect 11785 2855 11845 3045
rect 12185 2855 12245 3045
rect 12585 2855 12645 3045
rect 12985 2855 13045 3045
rect -225 2850 -145 2855
rect -225 2790 -215 2850
rect -155 2790 -145 2850
rect -225 2740 -145 2790
rect -225 2680 -215 2740
rect -155 2680 -145 2740
rect -225 2675 -145 2680
rect 175 2850 255 2855
rect 175 2790 185 2850
rect 245 2790 255 2850
rect 175 2740 255 2790
rect 175 2680 185 2740
rect 245 2680 255 2740
rect 175 2675 255 2680
rect 575 2850 655 2855
rect 575 2790 585 2850
rect 645 2790 655 2850
rect 575 2740 655 2790
rect 575 2680 585 2740
rect 645 2680 655 2740
rect 575 2675 655 2680
rect 975 2850 1055 2855
rect 975 2790 985 2850
rect 1045 2790 1055 2850
rect 975 2740 1055 2790
rect 975 2680 985 2740
rect 1045 2680 1055 2740
rect 975 2675 1055 2680
rect 1375 2850 1455 2855
rect 1375 2790 1385 2850
rect 1445 2790 1455 2850
rect 1375 2740 1455 2790
rect 1375 2680 1385 2740
rect 1445 2680 1455 2740
rect 1375 2675 1455 2680
rect 1775 2850 1855 2855
rect 1775 2790 1785 2850
rect 1845 2790 1855 2850
rect 1775 2740 1855 2790
rect 1775 2680 1785 2740
rect 1845 2680 1855 2740
rect 1775 2675 1855 2680
rect 2175 2850 2255 2855
rect 2175 2790 2185 2850
rect 2245 2790 2255 2850
rect 2175 2740 2255 2790
rect 2175 2680 2185 2740
rect 2245 2680 2255 2740
rect 2175 2675 2255 2680
rect 2575 2850 2655 2855
rect 2575 2790 2585 2850
rect 2645 2790 2655 2850
rect 2575 2740 2655 2790
rect 2575 2680 2585 2740
rect 2645 2680 2655 2740
rect 2575 2675 2655 2680
rect 2975 2850 3055 2855
rect 2975 2790 2985 2850
rect 3045 2790 3055 2850
rect 2975 2740 3055 2790
rect 2975 2680 2985 2740
rect 3045 2680 3055 2740
rect 2975 2675 3055 2680
rect 3375 2850 3455 2855
rect 3375 2790 3385 2850
rect 3445 2790 3455 2850
rect 3375 2740 3455 2790
rect 3375 2680 3385 2740
rect 3445 2680 3455 2740
rect 3375 2675 3455 2680
rect 3775 2850 3855 2855
rect 3775 2790 3785 2850
rect 3845 2790 3855 2850
rect 3775 2740 3855 2790
rect 3775 2680 3785 2740
rect 3845 2680 3855 2740
rect 3775 2675 3855 2680
rect 4175 2850 4255 2855
rect 4175 2790 4185 2850
rect 4245 2790 4255 2850
rect 4175 2740 4255 2790
rect 4175 2680 4185 2740
rect 4245 2680 4255 2740
rect 4175 2675 4255 2680
rect 4575 2850 4655 2855
rect 4575 2790 4585 2850
rect 4645 2790 4655 2850
rect 4575 2740 4655 2790
rect 4575 2680 4585 2740
rect 4645 2680 4655 2740
rect 4575 2675 4655 2680
rect 4975 2850 5055 2855
rect 4975 2790 4985 2850
rect 5045 2790 5055 2850
rect 4975 2740 5055 2790
rect 4975 2680 4985 2740
rect 5045 2680 5055 2740
rect 4975 2675 5055 2680
rect 5375 2850 5455 2855
rect 5375 2790 5385 2850
rect 5445 2790 5455 2850
rect 5375 2740 5455 2790
rect 5375 2680 5385 2740
rect 5445 2680 5455 2740
rect 5375 2675 5455 2680
rect 5775 2850 5855 2855
rect 5775 2790 5785 2850
rect 5845 2790 5855 2850
rect 5775 2740 5855 2790
rect 5775 2680 5785 2740
rect 5845 2680 5855 2740
rect 5775 2675 5855 2680
rect 6175 2850 6255 2855
rect 6175 2790 6185 2850
rect 6245 2790 6255 2850
rect 6175 2740 6255 2790
rect 6175 2680 6185 2740
rect 6245 2680 6255 2740
rect 6175 2675 6255 2680
rect 6575 2850 6655 2855
rect 6575 2790 6585 2850
rect 6645 2790 6655 2850
rect 6575 2740 6655 2790
rect 6575 2680 6585 2740
rect 6645 2680 6655 2740
rect 6575 2675 6655 2680
rect 6975 2850 7055 2855
rect 6975 2790 6985 2850
rect 7045 2790 7055 2850
rect 6975 2740 7055 2790
rect 6975 2680 6985 2740
rect 7045 2680 7055 2740
rect 6975 2675 7055 2680
rect 7375 2850 7455 2855
rect 7375 2790 7385 2850
rect 7445 2790 7455 2850
rect 7375 2740 7455 2790
rect 7375 2680 7385 2740
rect 7445 2680 7455 2740
rect 7375 2675 7455 2680
rect 7775 2850 7855 2855
rect 7775 2790 7785 2850
rect 7845 2790 7855 2850
rect 7775 2740 7855 2790
rect 7775 2680 7785 2740
rect 7845 2680 7855 2740
rect 7775 2675 7855 2680
rect 8175 2850 8255 2855
rect 8175 2790 8185 2850
rect 8245 2790 8255 2850
rect 8175 2740 8255 2790
rect 8175 2680 8185 2740
rect 8245 2680 8255 2740
rect 8175 2675 8255 2680
rect 8575 2850 8655 2855
rect 8575 2790 8585 2850
rect 8645 2790 8655 2850
rect 8575 2740 8655 2790
rect 8575 2680 8585 2740
rect 8645 2680 8655 2740
rect 8575 2675 8655 2680
rect 8975 2850 9055 2855
rect 8975 2790 8985 2850
rect 9045 2790 9055 2850
rect 8975 2740 9055 2790
rect 8975 2680 8985 2740
rect 9045 2680 9055 2740
rect 8975 2675 9055 2680
rect 9375 2850 9455 2855
rect 9375 2790 9385 2850
rect 9445 2790 9455 2850
rect 9375 2740 9455 2790
rect 9375 2680 9385 2740
rect 9445 2680 9455 2740
rect 9375 2675 9455 2680
rect 9775 2850 9855 2855
rect 9775 2790 9785 2850
rect 9845 2790 9855 2850
rect 9775 2740 9855 2790
rect 9775 2680 9785 2740
rect 9845 2680 9855 2740
rect 9775 2675 9855 2680
rect 10175 2850 10255 2855
rect 10175 2790 10185 2850
rect 10245 2790 10255 2850
rect 10175 2740 10255 2790
rect 10175 2680 10185 2740
rect 10245 2680 10255 2740
rect 10175 2675 10255 2680
rect 10575 2850 10655 2855
rect 10575 2790 10585 2850
rect 10645 2790 10655 2850
rect 10575 2740 10655 2790
rect 10575 2680 10585 2740
rect 10645 2680 10655 2740
rect 10575 2675 10655 2680
rect 10975 2850 11055 2855
rect 10975 2790 10985 2850
rect 11045 2790 11055 2850
rect 10975 2740 11055 2790
rect 10975 2680 10985 2740
rect 11045 2680 11055 2740
rect 10975 2675 11055 2680
rect 11375 2850 11455 2855
rect 11375 2790 11385 2850
rect 11445 2790 11455 2850
rect 11375 2740 11455 2790
rect 11375 2680 11385 2740
rect 11445 2680 11455 2740
rect 11375 2675 11455 2680
rect 11775 2850 11855 2855
rect 11775 2790 11785 2850
rect 11845 2790 11855 2850
rect 11775 2740 11855 2790
rect 11775 2680 11785 2740
rect 11845 2680 11855 2740
rect 11775 2675 11855 2680
rect 12175 2850 12255 2855
rect 12175 2790 12185 2850
rect 12245 2790 12255 2850
rect 12175 2740 12255 2790
rect 12175 2680 12185 2740
rect 12245 2680 12255 2740
rect 12175 2675 12255 2680
rect 12575 2850 12655 2855
rect 12575 2790 12585 2850
rect 12645 2790 12655 2850
rect 12575 2740 12655 2790
rect 12575 2680 12585 2740
rect 12645 2680 12655 2740
rect 12575 2675 12655 2680
rect 12975 2850 13055 2855
rect 12975 2790 12985 2850
rect 13045 2790 13055 2850
rect 12975 2740 13055 2790
rect 12975 2680 12985 2740
rect 13045 2680 13055 2740
rect 12975 2675 13055 2680
rect -215 2485 -155 2675
rect 185 2485 245 2675
rect 585 2485 645 2675
rect 985 2485 1045 2675
rect 1385 2485 1445 2675
rect 1785 2485 1845 2675
rect 2185 2485 2245 2675
rect 2585 2485 2645 2675
rect 2985 2485 3045 2675
rect 3385 2485 3445 2675
rect 3785 2485 3845 2675
rect 4185 2485 4245 2675
rect 4585 2485 4645 2675
rect 4985 2485 5045 2675
rect 5385 2485 5445 2675
rect 5785 2485 5845 2675
rect 6185 2485 6245 2675
rect 6585 2485 6645 2675
rect 6985 2485 7045 2675
rect 7385 2485 7445 2675
rect 7785 2485 7845 2675
rect 8185 2485 8245 2675
rect 8585 2485 8645 2675
rect 8985 2485 9045 2675
rect 9385 2485 9445 2675
rect 9785 2485 9845 2675
rect 10185 2485 10245 2675
rect 10585 2485 10645 2675
rect 10985 2485 11045 2675
rect 11385 2485 11445 2675
rect 11785 2485 11845 2675
rect 12185 2485 12245 2675
rect 12585 2485 12645 2675
rect 12985 2485 13045 2675
rect -225 2480 -145 2485
rect -225 2420 -215 2480
rect -155 2420 -145 2480
rect -225 2370 -145 2420
rect -225 2310 -215 2370
rect -155 2310 -145 2370
rect -225 2305 -145 2310
rect 175 2480 255 2485
rect 175 2420 185 2480
rect 245 2420 255 2480
rect 175 2370 255 2420
rect 175 2310 185 2370
rect 245 2310 255 2370
rect 175 2305 255 2310
rect 575 2480 655 2485
rect 575 2420 585 2480
rect 645 2420 655 2480
rect 575 2370 655 2420
rect 575 2310 585 2370
rect 645 2310 655 2370
rect 575 2305 655 2310
rect 975 2480 1055 2485
rect 975 2420 985 2480
rect 1045 2420 1055 2480
rect 975 2370 1055 2420
rect 975 2310 985 2370
rect 1045 2310 1055 2370
rect 975 2305 1055 2310
rect 1375 2480 1455 2485
rect 1375 2420 1385 2480
rect 1445 2420 1455 2480
rect 1375 2370 1455 2420
rect 1375 2310 1385 2370
rect 1445 2310 1455 2370
rect 1375 2305 1455 2310
rect 1775 2480 1855 2485
rect 1775 2420 1785 2480
rect 1845 2420 1855 2480
rect 1775 2370 1855 2420
rect 1775 2310 1785 2370
rect 1845 2310 1855 2370
rect 1775 2305 1855 2310
rect 2175 2480 2255 2485
rect 2175 2420 2185 2480
rect 2245 2420 2255 2480
rect 2175 2370 2255 2420
rect 2175 2310 2185 2370
rect 2245 2310 2255 2370
rect 2175 2305 2255 2310
rect 2575 2480 2655 2485
rect 2575 2420 2585 2480
rect 2645 2420 2655 2480
rect 2575 2370 2655 2420
rect 2575 2310 2585 2370
rect 2645 2310 2655 2370
rect 2575 2305 2655 2310
rect 2975 2480 3055 2485
rect 2975 2420 2985 2480
rect 3045 2420 3055 2480
rect 2975 2370 3055 2420
rect 2975 2310 2985 2370
rect 3045 2310 3055 2370
rect 2975 2305 3055 2310
rect 3375 2480 3455 2485
rect 3375 2420 3385 2480
rect 3445 2420 3455 2480
rect 3375 2370 3455 2420
rect 3375 2310 3385 2370
rect 3445 2310 3455 2370
rect 3375 2305 3455 2310
rect 3775 2480 3855 2485
rect 3775 2420 3785 2480
rect 3845 2420 3855 2480
rect 3775 2370 3855 2420
rect 3775 2310 3785 2370
rect 3845 2310 3855 2370
rect 3775 2305 3855 2310
rect 4175 2480 4255 2485
rect 4175 2420 4185 2480
rect 4245 2420 4255 2480
rect 4175 2370 4255 2420
rect 4175 2310 4185 2370
rect 4245 2310 4255 2370
rect 4175 2305 4255 2310
rect 4575 2480 4655 2485
rect 4575 2420 4585 2480
rect 4645 2420 4655 2480
rect 4575 2370 4655 2420
rect 4575 2310 4585 2370
rect 4645 2310 4655 2370
rect 4575 2305 4655 2310
rect 4975 2480 5055 2485
rect 4975 2420 4985 2480
rect 5045 2420 5055 2480
rect 4975 2370 5055 2420
rect 4975 2310 4985 2370
rect 5045 2310 5055 2370
rect 4975 2305 5055 2310
rect 5375 2480 5455 2485
rect 5375 2420 5385 2480
rect 5445 2420 5455 2480
rect 5375 2370 5455 2420
rect 5375 2310 5385 2370
rect 5445 2310 5455 2370
rect 5375 2305 5455 2310
rect 5775 2480 5855 2485
rect 5775 2420 5785 2480
rect 5845 2420 5855 2480
rect 5775 2370 5855 2420
rect 5775 2310 5785 2370
rect 5845 2310 5855 2370
rect 5775 2305 5855 2310
rect 6175 2480 6255 2485
rect 6175 2420 6185 2480
rect 6245 2420 6255 2480
rect 6175 2370 6255 2420
rect 6175 2310 6185 2370
rect 6245 2310 6255 2370
rect 6175 2305 6255 2310
rect 6575 2480 6655 2485
rect 6575 2420 6585 2480
rect 6645 2420 6655 2480
rect 6575 2370 6655 2420
rect 6575 2310 6585 2370
rect 6645 2310 6655 2370
rect 6575 2305 6655 2310
rect 6975 2480 7055 2485
rect 6975 2420 6985 2480
rect 7045 2420 7055 2480
rect 6975 2370 7055 2420
rect 6975 2310 6985 2370
rect 7045 2310 7055 2370
rect 6975 2305 7055 2310
rect 7375 2480 7455 2485
rect 7375 2420 7385 2480
rect 7445 2420 7455 2480
rect 7375 2370 7455 2420
rect 7375 2310 7385 2370
rect 7445 2310 7455 2370
rect 7375 2305 7455 2310
rect 7775 2480 7855 2485
rect 7775 2420 7785 2480
rect 7845 2420 7855 2480
rect 7775 2370 7855 2420
rect 7775 2310 7785 2370
rect 7845 2310 7855 2370
rect 7775 2305 7855 2310
rect 8175 2480 8255 2485
rect 8175 2420 8185 2480
rect 8245 2420 8255 2480
rect 8175 2370 8255 2420
rect 8175 2310 8185 2370
rect 8245 2310 8255 2370
rect 8175 2305 8255 2310
rect 8575 2480 8655 2485
rect 8575 2420 8585 2480
rect 8645 2420 8655 2480
rect 8575 2370 8655 2420
rect 8575 2310 8585 2370
rect 8645 2310 8655 2370
rect 8575 2305 8655 2310
rect 8975 2480 9055 2485
rect 8975 2420 8985 2480
rect 9045 2420 9055 2480
rect 8975 2370 9055 2420
rect 8975 2310 8985 2370
rect 9045 2310 9055 2370
rect 8975 2305 9055 2310
rect 9375 2480 9455 2485
rect 9375 2420 9385 2480
rect 9445 2420 9455 2480
rect 9375 2370 9455 2420
rect 9375 2310 9385 2370
rect 9445 2310 9455 2370
rect 9375 2305 9455 2310
rect 9775 2480 9855 2485
rect 9775 2420 9785 2480
rect 9845 2420 9855 2480
rect 9775 2370 9855 2420
rect 9775 2310 9785 2370
rect 9845 2310 9855 2370
rect 9775 2305 9855 2310
rect 10175 2480 10255 2485
rect 10175 2420 10185 2480
rect 10245 2420 10255 2480
rect 10175 2370 10255 2420
rect 10175 2310 10185 2370
rect 10245 2310 10255 2370
rect 10175 2305 10255 2310
rect 10575 2480 10655 2485
rect 10575 2420 10585 2480
rect 10645 2420 10655 2480
rect 10575 2370 10655 2420
rect 10575 2310 10585 2370
rect 10645 2310 10655 2370
rect 10575 2305 10655 2310
rect 10975 2480 11055 2485
rect 10975 2420 10985 2480
rect 11045 2420 11055 2480
rect 10975 2370 11055 2420
rect 10975 2310 10985 2370
rect 11045 2310 11055 2370
rect 10975 2305 11055 2310
rect 11375 2480 11455 2485
rect 11375 2420 11385 2480
rect 11445 2420 11455 2480
rect 11375 2370 11455 2420
rect 11375 2310 11385 2370
rect 11445 2310 11455 2370
rect 11375 2305 11455 2310
rect 11775 2480 11855 2485
rect 11775 2420 11785 2480
rect 11845 2420 11855 2480
rect 11775 2370 11855 2420
rect 11775 2310 11785 2370
rect 11845 2310 11855 2370
rect 11775 2305 11855 2310
rect 12175 2480 12255 2485
rect 12175 2420 12185 2480
rect 12245 2420 12255 2480
rect 12175 2370 12255 2420
rect 12175 2310 12185 2370
rect 12245 2310 12255 2370
rect 12175 2305 12255 2310
rect 12575 2480 12655 2485
rect 12575 2420 12585 2480
rect 12645 2420 12655 2480
rect 12575 2370 12655 2420
rect 12575 2310 12585 2370
rect 12645 2310 12655 2370
rect 12575 2305 12655 2310
rect 12975 2480 13055 2485
rect 12975 2420 12985 2480
rect 13045 2420 13055 2480
rect 12975 2370 13055 2420
rect 12975 2310 12985 2370
rect 13045 2310 13055 2370
rect 12975 2305 13055 2310
rect -215 2115 -155 2305
rect 185 2115 245 2305
rect 585 2115 645 2305
rect 985 2115 1045 2305
rect 1385 2115 1445 2305
rect 1785 2115 1845 2305
rect 2185 2115 2245 2305
rect 2585 2115 2645 2305
rect 2985 2115 3045 2305
rect 3385 2115 3445 2305
rect 3785 2115 3845 2305
rect 4185 2115 4245 2305
rect 4585 2115 4645 2305
rect 4985 2115 5045 2305
rect 5385 2115 5445 2305
rect 5785 2115 5845 2305
rect 6185 2115 6245 2305
rect 6585 2115 6645 2305
rect 6985 2115 7045 2305
rect 7385 2115 7445 2305
rect 7785 2115 7845 2305
rect 8185 2115 8245 2305
rect 8585 2115 8645 2305
rect 8985 2115 9045 2305
rect 9385 2115 9445 2305
rect 9785 2115 9845 2305
rect 10185 2115 10245 2305
rect 10585 2115 10645 2305
rect 10985 2115 11045 2305
rect 11385 2115 11445 2305
rect 11785 2115 11845 2305
rect 12185 2115 12245 2305
rect 12585 2115 12645 2305
rect 12985 2115 13045 2305
rect -225 2110 -145 2115
rect -225 2050 -215 2110
rect -155 2050 -145 2110
rect -225 2000 -145 2050
rect -225 1940 -215 2000
rect -155 1940 -145 2000
rect -225 1935 -145 1940
rect 175 2110 255 2115
rect 175 2050 185 2110
rect 245 2050 255 2110
rect 175 2000 255 2050
rect 175 1940 185 2000
rect 245 1940 255 2000
rect 175 1935 255 1940
rect 575 2110 655 2115
rect 575 2050 585 2110
rect 645 2050 655 2110
rect 575 2000 655 2050
rect 575 1940 585 2000
rect 645 1940 655 2000
rect 575 1935 655 1940
rect 975 2110 1055 2115
rect 975 2050 985 2110
rect 1045 2050 1055 2110
rect 975 2000 1055 2050
rect 975 1940 985 2000
rect 1045 1940 1055 2000
rect 975 1935 1055 1940
rect 1375 2110 1455 2115
rect 1375 2050 1385 2110
rect 1445 2050 1455 2110
rect 1375 2000 1455 2050
rect 1375 1940 1385 2000
rect 1445 1940 1455 2000
rect 1375 1935 1455 1940
rect 1775 2110 1855 2115
rect 1775 2050 1785 2110
rect 1845 2050 1855 2110
rect 1775 2000 1855 2050
rect 1775 1940 1785 2000
rect 1845 1940 1855 2000
rect 1775 1935 1855 1940
rect 2175 2110 2255 2115
rect 2175 2050 2185 2110
rect 2245 2050 2255 2110
rect 2175 2000 2255 2050
rect 2175 1940 2185 2000
rect 2245 1940 2255 2000
rect 2175 1935 2255 1940
rect 2575 2110 2655 2115
rect 2575 2050 2585 2110
rect 2645 2050 2655 2110
rect 2575 2000 2655 2050
rect 2575 1940 2585 2000
rect 2645 1940 2655 2000
rect 2575 1935 2655 1940
rect 2975 2110 3055 2115
rect 2975 2050 2985 2110
rect 3045 2050 3055 2110
rect 2975 2000 3055 2050
rect 2975 1940 2985 2000
rect 3045 1940 3055 2000
rect 2975 1935 3055 1940
rect 3375 2110 3455 2115
rect 3375 2050 3385 2110
rect 3445 2050 3455 2110
rect 3375 2000 3455 2050
rect 3375 1940 3385 2000
rect 3445 1940 3455 2000
rect 3375 1935 3455 1940
rect 3775 2110 3855 2115
rect 3775 2050 3785 2110
rect 3845 2050 3855 2110
rect 3775 2000 3855 2050
rect 3775 1940 3785 2000
rect 3845 1940 3855 2000
rect 3775 1935 3855 1940
rect 4175 2110 4255 2115
rect 4175 2050 4185 2110
rect 4245 2050 4255 2110
rect 4175 2000 4255 2050
rect 4175 1940 4185 2000
rect 4245 1940 4255 2000
rect 4175 1935 4255 1940
rect 4575 2110 4655 2115
rect 4575 2050 4585 2110
rect 4645 2050 4655 2110
rect 4575 2000 4655 2050
rect 4575 1940 4585 2000
rect 4645 1940 4655 2000
rect 4575 1935 4655 1940
rect 4975 2110 5055 2115
rect 4975 2050 4985 2110
rect 5045 2050 5055 2110
rect 4975 2000 5055 2050
rect 4975 1940 4985 2000
rect 5045 1940 5055 2000
rect 4975 1935 5055 1940
rect 5375 2110 5455 2115
rect 5375 2050 5385 2110
rect 5445 2050 5455 2110
rect 5375 2000 5455 2050
rect 5375 1940 5385 2000
rect 5445 1940 5455 2000
rect 5375 1935 5455 1940
rect 5775 2110 5855 2115
rect 5775 2050 5785 2110
rect 5845 2050 5855 2110
rect 5775 2000 5855 2050
rect 5775 1940 5785 2000
rect 5845 1940 5855 2000
rect 5775 1935 5855 1940
rect 6175 2110 6255 2115
rect 6175 2050 6185 2110
rect 6245 2050 6255 2110
rect 6175 2000 6255 2050
rect 6175 1940 6185 2000
rect 6245 1940 6255 2000
rect 6175 1935 6255 1940
rect 6575 2110 6655 2115
rect 6575 2050 6585 2110
rect 6645 2050 6655 2110
rect 6575 2000 6655 2050
rect 6575 1940 6585 2000
rect 6645 1940 6655 2000
rect 6575 1935 6655 1940
rect 6975 2110 7055 2115
rect 6975 2050 6985 2110
rect 7045 2050 7055 2110
rect 6975 2000 7055 2050
rect 6975 1940 6985 2000
rect 7045 1940 7055 2000
rect 6975 1935 7055 1940
rect 7375 2110 7455 2115
rect 7375 2050 7385 2110
rect 7445 2050 7455 2110
rect 7375 2000 7455 2050
rect 7375 1940 7385 2000
rect 7445 1940 7455 2000
rect 7375 1935 7455 1940
rect 7775 2110 7855 2115
rect 7775 2050 7785 2110
rect 7845 2050 7855 2110
rect 7775 2000 7855 2050
rect 7775 1940 7785 2000
rect 7845 1940 7855 2000
rect 7775 1935 7855 1940
rect 8175 2110 8255 2115
rect 8175 2050 8185 2110
rect 8245 2050 8255 2110
rect 8175 2000 8255 2050
rect 8175 1940 8185 2000
rect 8245 1940 8255 2000
rect 8175 1935 8255 1940
rect 8575 2110 8655 2115
rect 8575 2050 8585 2110
rect 8645 2050 8655 2110
rect 8575 2000 8655 2050
rect 8575 1940 8585 2000
rect 8645 1940 8655 2000
rect 8575 1935 8655 1940
rect 8975 2110 9055 2115
rect 8975 2050 8985 2110
rect 9045 2050 9055 2110
rect 8975 2000 9055 2050
rect 8975 1940 8985 2000
rect 9045 1940 9055 2000
rect 8975 1935 9055 1940
rect 9375 2110 9455 2115
rect 9375 2050 9385 2110
rect 9445 2050 9455 2110
rect 9375 2000 9455 2050
rect 9375 1940 9385 2000
rect 9445 1940 9455 2000
rect 9375 1935 9455 1940
rect 9775 2110 9855 2115
rect 9775 2050 9785 2110
rect 9845 2050 9855 2110
rect 9775 2000 9855 2050
rect 9775 1940 9785 2000
rect 9845 1940 9855 2000
rect 9775 1935 9855 1940
rect 10175 2110 10255 2115
rect 10175 2050 10185 2110
rect 10245 2050 10255 2110
rect 10175 2000 10255 2050
rect 10175 1940 10185 2000
rect 10245 1940 10255 2000
rect 10175 1935 10255 1940
rect 10575 2110 10655 2115
rect 10575 2050 10585 2110
rect 10645 2050 10655 2110
rect 10575 2000 10655 2050
rect 10575 1940 10585 2000
rect 10645 1940 10655 2000
rect 10575 1935 10655 1940
rect 10975 2110 11055 2115
rect 10975 2050 10985 2110
rect 11045 2050 11055 2110
rect 10975 2000 11055 2050
rect 10975 1940 10985 2000
rect 11045 1940 11055 2000
rect 10975 1935 11055 1940
rect 11375 2110 11455 2115
rect 11375 2050 11385 2110
rect 11445 2050 11455 2110
rect 11375 2000 11455 2050
rect 11375 1940 11385 2000
rect 11445 1940 11455 2000
rect 11375 1935 11455 1940
rect 11775 2110 11855 2115
rect 11775 2050 11785 2110
rect 11845 2050 11855 2110
rect 11775 2000 11855 2050
rect 11775 1940 11785 2000
rect 11845 1940 11855 2000
rect 11775 1935 11855 1940
rect 12175 2110 12255 2115
rect 12175 2050 12185 2110
rect 12245 2050 12255 2110
rect 12175 2000 12255 2050
rect 12175 1940 12185 2000
rect 12245 1940 12255 2000
rect 12175 1935 12255 1940
rect 12575 2110 12655 2115
rect 12575 2050 12585 2110
rect 12645 2050 12655 2110
rect 12575 2000 12655 2050
rect 12575 1940 12585 2000
rect 12645 1940 12655 2000
rect 12575 1935 12655 1940
rect 12975 2110 13055 2115
rect 12975 2050 12985 2110
rect 13045 2050 13055 2110
rect 12975 2000 13055 2050
rect 12975 1940 12985 2000
rect 13045 1940 13055 2000
rect 12975 1935 13055 1940
rect -215 1745 -155 1935
rect 185 1745 245 1935
rect 585 1745 645 1935
rect 985 1745 1045 1935
rect 1385 1745 1445 1935
rect 1785 1745 1845 1935
rect 2185 1745 2245 1935
rect 2585 1745 2645 1935
rect 2985 1745 3045 1935
rect 3385 1745 3445 1935
rect 3785 1745 3845 1935
rect 4185 1745 4245 1935
rect 4585 1745 4645 1935
rect 4985 1745 5045 1935
rect 5385 1745 5445 1935
rect 5785 1745 5845 1935
rect 6185 1745 6245 1935
rect 6585 1745 6645 1935
rect 6985 1745 7045 1935
rect 7385 1745 7445 1935
rect 7785 1745 7845 1935
rect 8185 1745 8245 1935
rect 8585 1745 8645 1935
rect 8985 1745 9045 1935
rect 9385 1745 9445 1935
rect 9785 1745 9845 1935
rect 10185 1745 10245 1935
rect 10585 1745 10645 1935
rect 10985 1745 11045 1935
rect 11385 1745 11445 1935
rect 11785 1745 11845 1935
rect 12185 1745 12245 1935
rect 12585 1745 12645 1935
rect 12985 1745 13045 1935
rect -225 1740 -145 1745
rect -225 1680 -215 1740
rect -155 1680 -145 1740
rect -225 1630 -145 1680
rect -225 1570 -215 1630
rect -155 1570 -145 1630
rect -225 1565 -145 1570
rect 175 1740 255 1745
rect 175 1680 185 1740
rect 245 1680 255 1740
rect 175 1630 255 1680
rect 175 1570 185 1630
rect 245 1570 255 1630
rect 175 1565 255 1570
rect 575 1740 655 1745
rect 575 1680 585 1740
rect 645 1680 655 1740
rect 575 1630 655 1680
rect 575 1570 585 1630
rect 645 1570 655 1630
rect 575 1565 655 1570
rect 975 1740 1055 1745
rect 975 1680 985 1740
rect 1045 1680 1055 1740
rect 975 1630 1055 1680
rect 975 1570 985 1630
rect 1045 1570 1055 1630
rect 975 1565 1055 1570
rect 1375 1740 1455 1745
rect 1375 1680 1385 1740
rect 1445 1680 1455 1740
rect 1375 1630 1455 1680
rect 1375 1570 1385 1630
rect 1445 1570 1455 1630
rect 1375 1565 1455 1570
rect 1775 1740 1855 1745
rect 1775 1680 1785 1740
rect 1845 1680 1855 1740
rect 1775 1630 1855 1680
rect 1775 1570 1785 1630
rect 1845 1570 1855 1630
rect 1775 1565 1855 1570
rect 2175 1740 2255 1745
rect 2175 1680 2185 1740
rect 2245 1680 2255 1740
rect 2175 1630 2255 1680
rect 2175 1570 2185 1630
rect 2245 1570 2255 1630
rect 2175 1565 2255 1570
rect 2575 1740 2655 1745
rect 2575 1680 2585 1740
rect 2645 1680 2655 1740
rect 2575 1630 2655 1680
rect 2575 1570 2585 1630
rect 2645 1570 2655 1630
rect 2575 1565 2655 1570
rect 2975 1740 3055 1745
rect 2975 1680 2985 1740
rect 3045 1680 3055 1740
rect 2975 1630 3055 1680
rect 2975 1570 2985 1630
rect 3045 1570 3055 1630
rect 2975 1565 3055 1570
rect 3375 1740 3455 1745
rect 3375 1680 3385 1740
rect 3445 1680 3455 1740
rect 3375 1630 3455 1680
rect 3375 1570 3385 1630
rect 3445 1570 3455 1630
rect 3375 1565 3455 1570
rect 3775 1740 3855 1745
rect 3775 1680 3785 1740
rect 3845 1680 3855 1740
rect 3775 1630 3855 1680
rect 3775 1570 3785 1630
rect 3845 1570 3855 1630
rect 3775 1565 3855 1570
rect 4175 1740 4255 1745
rect 4175 1680 4185 1740
rect 4245 1680 4255 1740
rect 4175 1630 4255 1680
rect 4175 1570 4185 1630
rect 4245 1570 4255 1630
rect 4175 1565 4255 1570
rect 4575 1740 4655 1745
rect 4575 1680 4585 1740
rect 4645 1680 4655 1740
rect 4575 1630 4655 1680
rect 4575 1570 4585 1630
rect 4645 1570 4655 1630
rect 4575 1565 4655 1570
rect 4975 1740 5055 1745
rect 4975 1680 4985 1740
rect 5045 1680 5055 1740
rect 4975 1630 5055 1680
rect 4975 1570 4985 1630
rect 5045 1570 5055 1630
rect 4975 1565 5055 1570
rect 5375 1740 5455 1745
rect 5375 1680 5385 1740
rect 5445 1680 5455 1740
rect 5375 1630 5455 1680
rect 5375 1570 5385 1630
rect 5445 1570 5455 1630
rect 5375 1565 5455 1570
rect 5775 1740 5855 1745
rect 5775 1680 5785 1740
rect 5845 1680 5855 1740
rect 5775 1630 5855 1680
rect 5775 1570 5785 1630
rect 5845 1570 5855 1630
rect 5775 1565 5855 1570
rect 6175 1740 6255 1745
rect 6175 1680 6185 1740
rect 6245 1680 6255 1740
rect 6175 1630 6255 1680
rect 6175 1570 6185 1630
rect 6245 1570 6255 1630
rect 6175 1565 6255 1570
rect 6575 1740 6655 1745
rect 6575 1680 6585 1740
rect 6645 1680 6655 1740
rect 6575 1630 6655 1680
rect 6575 1570 6585 1630
rect 6645 1570 6655 1630
rect 6575 1565 6655 1570
rect 6975 1740 7055 1745
rect 6975 1680 6985 1740
rect 7045 1680 7055 1740
rect 6975 1630 7055 1680
rect 6975 1570 6985 1630
rect 7045 1570 7055 1630
rect 6975 1565 7055 1570
rect 7375 1740 7455 1745
rect 7375 1680 7385 1740
rect 7445 1680 7455 1740
rect 7375 1630 7455 1680
rect 7375 1570 7385 1630
rect 7445 1570 7455 1630
rect 7375 1565 7455 1570
rect 7775 1740 7855 1745
rect 7775 1680 7785 1740
rect 7845 1680 7855 1740
rect 7775 1630 7855 1680
rect 7775 1570 7785 1630
rect 7845 1570 7855 1630
rect 7775 1565 7855 1570
rect 8175 1740 8255 1745
rect 8175 1680 8185 1740
rect 8245 1680 8255 1740
rect 8175 1630 8255 1680
rect 8175 1570 8185 1630
rect 8245 1570 8255 1630
rect 8175 1565 8255 1570
rect 8575 1740 8655 1745
rect 8575 1680 8585 1740
rect 8645 1680 8655 1740
rect 8575 1630 8655 1680
rect 8575 1570 8585 1630
rect 8645 1570 8655 1630
rect 8575 1565 8655 1570
rect 8975 1740 9055 1745
rect 8975 1680 8985 1740
rect 9045 1680 9055 1740
rect 8975 1630 9055 1680
rect 8975 1570 8985 1630
rect 9045 1570 9055 1630
rect 8975 1565 9055 1570
rect 9375 1740 9455 1745
rect 9375 1680 9385 1740
rect 9445 1680 9455 1740
rect 9375 1630 9455 1680
rect 9375 1570 9385 1630
rect 9445 1570 9455 1630
rect 9375 1565 9455 1570
rect 9775 1740 9855 1745
rect 9775 1680 9785 1740
rect 9845 1680 9855 1740
rect 9775 1630 9855 1680
rect 9775 1570 9785 1630
rect 9845 1570 9855 1630
rect 9775 1565 9855 1570
rect 10175 1740 10255 1745
rect 10175 1680 10185 1740
rect 10245 1680 10255 1740
rect 10175 1630 10255 1680
rect 10175 1570 10185 1630
rect 10245 1570 10255 1630
rect 10175 1565 10255 1570
rect 10575 1740 10655 1745
rect 10575 1680 10585 1740
rect 10645 1680 10655 1740
rect 10575 1630 10655 1680
rect 10575 1570 10585 1630
rect 10645 1570 10655 1630
rect 10575 1565 10655 1570
rect 10975 1740 11055 1745
rect 10975 1680 10985 1740
rect 11045 1680 11055 1740
rect 10975 1630 11055 1680
rect 10975 1570 10985 1630
rect 11045 1570 11055 1630
rect 10975 1565 11055 1570
rect 11375 1740 11455 1745
rect 11375 1680 11385 1740
rect 11445 1680 11455 1740
rect 11375 1630 11455 1680
rect 11375 1570 11385 1630
rect 11445 1570 11455 1630
rect 11375 1565 11455 1570
rect 11775 1740 11855 1745
rect 11775 1680 11785 1740
rect 11845 1680 11855 1740
rect 11775 1630 11855 1680
rect 11775 1570 11785 1630
rect 11845 1570 11855 1630
rect 11775 1565 11855 1570
rect 12175 1740 12255 1745
rect 12175 1680 12185 1740
rect 12245 1680 12255 1740
rect 12175 1630 12255 1680
rect 12175 1570 12185 1630
rect 12245 1570 12255 1630
rect 12175 1565 12255 1570
rect 12575 1740 12655 1745
rect 12575 1680 12585 1740
rect 12645 1680 12655 1740
rect 12575 1630 12655 1680
rect 12575 1570 12585 1630
rect 12645 1570 12655 1630
rect 12575 1565 12655 1570
rect 12975 1740 13055 1745
rect 12975 1680 12985 1740
rect 13045 1680 13055 1740
rect 12975 1630 13055 1680
rect 12975 1570 12985 1630
rect 13045 1570 13055 1630
rect 12975 1565 13055 1570
rect -215 1375 -155 1565
rect 185 1375 245 1565
rect 585 1375 645 1565
rect 985 1375 1045 1565
rect 1385 1375 1445 1565
rect 1785 1375 1845 1565
rect 2185 1375 2245 1565
rect 2585 1375 2645 1565
rect 2985 1375 3045 1565
rect 3385 1375 3445 1565
rect 3785 1375 3845 1565
rect 4185 1375 4245 1565
rect 4585 1375 4645 1565
rect 4985 1375 5045 1565
rect 5385 1375 5445 1565
rect 5785 1375 5845 1565
rect 6185 1375 6245 1565
rect 6585 1375 6645 1565
rect 6985 1375 7045 1565
rect 7385 1375 7445 1565
rect 7785 1375 7845 1565
rect 8185 1375 8245 1565
rect 8585 1375 8645 1565
rect 8985 1375 9045 1565
rect 9385 1375 9445 1565
rect 9785 1375 9845 1565
rect 10185 1375 10245 1565
rect 10585 1375 10645 1565
rect 10985 1375 11045 1565
rect 11385 1375 11445 1565
rect 11785 1375 11845 1565
rect 12185 1375 12245 1565
rect 12585 1375 12645 1565
rect 12985 1375 13045 1565
rect -225 1370 -145 1375
rect -225 1310 -215 1370
rect -155 1310 -145 1370
rect -225 1260 -145 1310
rect -225 1200 -215 1260
rect -155 1200 -145 1260
rect -225 1195 -145 1200
rect 175 1370 255 1375
rect 175 1310 185 1370
rect 245 1310 255 1370
rect 175 1260 255 1310
rect 175 1200 185 1260
rect 245 1200 255 1260
rect 175 1195 255 1200
rect 575 1370 655 1375
rect 575 1310 585 1370
rect 645 1310 655 1370
rect 575 1260 655 1310
rect 575 1200 585 1260
rect 645 1200 655 1260
rect 575 1195 655 1200
rect 975 1370 1055 1375
rect 975 1310 985 1370
rect 1045 1310 1055 1370
rect 975 1260 1055 1310
rect 975 1200 985 1260
rect 1045 1200 1055 1260
rect 975 1195 1055 1200
rect 1375 1370 1455 1375
rect 1375 1310 1385 1370
rect 1445 1310 1455 1370
rect 1375 1260 1455 1310
rect 1375 1200 1385 1260
rect 1445 1200 1455 1260
rect 1375 1195 1455 1200
rect 1775 1370 1855 1375
rect 1775 1310 1785 1370
rect 1845 1310 1855 1370
rect 1775 1260 1855 1310
rect 1775 1200 1785 1260
rect 1845 1200 1855 1260
rect 1775 1195 1855 1200
rect 2175 1370 2255 1375
rect 2175 1310 2185 1370
rect 2245 1310 2255 1370
rect 2175 1260 2255 1310
rect 2175 1200 2185 1260
rect 2245 1200 2255 1260
rect 2175 1195 2255 1200
rect 2575 1370 2655 1375
rect 2575 1310 2585 1370
rect 2645 1310 2655 1370
rect 2575 1260 2655 1310
rect 2575 1200 2585 1260
rect 2645 1200 2655 1260
rect 2575 1195 2655 1200
rect 2975 1370 3055 1375
rect 2975 1310 2985 1370
rect 3045 1310 3055 1370
rect 2975 1260 3055 1310
rect 2975 1200 2985 1260
rect 3045 1200 3055 1260
rect 2975 1195 3055 1200
rect 3375 1370 3455 1375
rect 3375 1310 3385 1370
rect 3445 1310 3455 1370
rect 3375 1260 3455 1310
rect 3375 1200 3385 1260
rect 3445 1200 3455 1260
rect 3375 1195 3455 1200
rect 3775 1370 3855 1375
rect 3775 1310 3785 1370
rect 3845 1310 3855 1370
rect 3775 1260 3855 1310
rect 3775 1200 3785 1260
rect 3845 1200 3855 1260
rect 3775 1195 3855 1200
rect 4175 1370 4255 1375
rect 4175 1310 4185 1370
rect 4245 1310 4255 1370
rect 4175 1260 4255 1310
rect 4175 1200 4185 1260
rect 4245 1200 4255 1260
rect 4175 1195 4255 1200
rect 4575 1370 4655 1375
rect 4575 1310 4585 1370
rect 4645 1310 4655 1370
rect 4575 1260 4655 1310
rect 4575 1200 4585 1260
rect 4645 1200 4655 1260
rect 4575 1195 4655 1200
rect 4975 1370 5055 1375
rect 4975 1310 4985 1370
rect 5045 1310 5055 1370
rect 4975 1260 5055 1310
rect 4975 1200 4985 1260
rect 5045 1200 5055 1260
rect 4975 1195 5055 1200
rect 5375 1370 5455 1375
rect 5375 1310 5385 1370
rect 5445 1310 5455 1370
rect 5375 1260 5455 1310
rect 5375 1200 5385 1260
rect 5445 1200 5455 1260
rect 5375 1195 5455 1200
rect 5775 1370 5855 1375
rect 5775 1310 5785 1370
rect 5845 1310 5855 1370
rect 5775 1260 5855 1310
rect 5775 1200 5785 1260
rect 5845 1200 5855 1260
rect 5775 1195 5855 1200
rect 6175 1370 6255 1375
rect 6175 1310 6185 1370
rect 6245 1310 6255 1370
rect 6175 1260 6255 1310
rect 6175 1200 6185 1260
rect 6245 1200 6255 1260
rect 6175 1195 6255 1200
rect 6575 1370 6655 1375
rect 6575 1310 6585 1370
rect 6645 1310 6655 1370
rect 6575 1260 6655 1310
rect 6575 1200 6585 1260
rect 6645 1200 6655 1260
rect 6575 1195 6655 1200
rect 6975 1370 7055 1375
rect 6975 1310 6985 1370
rect 7045 1310 7055 1370
rect 6975 1260 7055 1310
rect 6975 1200 6985 1260
rect 7045 1200 7055 1260
rect 6975 1195 7055 1200
rect 7375 1370 7455 1375
rect 7375 1310 7385 1370
rect 7445 1310 7455 1370
rect 7375 1260 7455 1310
rect 7375 1200 7385 1260
rect 7445 1200 7455 1260
rect 7375 1195 7455 1200
rect 7775 1370 7855 1375
rect 7775 1310 7785 1370
rect 7845 1310 7855 1370
rect 7775 1260 7855 1310
rect 7775 1200 7785 1260
rect 7845 1200 7855 1260
rect 7775 1195 7855 1200
rect 8175 1370 8255 1375
rect 8175 1310 8185 1370
rect 8245 1310 8255 1370
rect 8175 1260 8255 1310
rect 8175 1200 8185 1260
rect 8245 1200 8255 1260
rect 8175 1195 8255 1200
rect 8575 1370 8655 1375
rect 8575 1310 8585 1370
rect 8645 1310 8655 1370
rect 8575 1260 8655 1310
rect 8575 1200 8585 1260
rect 8645 1200 8655 1260
rect 8575 1195 8655 1200
rect 8975 1370 9055 1375
rect 8975 1310 8985 1370
rect 9045 1310 9055 1370
rect 8975 1260 9055 1310
rect 8975 1200 8985 1260
rect 9045 1200 9055 1260
rect 8975 1195 9055 1200
rect 9375 1370 9455 1375
rect 9375 1310 9385 1370
rect 9445 1310 9455 1370
rect 9375 1260 9455 1310
rect 9375 1200 9385 1260
rect 9445 1200 9455 1260
rect 9375 1195 9455 1200
rect 9775 1370 9855 1375
rect 9775 1310 9785 1370
rect 9845 1310 9855 1370
rect 9775 1260 9855 1310
rect 9775 1200 9785 1260
rect 9845 1200 9855 1260
rect 9775 1195 9855 1200
rect 10175 1370 10255 1375
rect 10175 1310 10185 1370
rect 10245 1310 10255 1370
rect 10175 1260 10255 1310
rect 10175 1200 10185 1260
rect 10245 1200 10255 1260
rect 10175 1195 10255 1200
rect 10575 1370 10655 1375
rect 10575 1310 10585 1370
rect 10645 1310 10655 1370
rect 10575 1260 10655 1310
rect 10575 1200 10585 1260
rect 10645 1200 10655 1260
rect 10575 1195 10655 1200
rect 10975 1370 11055 1375
rect 10975 1310 10985 1370
rect 11045 1310 11055 1370
rect 10975 1260 11055 1310
rect 10975 1200 10985 1260
rect 11045 1200 11055 1260
rect 10975 1195 11055 1200
rect 11375 1370 11455 1375
rect 11375 1310 11385 1370
rect 11445 1310 11455 1370
rect 11375 1260 11455 1310
rect 11375 1200 11385 1260
rect 11445 1200 11455 1260
rect 11375 1195 11455 1200
rect 11775 1370 11855 1375
rect 11775 1310 11785 1370
rect 11845 1310 11855 1370
rect 11775 1260 11855 1310
rect 11775 1200 11785 1260
rect 11845 1200 11855 1260
rect 11775 1195 11855 1200
rect 12175 1370 12255 1375
rect 12175 1310 12185 1370
rect 12245 1310 12255 1370
rect 12175 1260 12255 1310
rect 12175 1200 12185 1260
rect 12245 1200 12255 1260
rect 12175 1195 12255 1200
rect 12575 1370 12655 1375
rect 12575 1310 12585 1370
rect 12645 1310 12655 1370
rect 12575 1260 12655 1310
rect 12575 1200 12585 1260
rect 12645 1200 12655 1260
rect 12575 1195 12655 1200
rect 12975 1370 13055 1375
rect 12975 1310 12985 1370
rect 13045 1310 13055 1370
rect 12975 1260 13055 1310
rect 12975 1200 12985 1260
rect 13045 1200 13055 1260
rect 12975 1195 13055 1200
rect -215 1005 -155 1195
rect 185 1005 245 1195
rect 585 1005 645 1195
rect 985 1005 1045 1195
rect 1385 1005 1445 1195
rect 1785 1005 1845 1195
rect 2185 1005 2245 1195
rect 2585 1005 2645 1195
rect 2985 1005 3045 1195
rect 3385 1005 3445 1195
rect 3785 1005 3845 1195
rect 4185 1005 4245 1195
rect 4585 1005 4645 1195
rect 4985 1005 5045 1195
rect 5385 1005 5445 1195
rect 5785 1005 5845 1195
rect 6185 1005 6245 1195
rect 6585 1005 6645 1195
rect 6985 1005 7045 1195
rect 7385 1005 7445 1195
rect 7785 1005 7845 1195
rect 8185 1005 8245 1195
rect 8585 1005 8645 1195
rect 8985 1005 9045 1195
rect 9385 1005 9445 1195
rect 9785 1005 9845 1195
rect 10185 1005 10245 1195
rect 10585 1005 10645 1195
rect 10985 1005 11045 1195
rect 11385 1005 11445 1195
rect 11785 1005 11845 1195
rect 12185 1005 12245 1195
rect 12585 1005 12645 1195
rect 12985 1005 13045 1195
rect -225 1000 -145 1005
rect -225 940 -215 1000
rect -155 940 -145 1000
rect -225 890 -145 940
rect -225 830 -215 890
rect -155 830 -145 890
rect -225 825 -145 830
rect 175 1000 255 1005
rect 175 940 185 1000
rect 245 940 255 1000
rect 175 890 255 940
rect 175 830 185 890
rect 245 830 255 890
rect 175 825 255 830
rect 575 1000 655 1005
rect 575 940 585 1000
rect 645 940 655 1000
rect 575 890 655 940
rect 575 830 585 890
rect 645 830 655 890
rect 575 825 655 830
rect 975 1000 1055 1005
rect 975 940 985 1000
rect 1045 940 1055 1000
rect 975 890 1055 940
rect 975 830 985 890
rect 1045 830 1055 890
rect 975 825 1055 830
rect 1375 1000 1455 1005
rect 1375 940 1385 1000
rect 1445 940 1455 1000
rect 1375 890 1455 940
rect 1375 830 1385 890
rect 1445 830 1455 890
rect 1375 825 1455 830
rect 1775 1000 1855 1005
rect 1775 940 1785 1000
rect 1845 940 1855 1000
rect 1775 890 1855 940
rect 1775 830 1785 890
rect 1845 830 1855 890
rect 1775 825 1855 830
rect 2175 1000 2255 1005
rect 2175 940 2185 1000
rect 2245 940 2255 1000
rect 2175 890 2255 940
rect 2175 830 2185 890
rect 2245 830 2255 890
rect 2175 825 2255 830
rect 2575 1000 2655 1005
rect 2575 940 2585 1000
rect 2645 940 2655 1000
rect 2575 890 2655 940
rect 2575 830 2585 890
rect 2645 830 2655 890
rect 2575 825 2655 830
rect 2975 1000 3055 1005
rect 2975 940 2985 1000
rect 3045 940 3055 1000
rect 2975 890 3055 940
rect 2975 830 2985 890
rect 3045 830 3055 890
rect 2975 825 3055 830
rect 3375 1000 3455 1005
rect 3375 940 3385 1000
rect 3445 940 3455 1000
rect 3375 890 3455 940
rect 3375 830 3385 890
rect 3445 830 3455 890
rect 3375 825 3455 830
rect 3775 1000 3855 1005
rect 3775 940 3785 1000
rect 3845 940 3855 1000
rect 3775 890 3855 940
rect 3775 830 3785 890
rect 3845 830 3855 890
rect 3775 825 3855 830
rect 4175 1000 4255 1005
rect 4175 940 4185 1000
rect 4245 940 4255 1000
rect 4175 890 4255 940
rect 4175 830 4185 890
rect 4245 830 4255 890
rect 4175 825 4255 830
rect 4575 1000 4655 1005
rect 4575 940 4585 1000
rect 4645 940 4655 1000
rect 4575 890 4655 940
rect 4575 830 4585 890
rect 4645 830 4655 890
rect 4575 825 4655 830
rect 4975 1000 5055 1005
rect 4975 940 4985 1000
rect 5045 940 5055 1000
rect 4975 890 5055 940
rect 4975 830 4985 890
rect 5045 830 5055 890
rect 4975 825 5055 830
rect 5375 1000 5455 1005
rect 5375 940 5385 1000
rect 5445 940 5455 1000
rect 5375 890 5455 940
rect 5375 830 5385 890
rect 5445 830 5455 890
rect 5375 825 5455 830
rect 5775 1000 5855 1005
rect 5775 940 5785 1000
rect 5845 940 5855 1000
rect 5775 890 5855 940
rect 5775 830 5785 890
rect 5845 830 5855 890
rect 5775 825 5855 830
rect 6175 1000 6255 1005
rect 6175 940 6185 1000
rect 6245 940 6255 1000
rect 6175 890 6255 940
rect 6175 830 6185 890
rect 6245 830 6255 890
rect 6175 825 6255 830
rect 6575 1000 6655 1005
rect 6575 940 6585 1000
rect 6645 940 6655 1000
rect 6575 890 6655 940
rect 6575 830 6585 890
rect 6645 830 6655 890
rect 6575 825 6655 830
rect 6975 1000 7055 1005
rect 6975 940 6985 1000
rect 7045 940 7055 1000
rect 6975 890 7055 940
rect 6975 830 6985 890
rect 7045 830 7055 890
rect 6975 825 7055 830
rect 7375 1000 7455 1005
rect 7375 940 7385 1000
rect 7445 940 7455 1000
rect 7375 890 7455 940
rect 7375 830 7385 890
rect 7445 830 7455 890
rect 7375 825 7455 830
rect 7775 1000 7855 1005
rect 7775 940 7785 1000
rect 7845 940 7855 1000
rect 7775 890 7855 940
rect 7775 830 7785 890
rect 7845 830 7855 890
rect 7775 825 7855 830
rect 8175 1000 8255 1005
rect 8175 940 8185 1000
rect 8245 940 8255 1000
rect 8175 890 8255 940
rect 8175 830 8185 890
rect 8245 830 8255 890
rect 8175 825 8255 830
rect 8575 1000 8655 1005
rect 8575 940 8585 1000
rect 8645 940 8655 1000
rect 8575 890 8655 940
rect 8575 830 8585 890
rect 8645 830 8655 890
rect 8575 825 8655 830
rect 8975 1000 9055 1005
rect 8975 940 8985 1000
rect 9045 940 9055 1000
rect 8975 890 9055 940
rect 8975 830 8985 890
rect 9045 830 9055 890
rect 8975 825 9055 830
rect 9375 1000 9455 1005
rect 9375 940 9385 1000
rect 9445 940 9455 1000
rect 9375 890 9455 940
rect 9375 830 9385 890
rect 9445 830 9455 890
rect 9375 825 9455 830
rect 9775 1000 9855 1005
rect 9775 940 9785 1000
rect 9845 940 9855 1000
rect 9775 890 9855 940
rect 9775 830 9785 890
rect 9845 830 9855 890
rect 9775 825 9855 830
rect 10175 1000 10255 1005
rect 10175 940 10185 1000
rect 10245 940 10255 1000
rect 10175 890 10255 940
rect 10175 830 10185 890
rect 10245 830 10255 890
rect 10175 825 10255 830
rect 10575 1000 10655 1005
rect 10575 940 10585 1000
rect 10645 940 10655 1000
rect 10575 890 10655 940
rect 10575 830 10585 890
rect 10645 830 10655 890
rect 10575 825 10655 830
rect 10975 1000 11055 1005
rect 10975 940 10985 1000
rect 11045 940 11055 1000
rect 10975 890 11055 940
rect 10975 830 10985 890
rect 11045 830 11055 890
rect 10975 825 11055 830
rect 11375 1000 11455 1005
rect 11375 940 11385 1000
rect 11445 940 11455 1000
rect 11375 890 11455 940
rect 11375 830 11385 890
rect 11445 830 11455 890
rect 11375 825 11455 830
rect 11775 1000 11855 1005
rect 11775 940 11785 1000
rect 11845 940 11855 1000
rect 11775 890 11855 940
rect 11775 830 11785 890
rect 11845 830 11855 890
rect 11775 825 11855 830
rect 12175 1000 12255 1005
rect 12175 940 12185 1000
rect 12245 940 12255 1000
rect 12175 890 12255 940
rect 12175 830 12185 890
rect 12245 830 12255 890
rect 12175 825 12255 830
rect 12575 1000 12655 1005
rect 12575 940 12585 1000
rect 12645 940 12655 1000
rect 12575 890 12655 940
rect 12575 830 12585 890
rect 12645 830 12655 890
rect 12575 825 12655 830
rect 12975 1000 13055 1005
rect 12975 940 12985 1000
rect 13045 940 13055 1000
rect 12975 890 13055 940
rect 12975 830 12985 890
rect 13045 830 13055 890
rect 12975 825 13055 830
rect -215 635 -155 825
rect 185 635 245 825
rect 585 635 645 825
rect 985 635 1045 825
rect 1385 635 1445 825
rect 1785 635 1845 825
rect 2185 635 2245 825
rect 2585 635 2645 825
rect 2985 635 3045 825
rect 3385 635 3445 825
rect 3785 635 3845 825
rect 4185 635 4245 825
rect 4585 635 4645 825
rect 4985 635 5045 825
rect 5385 635 5445 825
rect 5785 635 5845 825
rect 6185 635 6245 825
rect 6585 635 6645 825
rect 6985 635 7045 825
rect 7385 635 7445 825
rect 7785 635 7845 825
rect 8185 635 8245 825
rect 8585 635 8645 825
rect 8985 635 9045 825
rect 9385 635 9445 825
rect 9785 635 9845 825
rect 10185 635 10245 825
rect 10585 635 10645 825
rect 10985 635 11045 825
rect 11385 635 11445 825
rect 11785 635 11845 825
rect 12185 635 12245 825
rect 12585 635 12645 825
rect 12985 635 13045 825
rect -225 630 -145 635
rect -225 570 -215 630
rect -155 570 -145 630
rect -225 520 -145 570
rect -225 460 -215 520
rect -155 460 -145 520
rect -225 455 -145 460
rect 175 630 255 635
rect 175 570 185 630
rect 245 570 255 630
rect 175 520 255 570
rect 175 460 185 520
rect 245 460 255 520
rect 175 455 255 460
rect 575 630 655 635
rect 575 570 585 630
rect 645 570 655 630
rect 575 520 655 570
rect 575 460 585 520
rect 645 460 655 520
rect 575 455 655 460
rect 975 630 1055 635
rect 975 570 985 630
rect 1045 570 1055 630
rect 975 520 1055 570
rect 975 460 985 520
rect 1045 460 1055 520
rect 975 455 1055 460
rect 1375 630 1455 635
rect 1375 570 1385 630
rect 1445 570 1455 630
rect 1375 520 1455 570
rect 1375 460 1385 520
rect 1445 460 1455 520
rect 1375 455 1455 460
rect 1775 630 1855 635
rect 1775 570 1785 630
rect 1845 570 1855 630
rect 1775 520 1855 570
rect 1775 460 1785 520
rect 1845 460 1855 520
rect 1775 455 1855 460
rect 2175 630 2255 635
rect 2175 570 2185 630
rect 2245 570 2255 630
rect 2175 520 2255 570
rect 2175 460 2185 520
rect 2245 460 2255 520
rect 2175 455 2255 460
rect 2575 630 2655 635
rect 2575 570 2585 630
rect 2645 570 2655 630
rect 2575 520 2655 570
rect 2575 460 2585 520
rect 2645 460 2655 520
rect 2575 455 2655 460
rect 2975 630 3055 635
rect 2975 570 2985 630
rect 3045 570 3055 630
rect 2975 520 3055 570
rect 2975 460 2985 520
rect 3045 460 3055 520
rect 2975 455 3055 460
rect 3375 630 3455 635
rect 3375 570 3385 630
rect 3445 570 3455 630
rect 3375 520 3455 570
rect 3375 460 3385 520
rect 3445 460 3455 520
rect 3375 455 3455 460
rect 3775 630 3855 635
rect 3775 570 3785 630
rect 3845 570 3855 630
rect 3775 520 3855 570
rect 3775 460 3785 520
rect 3845 460 3855 520
rect 3775 455 3855 460
rect 4175 630 4255 635
rect 4175 570 4185 630
rect 4245 570 4255 630
rect 4175 520 4255 570
rect 4175 460 4185 520
rect 4245 460 4255 520
rect 4175 455 4255 460
rect 4575 630 4655 635
rect 4575 570 4585 630
rect 4645 570 4655 630
rect 4575 520 4655 570
rect 4575 460 4585 520
rect 4645 460 4655 520
rect 4575 455 4655 460
rect 4975 630 5055 635
rect 4975 570 4985 630
rect 5045 570 5055 630
rect 4975 520 5055 570
rect 4975 460 4985 520
rect 5045 460 5055 520
rect 4975 455 5055 460
rect 5375 630 5455 635
rect 5375 570 5385 630
rect 5445 570 5455 630
rect 5375 520 5455 570
rect 5375 460 5385 520
rect 5445 460 5455 520
rect 5375 455 5455 460
rect 5775 630 5855 635
rect 5775 570 5785 630
rect 5845 570 5855 630
rect 5775 520 5855 570
rect 5775 460 5785 520
rect 5845 460 5855 520
rect 5775 455 5855 460
rect 6175 630 6255 635
rect 6175 570 6185 630
rect 6245 570 6255 630
rect 6175 520 6255 570
rect 6175 460 6185 520
rect 6245 460 6255 520
rect 6175 455 6255 460
rect 6575 630 6655 635
rect 6575 570 6585 630
rect 6645 570 6655 630
rect 6575 520 6655 570
rect 6575 460 6585 520
rect 6645 460 6655 520
rect 6575 455 6655 460
rect 6975 630 7055 635
rect 6975 570 6985 630
rect 7045 570 7055 630
rect 6975 520 7055 570
rect 6975 460 6985 520
rect 7045 460 7055 520
rect 6975 455 7055 460
rect 7375 630 7455 635
rect 7375 570 7385 630
rect 7445 570 7455 630
rect 7375 520 7455 570
rect 7375 460 7385 520
rect 7445 460 7455 520
rect 7375 455 7455 460
rect 7775 630 7855 635
rect 7775 570 7785 630
rect 7845 570 7855 630
rect 7775 520 7855 570
rect 7775 460 7785 520
rect 7845 460 7855 520
rect 7775 455 7855 460
rect 8175 630 8255 635
rect 8175 570 8185 630
rect 8245 570 8255 630
rect 8175 520 8255 570
rect 8175 460 8185 520
rect 8245 460 8255 520
rect 8175 455 8255 460
rect 8575 630 8655 635
rect 8575 570 8585 630
rect 8645 570 8655 630
rect 8575 520 8655 570
rect 8575 460 8585 520
rect 8645 460 8655 520
rect 8575 455 8655 460
rect 8975 630 9055 635
rect 8975 570 8985 630
rect 9045 570 9055 630
rect 8975 520 9055 570
rect 8975 460 8985 520
rect 9045 460 9055 520
rect 8975 455 9055 460
rect 9375 630 9455 635
rect 9375 570 9385 630
rect 9445 570 9455 630
rect 9375 520 9455 570
rect 9375 460 9385 520
rect 9445 460 9455 520
rect 9375 455 9455 460
rect 9775 630 9855 635
rect 9775 570 9785 630
rect 9845 570 9855 630
rect 9775 520 9855 570
rect 9775 460 9785 520
rect 9845 460 9855 520
rect 9775 455 9855 460
rect 10175 630 10255 635
rect 10175 570 10185 630
rect 10245 570 10255 630
rect 10175 520 10255 570
rect 10175 460 10185 520
rect 10245 460 10255 520
rect 10175 455 10255 460
rect 10575 630 10655 635
rect 10575 570 10585 630
rect 10645 570 10655 630
rect 10575 520 10655 570
rect 10575 460 10585 520
rect 10645 460 10655 520
rect 10575 455 10655 460
rect 10975 630 11055 635
rect 10975 570 10985 630
rect 11045 570 11055 630
rect 10975 520 11055 570
rect 10975 460 10985 520
rect 11045 460 11055 520
rect 10975 455 11055 460
rect 11375 630 11455 635
rect 11375 570 11385 630
rect 11445 570 11455 630
rect 11375 520 11455 570
rect 11375 460 11385 520
rect 11445 460 11455 520
rect 11375 455 11455 460
rect 11775 630 11855 635
rect 11775 570 11785 630
rect 11845 570 11855 630
rect 11775 520 11855 570
rect 11775 460 11785 520
rect 11845 460 11855 520
rect 11775 455 11855 460
rect 12175 630 12255 635
rect 12175 570 12185 630
rect 12245 570 12255 630
rect 12175 520 12255 570
rect 12175 460 12185 520
rect 12245 460 12255 520
rect 12175 455 12255 460
rect 12575 630 12655 635
rect 12575 570 12585 630
rect 12645 570 12655 630
rect 12575 520 12655 570
rect 12575 460 12585 520
rect 12645 460 12655 520
rect 12575 455 12655 460
rect 12975 630 13055 635
rect 12975 570 12985 630
rect 13045 570 13055 630
rect 12975 520 13055 570
rect 12975 460 12985 520
rect 13045 460 13055 520
rect 12975 455 13055 460
rect -215 265 -155 455
rect 185 265 245 455
rect 585 265 645 455
rect 985 265 1045 455
rect 1385 265 1445 455
rect 1785 265 1845 455
rect 2185 265 2245 455
rect 2585 265 2645 455
rect 2985 265 3045 455
rect 3385 265 3445 455
rect 3785 265 3845 455
rect 4185 265 4245 455
rect 4585 265 4645 455
rect 4985 265 5045 455
rect 5385 265 5445 455
rect 5785 265 5845 455
rect 6185 265 6245 455
rect 6585 265 6645 455
rect 6985 265 7045 455
rect 7385 265 7445 455
rect 7785 265 7845 455
rect 8185 265 8245 455
rect 8585 265 8645 455
rect 8985 265 9045 455
rect 9385 265 9445 455
rect 9785 265 9845 455
rect 10185 265 10245 455
rect 10585 265 10645 455
rect 10985 265 11045 455
rect 11385 265 11445 455
rect 11785 265 11845 455
rect 12185 265 12245 455
rect 12585 265 12645 455
rect 12985 265 13045 455
rect -225 260 -145 265
rect -225 200 -215 260
rect -155 200 -145 260
rect -225 150 -145 200
rect -225 90 -215 150
rect -155 90 -145 150
rect -225 85 -145 90
rect 175 260 255 265
rect 175 200 185 260
rect 245 200 255 260
rect 175 150 255 200
rect 175 90 185 150
rect 245 90 255 150
rect 175 85 255 90
rect 575 260 655 265
rect 575 200 585 260
rect 645 200 655 260
rect 575 150 655 200
rect 575 90 585 150
rect 645 90 655 150
rect 575 85 655 90
rect 975 260 1055 265
rect 975 200 985 260
rect 1045 200 1055 260
rect 975 150 1055 200
rect 975 90 985 150
rect 1045 90 1055 150
rect 975 85 1055 90
rect 1375 260 1455 265
rect 1375 200 1385 260
rect 1445 200 1455 260
rect 1375 150 1455 200
rect 1375 90 1385 150
rect 1445 90 1455 150
rect 1375 85 1455 90
rect 1775 260 1855 265
rect 1775 200 1785 260
rect 1845 200 1855 260
rect 1775 150 1855 200
rect 1775 90 1785 150
rect 1845 90 1855 150
rect 1775 85 1855 90
rect 2175 260 2255 265
rect 2175 200 2185 260
rect 2245 200 2255 260
rect 2175 150 2255 200
rect 2175 90 2185 150
rect 2245 90 2255 150
rect 2175 85 2255 90
rect 2575 260 2655 265
rect 2575 200 2585 260
rect 2645 200 2655 260
rect 2575 150 2655 200
rect 2575 90 2585 150
rect 2645 90 2655 150
rect 2575 85 2655 90
rect 2975 260 3055 265
rect 2975 200 2985 260
rect 3045 200 3055 260
rect 2975 150 3055 200
rect 2975 90 2985 150
rect 3045 90 3055 150
rect 2975 85 3055 90
rect 3375 260 3455 265
rect 3375 200 3385 260
rect 3445 200 3455 260
rect 3375 150 3455 200
rect 3375 90 3385 150
rect 3445 90 3455 150
rect 3375 85 3455 90
rect 3775 260 3855 265
rect 3775 200 3785 260
rect 3845 200 3855 260
rect 3775 150 3855 200
rect 3775 90 3785 150
rect 3845 90 3855 150
rect 3775 85 3855 90
rect 4175 260 4255 265
rect 4175 200 4185 260
rect 4245 200 4255 260
rect 4175 150 4255 200
rect 4175 90 4185 150
rect 4245 90 4255 150
rect 4175 85 4255 90
rect 4575 260 4655 265
rect 4575 200 4585 260
rect 4645 200 4655 260
rect 4575 150 4655 200
rect 4575 90 4585 150
rect 4645 90 4655 150
rect 4575 85 4655 90
rect 4975 260 5055 265
rect 4975 200 4985 260
rect 5045 200 5055 260
rect 4975 150 5055 200
rect 4975 90 4985 150
rect 5045 90 5055 150
rect 4975 85 5055 90
rect 5375 260 5455 265
rect 5375 200 5385 260
rect 5445 200 5455 260
rect 5375 150 5455 200
rect 5375 90 5385 150
rect 5445 90 5455 150
rect 5375 85 5455 90
rect 5775 260 5855 265
rect 5775 200 5785 260
rect 5845 200 5855 260
rect 5775 150 5855 200
rect 5775 90 5785 150
rect 5845 90 5855 150
rect 5775 85 5855 90
rect 6175 260 6255 265
rect 6175 200 6185 260
rect 6245 200 6255 260
rect 6175 150 6255 200
rect 6175 90 6185 150
rect 6245 90 6255 150
rect 6175 85 6255 90
rect 6575 260 6655 265
rect 6575 200 6585 260
rect 6645 200 6655 260
rect 6575 150 6655 200
rect 6575 90 6585 150
rect 6645 90 6655 150
rect 6575 85 6655 90
rect 6975 260 7055 265
rect 6975 200 6985 260
rect 7045 200 7055 260
rect 6975 150 7055 200
rect 6975 90 6985 150
rect 7045 90 7055 150
rect 6975 85 7055 90
rect 7375 260 7455 265
rect 7375 200 7385 260
rect 7445 200 7455 260
rect 7375 150 7455 200
rect 7375 90 7385 150
rect 7445 90 7455 150
rect 7375 85 7455 90
rect 7775 260 7855 265
rect 7775 200 7785 260
rect 7845 200 7855 260
rect 7775 150 7855 200
rect 7775 90 7785 150
rect 7845 90 7855 150
rect 7775 85 7855 90
rect 8175 260 8255 265
rect 8175 200 8185 260
rect 8245 200 8255 260
rect 8175 150 8255 200
rect 8175 90 8185 150
rect 8245 90 8255 150
rect 8175 85 8255 90
rect 8575 260 8655 265
rect 8575 200 8585 260
rect 8645 200 8655 260
rect 8575 150 8655 200
rect 8575 90 8585 150
rect 8645 90 8655 150
rect 8575 85 8655 90
rect 8975 260 9055 265
rect 8975 200 8985 260
rect 9045 200 9055 260
rect 8975 150 9055 200
rect 8975 90 8985 150
rect 9045 90 9055 150
rect 8975 85 9055 90
rect 9375 260 9455 265
rect 9375 200 9385 260
rect 9445 200 9455 260
rect 9375 150 9455 200
rect 9375 90 9385 150
rect 9445 90 9455 150
rect 9375 85 9455 90
rect 9775 260 9855 265
rect 9775 200 9785 260
rect 9845 200 9855 260
rect 9775 150 9855 200
rect 9775 90 9785 150
rect 9845 90 9855 150
rect 9775 85 9855 90
rect 10175 260 10255 265
rect 10175 200 10185 260
rect 10245 200 10255 260
rect 10175 150 10255 200
rect 10175 90 10185 150
rect 10245 90 10255 150
rect 10175 85 10255 90
rect 10575 260 10655 265
rect 10575 200 10585 260
rect 10645 200 10655 260
rect 10575 150 10655 200
rect 10575 90 10585 150
rect 10645 90 10655 150
rect 10575 85 10655 90
rect 10975 260 11055 265
rect 10975 200 10985 260
rect 11045 200 11055 260
rect 10975 150 11055 200
rect 10975 90 10985 150
rect 11045 90 11055 150
rect 10975 85 11055 90
rect 11375 260 11455 265
rect 11375 200 11385 260
rect 11445 200 11455 260
rect 11375 150 11455 200
rect 11375 90 11385 150
rect 11445 90 11455 150
rect 11375 85 11455 90
rect 11775 260 11855 265
rect 11775 200 11785 260
rect 11845 200 11855 260
rect 11775 150 11855 200
rect 11775 90 11785 150
rect 11845 90 11855 150
rect 11775 85 11855 90
rect 12175 260 12255 265
rect 12175 200 12185 260
rect 12245 200 12255 260
rect 12175 150 12255 200
rect 12175 90 12185 150
rect 12245 90 12255 150
rect 12175 85 12255 90
rect 12575 260 12655 265
rect 12575 200 12585 260
rect 12645 200 12655 260
rect 12575 150 12655 200
rect 12575 90 12585 150
rect 12645 90 12655 150
rect 12575 85 12655 90
rect 12975 260 13055 265
rect 12975 200 12985 260
rect 13045 200 13055 260
rect 12975 150 13055 200
rect 12975 90 12985 150
rect 13045 90 13055 150
rect 12975 85 13055 90
rect -215 -105 -155 85
rect 185 -105 245 85
rect 585 -105 645 85
rect 985 -105 1045 85
rect 1385 -105 1445 85
rect 1785 -105 1845 85
rect 2185 -105 2245 85
rect 2585 -105 2645 85
rect 2985 -105 3045 85
rect 3385 -105 3445 85
rect 3785 -105 3845 85
rect 4185 -105 4245 85
rect 4585 -105 4645 85
rect 4985 -105 5045 85
rect 5385 -105 5445 85
rect 5785 -105 5845 85
rect 6185 -105 6245 85
rect 6585 -105 6645 85
rect 6985 -105 7045 85
rect 7385 -105 7445 85
rect 7785 -105 7845 85
rect 8185 -105 8245 85
rect 8585 -105 8645 85
rect 8985 -105 9045 85
rect 9385 -105 9445 85
rect 9785 -105 9845 85
rect 10185 -105 10245 85
rect 10585 -105 10645 85
rect 10985 -105 11045 85
rect 11385 -105 11445 85
rect 11785 -105 11845 85
rect 12185 -105 12245 85
rect 12585 -105 12645 85
rect 12985 -105 13045 85
rect -225 -110 -145 -105
rect -225 -170 -215 -110
rect -155 -170 -145 -110
rect -225 -220 -145 -170
rect -225 -280 -215 -220
rect -155 -280 -145 -220
rect -225 -285 -145 -280
rect 175 -110 255 -105
rect 175 -170 185 -110
rect 245 -170 255 -110
rect 175 -220 255 -170
rect 175 -280 185 -220
rect 245 -280 255 -220
rect 175 -285 255 -280
rect 575 -110 655 -105
rect 575 -170 585 -110
rect 645 -170 655 -110
rect 575 -220 655 -170
rect 575 -280 585 -220
rect 645 -280 655 -220
rect 575 -285 655 -280
rect 975 -110 1055 -105
rect 975 -170 985 -110
rect 1045 -170 1055 -110
rect 975 -220 1055 -170
rect 975 -280 985 -220
rect 1045 -280 1055 -220
rect 975 -285 1055 -280
rect 1375 -110 1455 -105
rect 1375 -170 1385 -110
rect 1445 -170 1455 -110
rect 1375 -220 1455 -170
rect 1375 -280 1385 -220
rect 1445 -280 1455 -220
rect 1375 -285 1455 -280
rect 1775 -110 1855 -105
rect 1775 -170 1785 -110
rect 1845 -170 1855 -110
rect 1775 -220 1855 -170
rect 1775 -280 1785 -220
rect 1845 -280 1855 -220
rect 1775 -285 1855 -280
rect 2175 -110 2255 -105
rect 2175 -170 2185 -110
rect 2245 -170 2255 -110
rect 2175 -220 2255 -170
rect 2175 -280 2185 -220
rect 2245 -280 2255 -220
rect 2175 -285 2255 -280
rect 2575 -110 2655 -105
rect 2575 -170 2585 -110
rect 2645 -170 2655 -110
rect 2575 -220 2655 -170
rect 2575 -280 2585 -220
rect 2645 -280 2655 -220
rect 2575 -285 2655 -280
rect 2975 -110 3055 -105
rect 2975 -170 2985 -110
rect 3045 -170 3055 -110
rect 2975 -220 3055 -170
rect 2975 -280 2985 -220
rect 3045 -280 3055 -220
rect 2975 -285 3055 -280
rect 3375 -110 3455 -105
rect 3375 -170 3385 -110
rect 3445 -170 3455 -110
rect 3375 -220 3455 -170
rect 3375 -280 3385 -220
rect 3445 -280 3455 -220
rect 3375 -285 3455 -280
rect 3775 -110 3855 -105
rect 3775 -170 3785 -110
rect 3845 -170 3855 -110
rect 3775 -220 3855 -170
rect 3775 -280 3785 -220
rect 3845 -280 3855 -220
rect 3775 -285 3855 -280
rect 4175 -110 4255 -105
rect 4175 -170 4185 -110
rect 4245 -170 4255 -110
rect 4175 -220 4255 -170
rect 4175 -280 4185 -220
rect 4245 -280 4255 -220
rect 4175 -285 4255 -280
rect 4575 -110 4655 -105
rect 4575 -170 4585 -110
rect 4645 -170 4655 -110
rect 4575 -220 4655 -170
rect 4575 -280 4585 -220
rect 4645 -280 4655 -220
rect 4575 -285 4655 -280
rect 4975 -110 5055 -105
rect 4975 -170 4985 -110
rect 5045 -170 5055 -110
rect 4975 -220 5055 -170
rect 4975 -280 4985 -220
rect 5045 -280 5055 -220
rect 4975 -285 5055 -280
rect 5375 -110 5455 -105
rect 5375 -170 5385 -110
rect 5445 -170 5455 -110
rect 5375 -220 5455 -170
rect 5375 -280 5385 -220
rect 5445 -280 5455 -220
rect 5375 -285 5455 -280
rect 5775 -110 5855 -105
rect 5775 -170 5785 -110
rect 5845 -170 5855 -110
rect 5775 -220 5855 -170
rect 5775 -280 5785 -220
rect 5845 -280 5855 -220
rect 5775 -285 5855 -280
rect 6175 -110 6255 -105
rect 6175 -170 6185 -110
rect 6245 -170 6255 -110
rect 6175 -220 6255 -170
rect 6175 -280 6185 -220
rect 6245 -280 6255 -220
rect 6175 -285 6255 -280
rect 6575 -110 6655 -105
rect 6575 -170 6585 -110
rect 6645 -170 6655 -110
rect 6575 -220 6655 -170
rect 6575 -280 6585 -220
rect 6645 -280 6655 -220
rect 6575 -285 6655 -280
rect 6975 -110 7055 -105
rect 6975 -170 6985 -110
rect 7045 -170 7055 -110
rect 6975 -220 7055 -170
rect 6975 -280 6985 -220
rect 7045 -280 7055 -220
rect 6975 -285 7055 -280
rect 7375 -110 7455 -105
rect 7375 -170 7385 -110
rect 7445 -170 7455 -110
rect 7375 -220 7455 -170
rect 7375 -280 7385 -220
rect 7445 -280 7455 -220
rect 7375 -285 7455 -280
rect 7775 -110 7855 -105
rect 7775 -170 7785 -110
rect 7845 -170 7855 -110
rect 7775 -220 7855 -170
rect 7775 -280 7785 -220
rect 7845 -280 7855 -220
rect 7775 -285 7855 -280
rect 8175 -110 8255 -105
rect 8175 -170 8185 -110
rect 8245 -170 8255 -110
rect 8175 -220 8255 -170
rect 8175 -280 8185 -220
rect 8245 -280 8255 -220
rect 8175 -285 8255 -280
rect 8575 -110 8655 -105
rect 8575 -170 8585 -110
rect 8645 -170 8655 -110
rect 8575 -220 8655 -170
rect 8575 -280 8585 -220
rect 8645 -280 8655 -220
rect 8575 -285 8655 -280
rect 8975 -110 9055 -105
rect 8975 -170 8985 -110
rect 9045 -170 9055 -110
rect 8975 -220 9055 -170
rect 8975 -280 8985 -220
rect 9045 -280 9055 -220
rect 8975 -285 9055 -280
rect 9375 -110 9455 -105
rect 9375 -170 9385 -110
rect 9445 -170 9455 -110
rect 9375 -220 9455 -170
rect 9375 -280 9385 -220
rect 9445 -280 9455 -220
rect 9375 -285 9455 -280
rect 9775 -110 9855 -105
rect 9775 -170 9785 -110
rect 9845 -170 9855 -110
rect 9775 -220 9855 -170
rect 9775 -280 9785 -220
rect 9845 -280 9855 -220
rect 9775 -285 9855 -280
rect 10175 -110 10255 -105
rect 10175 -170 10185 -110
rect 10245 -170 10255 -110
rect 10175 -220 10255 -170
rect 10175 -280 10185 -220
rect 10245 -280 10255 -220
rect 10175 -285 10255 -280
rect 10575 -110 10655 -105
rect 10575 -170 10585 -110
rect 10645 -170 10655 -110
rect 10575 -220 10655 -170
rect 10575 -280 10585 -220
rect 10645 -280 10655 -220
rect 10575 -285 10655 -280
rect 10975 -110 11055 -105
rect 10975 -170 10985 -110
rect 11045 -170 11055 -110
rect 10975 -220 11055 -170
rect 10975 -280 10985 -220
rect 11045 -280 11055 -220
rect 10975 -285 11055 -280
rect 11375 -110 11455 -105
rect 11375 -170 11385 -110
rect 11445 -170 11455 -110
rect 11375 -220 11455 -170
rect 11375 -280 11385 -220
rect 11445 -280 11455 -220
rect 11375 -285 11455 -280
rect 11775 -110 11855 -105
rect 11775 -170 11785 -110
rect 11845 -170 11855 -110
rect 11775 -220 11855 -170
rect 11775 -280 11785 -220
rect 11845 -280 11855 -220
rect 11775 -285 11855 -280
rect 12175 -110 12255 -105
rect 12175 -170 12185 -110
rect 12245 -170 12255 -110
rect 12175 -220 12255 -170
rect 12175 -280 12185 -220
rect 12245 -280 12255 -220
rect 12175 -285 12255 -280
rect 12575 -110 12655 -105
rect 12575 -170 12585 -110
rect 12645 -170 12655 -110
rect 12575 -220 12655 -170
rect 12575 -280 12585 -220
rect 12645 -280 12655 -220
rect 12575 -285 12655 -280
rect 12975 -110 13055 -105
rect 12975 -170 12985 -110
rect 13045 -170 13055 -110
rect 12975 -220 13055 -170
rect 12975 -280 12985 -220
rect 13045 -280 13055 -220
rect 12975 -285 13055 -280
rect -215 -380 -155 -285
rect 185 -380 245 -285
rect 585 -380 645 -285
rect 985 -380 1045 -285
rect 1385 -380 1445 -285
rect 1785 -380 1845 -285
rect 2185 -380 2245 -285
rect 2585 -380 2645 -285
rect 2985 -380 3045 -285
rect 3385 -380 3445 -285
rect 3785 -380 3845 -285
rect 4185 -380 4245 -285
rect 4585 -380 4645 -285
rect 4985 -380 5045 -285
rect 5385 -380 5445 -285
rect 5785 -380 5845 -285
rect 6185 -380 6245 -285
rect 6585 -380 6645 -285
rect 6985 -380 7045 -285
rect 7385 -380 7445 -285
rect 7785 -380 7845 -285
rect 8185 -380 8245 -285
rect 8585 -380 8645 -285
rect 8985 -380 9045 -285
rect 9385 -380 9445 -285
rect 9785 -380 9845 -285
rect 10185 -380 10245 -285
rect 10585 -380 10645 -285
rect 10985 -380 11045 -285
rect 11385 -380 11445 -285
rect 11785 -380 11845 -285
rect 12185 -380 12245 -285
rect 12585 -380 12645 -285
rect 12985 -380 13045 -285
<< via3 >>
rect 12905 24125 12985 24135
rect 12905 24065 12915 24125
rect 12915 24065 12975 24125
rect 12975 24065 12985 24125
rect 12905 24055 12985 24065
rect 13035 24125 13115 24135
rect 13035 24065 13045 24125
rect 13045 24065 13105 24125
rect 13105 24065 13115 24125
rect 13035 24055 13115 24065
rect 180 23940 250 23945
rect 180 23880 185 23940
rect 185 23880 245 23940
rect 245 23880 250 23940
rect 180 23875 250 23880
rect 580 23940 650 23945
rect 580 23880 585 23940
rect 585 23880 645 23940
rect 645 23880 650 23940
rect 580 23875 650 23880
rect 980 23940 1050 23945
rect 980 23880 985 23940
rect 985 23880 1045 23940
rect 1045 23880 1050 23940
rect 980 23875 1050 23880
rect 1380 23940 1450 23945
rect 1380 23880 1385 23940
rect 1385 23880 1445 23940
rect 1445 23880 1450 23940
rect 1380 23875 1450 23880
rect 1780 23940 1850 23945
rect 1780 23880 1785 23940
rect 1785 23880 1845 23940
rect 1845 23880 1850 23940
rect 1780 23875 1850 23880
rect 2180 23940 2250 23945
rect 2180 23880 2185 23940
rect 2185 23880 2245 23940
rect 2245 23880 2250 23940
rect 2180 23875 2250 23880
rect 2580 23940 2650 23945
rect 2580 23880 2585 23940
rect 2585 23880 2645 23940
rect 2645 23880 2650 23940
rect 2580 23875 2650 23880
rect 2980 23940 3050 23945
rect 2980 23880 2985 23940
rect 2985 23880 3045 23940
rect 3045 23880 3050 23940
rect 2980 23875 3050 23880
rect 3380 23940 3450 23945
rect 3380 23880 3385 23940
rect 3385 23880 3445 23940
rect 3445 23880 3450 23940
rect 3380 23875 3450 23880
rect 3780 23940 3850 23945
rect 3780 23880 3785 23940
rect 3785 23880 3845 23940
rect 3845 23880 3850 23940
rect 3780 23875 3850 23880
rect 4180 23940 4250 23945
rect 4180 23880 4185 23940
rect 4185 23880 4245 23940
rect 4245 23880 4250 23940
rect 4180 23875 4250 23880
rect 4580 23940 4650 23945
rect 4580 23880 4585 23940
rect 4585 23880 4645 23940
rect 4645 23880 4650 23940
rect 4580 23875 4650 23880
rect 4980 23940 5050 23945
rect 4980 23880 4985 23940
rect 4985 23880 5045 23940
rect 5045 23880 5050 23940
rect 4980 23875 5050 23880
rect 5380 23940 5450 23945
rect 5380 23880 5385 23940
rect 5385 23880 5445 23940
rect 5445 23880 5450 23940
rect 5380 23875 5450 23880
rect 5780 23940 5850 23945
rect 5780 23880 5785 23940
rect 5785 23880 5845 23940
rect 5845 23880 5850 23940
rect 5780 23875 5850 23880
rect 6180 23940 6250 23945
rect 6180 23880 6185 23940
rect 6185 23880 6245 23940
rect 6245 23880 6250 23940
rect 6180 23875 6250 23880
rect 6580 23940 6650 23945
rect 6580 23880 6585 23940
rect 6585 23880 6645 23940
rect 6645 23880 6650 23940
rect 6580 23875 6650 23880
rect 6980 23940 7050 23945
rect 6980 23880 6985 23940
rect 6985 23880 7045 23940
rect 7045 23880 7050 23940
rect 6980 23875 7050 23880
rect 7380 23940 7450 23945
rect 7380 23880 7385 23940
rect 7385 23880 7445 23940
rect 7445 23880 7450 23940
rect 7380 23875 7450 23880
rect 7780 23940 7850 23945
rect 7780 23880 7785 23940
rect 7785 23880 7845 23940
rect 7845 23880 7850 23940
rect 7780 23875 7850 23880
rect 8180 23940 8250 23945
rect 8180 23880 8185 23940
rect 8185 23880 8245 23940
rect 8245 23880 8250 23940
rect 8180 23875 8250 23880
rect 8580 23940 8650 23945
rect 8580 23880 8585 23940
rect 8585 23880 8645 23940
rect 8645 23880 8650 23940
rect 8580 23875 8650 23880
rect 8980 23940 9050 23945
rect 8980 23880 8985 23940
rect 8985 23880 9045 23940
rect 9045 23880 9050 23940
rect 8980 23875 9050 23880
rect 9380 23940 9450 23945
rect 9380 23880 9385 23940
rect 9385 23880 9445 23940
rect 9445 23880 9450 23940
rect 9380 23875 9450 23880
rect 9780 23940 9850 23945
rect 9780 23880 9785 23940
rect 9785 23880 9845 23940
rect 9845 23880 9850 23940
rect 9780 23875 9850 23880
rect 10180 23940 10250 23945
rect 10180 23880 10185 23940
rect 10185 23880 10245 23940
rect 10245 23880 10250 23940
rect 10180 23875 10250 23880
rect 10580 23940 10650 23945
rect 10580 23880 10585 23940
rect 10585 23880 10645 23940
rect 10645 23880 10650 23940
rect 10580 23875 10650 23880
rect 10980 23940 11050 23945
rect 10980 23880 10985 23940
rect 10985 23880 11045 23940
rect 11045 23880 11050 23940
rect 10980 23875 11050 23880
rect 11380 23940 11450 23945
rect 11380 23880 11385 23940
rect 11385 23880 11445 23940
rect 11445 23880 11450 23940
rect 11380 23875 11450 23880
rect 11780 23940 11850 23945
rect 11780 23880 11785 23940
rect 11785 23880 11845 23940
rect 11845 23880 11850 23940
rect 11780 23875 11850 23880
rect 12180 23940 12250 23945
rect 12180 23880 12185 23940
rect 12185 23880 12245 23940
rect 12245 23880 12250 23940
rect 12180 23875 12250 23880
rect 12580 23940 12650 23945
rect 12580 23880 12585 23940
rect 12585 23880 12645 23940
rect 12645 23880 12650 23940
rect 12580 23875 12650 23880
<< metal4 >>
rect 180 24075 12650 24145
rect 180 23946 250 24075
rect 580 23946 650 24075
rect 980 23946 1050 24075
rect 1380 23946 1450 24075
rect 1780 23946 1850 24075
rect 2180 23946 2250 24075
rect 2580 23946 2650 24075
rect 2980 23946 3050 24075
rect 3380 23946 3450 24075
rect 3780 23946 3850 24075
rect 4180 23946 4250 24075
rect 4580 23946 4650 24075
rect 4980 23946 5050 24075
rect 5380 23946 5450 24075
rect 5780 23946 5850 24075
rect 6180 23946 6250 24075
rect 6580 23946 6650 24075
rect 6980 23946 7050 24075
rect 7380 23946 7450 24075
rect 7780 23946 7850 24075
rect 8180 23946 8250 24075
rect 8580 23946 8650 24075
rect 8980 23946 9050 24075
rect 9380 23946 9450 24075
rect 9780 23946 9850 24075
rect 10180 23946 10250 24075
rect 10580 23946 10650 24075
rect 10980 23946 11050 24075
rect 11380 23946 11450 24075
rect 11780 23946 11850 24075
rect 12180 23946 12250 24075
rect 12580 23946 12650 24075
rect 12895 24135 13125 24145
rect 12895 24055 12905 24135
rect 12985 24055 13035 24135
rect 13115 24055 13125 24135
rect 12895 24045 13125 24055
rect 179 23945 251 23946
rect 179 23875 180 23945
rect 250 23875 251 23945
rect 179 23874 251 23875
rect 579 23945 651 23946
rect 579 23875 580 23945
rect 650 23875 651 23945
rect 579 23874 651 23875
rect 979 23945 1051 23946
rect 979 23875 980 23945
rect 1050 23875 1051 23945
rect 979 23874 1051 23875
rect 1379 23945 1451 23946
rect 1379 23875 1380 23945
rect 1450 23875 1451 23945
rect 1379 23874 1451 23875
rect 1779 23945 1851 23946
rect 1779 23875 1780 23945
rect 1850 23875 1851 23945
rect 1779 23874 1851 23875
rect 2179 23945 2251 23946
rect 2179 23875 2180 23945
rect 2250 23875 2251 23945
rect 2179 23874 2251 23875
rect 2579 23945 2651 23946
rect 2579 23875 2580 23945
rect 2650 23875 2651 23945
rect 2579 23874 2651 23875
rect 2979 23945 3051 23946
rect 2979 23875 2980 23945
rect 3050 23875 3051 23945
rect 2979 23874 3051 23875
rect 3379 23945 3451 23946
rect 3379 23875 3380 23945
rect 3450 23875 3451 23945
rect 3379 23874 3451 23875
rect 3779 23945 3851 23946
rect 3779 23875 3780 23945
rect 3850 23875 3851 23945
rect 3779 23874 3851 23875
rect 4179 23945 4251 23946
rect 4179 23875 4180 23945
rect 4250 23875 4251 23945
rect 4179 23874 4251 23875
rect 4579 23945 4651 23946
rect 4579 23875 4580 23945
rect 4650 23875 4651 23945
rect 4579 23874 4651 23875
rect 4979 23945 5051 23946
rect 4979 23875 4980 23945
rect 5050 23875 5051 23945
rect 4979 23874 5051 23875
rect 5379 23945 5451 23946
rect 5379 23875 5380 23945
rect 5450 23875 5451 23945
rect 5379 23874 5451 23875
rect 5779 23945 5851 23946
rect 5779 23875 5780 23945
rect 5850 23875 5851 23945
rect 5779 23874 5851 23875
rect 6179 23945 6251 23946
rect 6179 23875 6180 23945
rect 6250 23875 6251 23945
rect 6179 23874 6251 23875
rect 6579 23945 6651 23946
rect 6579 23875 6580 23945
rect 6650 23875 6651 23945
rect 6579 23874 6651 23875
rect 6979 23945 7051 23946
rect 6979 23875 6980 23945
rect 7050 23875 7051 23945
rect 6979 23874 7051 23875
rect 7379 23945 7451 23946
rect 7379 23875 7380 23945
rect 7450 23875 7451 23945
rect 7379 23874 7451 23875
rect 7779 23945 7851 23946
rect 7779 23875 7780 23945
rect 7850 23875 7851 23945
rect 7779 23874 7851 23875
rect 8179 23945 8251 23946
rect 8179 23875 8180 23945
rect 8250 23875 8251 23945
rect 8179 23874 8251 23875
rect 8579 23945 8651 23946
rect 8579 23875 8580 23945
rect 8650 23875 8651 23945
rect 8579 23874 8651 23875
rect 8979 23945 9051 23946
rect 8979 23875 8980 23945
rect 9050 23875 9051 23945
rect 8979 23874 9051 23875
rect 9379 23945 9451 23946
rect 9379 23875 9380 23945
rect 9450 23875 9451 23945
rect 9379 23874 9451 23875
rect 9779 23945 9851 23946
rect 9779 23875 9780 23945
rect 9850 23875 9851 23945
rect 9779 23874 9851 23875
rect 10179 23945 10251 23946
rect 10179 23875 10180 23945
rect 10250 23875 10251 23945
rect 10179 23874 10251 23875
rect 10579 23945 10651 23946
rect 10579 23875 10580 23945
rect 10650 23875 10651 23945
rect 10579 23874 10651 23875
rect 10979 23945 11051 23946
rect 10979 23875 10980 23945
rect 11050 23875 11051 23945
rect 10979 23874 11051 23875
rect 11379 23945 11451 23946
rect 11379 23875 11380 23945
rect 11450 23875 11451 23945
rect 11379 23874 11451 23875
rect 11779 23945 11851 23946
rect 11779 23875 11780 23945
rect 11850 23875 11851 23945
rect 11779 23874 11851 23875
rect 12179 23945 12251 23946
rect 12179 23875 12180 23945
rect 12250 23875 12251 23945
rect 12179 23874 12251 23875
rect 12579 23945 12651 23946
rect 12579 23875 12580 23945
rect 12650 23875 12651 23945
rect 12579 23874 12651 23875
<< labels >>
rlabel metal1 13360 3870 13380 3890 1 C10
port 12 n
rlabel metal1 13360 6090 13380 6110 1 C9
port 11 n
rlabel metal1 13360 7940 13380 7960 1 C8
port 10 n
rlabel metal1 13360 9050 13380 9070 1 C7
port 9 n
rlabel metal1 13360 9790 13380 9810 1 C6
port 8 n
rlabel metal1 13360 10160 13380 10180 1 C5
port 7 n
rlabel metal1 13360 10900 13380 10920 1 C4
port 6 n
rlabel metal1 13360 12750 13380 12770 1 C3
port 5 n
rlabel metal1 13360 11270 13380 11290 1 C2
port 4 n
rlabel metal1 13360 12380 13380 12400 1 C1
port 3 n
rlabel metal1 13360 12010 13380 12030 1 C0
port 2 n
rlabel metal1 13360 11640 13380 11660 1 C0_dummy
port 1 n
rlabel metal4 12975 24065 13035 24125 1 VSS
port 15 n
rlabel metal4 12390 24090 12495 24135 1 Ctop
port 14 n
<< end >>
