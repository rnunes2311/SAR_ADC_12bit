magic
tech sky130A
magscale 1 2
timestamp 1711796880
<< error_p >>
rect -415 481 -353 487
rect -287 481 -225 487
rect -159 481 -97 487
rect -31 481 31 487
rect 97 481 159 487
rect 225 481 287 487
rect 353 481 415 487
rect -415 447 -403 481
rect -287 447 -275 481
rect -159 447 -147 481
rect -31 447 -19 481
rect 97 447 109 481
rect 225 447 237 481
rect 353 447 365 481
rect -415 441 -353 447
rect -287 441 -225 447
rect -159 441 -97 447
rect -31 441 31 447
rect 97 441 159 447
rect 225 441 287 447
rect 353 441 415 447
rect -415 -447 -353 -441
rect -287 -447 -225 -441
rect -159 -447 -97 -441
rect -31 -447 31 -441
rect 97 -447 159 -441
rect 225 -447 287 -441
rect 353 -447 415 -441
rect -415 -481 -403 -447
rect -287 -481 -275 -447
rect -159 -481 -147 -447
rect -31 -481 -19 -447
rect 97 -481 109 -447
rect 225 -481 237 -447
rect 353 -481 365 -447
rect -415 -487 -353 -481
rect -287 -487 -225 -481
rect -159 -487 -97 -481
rect -31 -487 31 -481
rect 97 -487 159 -481
rect 225 -487 287 -481
rect 353 -487 415 -481
<< nwell >>
rect -513 -500 513 500
<< pmoslvt >>
rect -419 -400 -349 400
rect -291 -400 -221 400
rect -163 -400 -93 400
rect -35 -400 35 400
rect 93 -400 163 400
rect 221 -400 291 400
rect 349 -400 419 400
<< pdiff >>
rect -477 388 -419 400
rect -477 -388 -465 388
rect -431 -388 -419 388
rect -477 -400 -419 -388
rect -349 388 -291 400
rect -349 -388 -337 388
rect -303 -388 -291 388
rect -349 -400 -291 -388
rect -221 388 -163 400
rect -221 -388 -209 388
rect -175 -388 -163 388
rect -221 -400 -163 -388
rect -93 388 -35 400
rect -93 -388 -81 388
rect -47 -388 -35 388
rect -93 -400 -35 -388
rect 35 388 93 400
rect 35 -388 47 388
rect 81 -388 93 388
rect 35 -400 93 -388
rect 163 388 221 400
rect 163 -388 175 388
rect 209 -388 221 388
rect 163 -400 221 -388
rect 291 388 349 400
rect 291 -388 303 388
rect 337 -388 349 388
rect 291 -400 349 -388
rect 419 388 477 400
rect 419 -388 431 388
rect 465 -388 477 388
rect 419 -400 477 -388
<< pdiffc >>
rect -465 -388 -431 388
rect -337 -388 -303 388
rect -209 -388 -175 388
rect -81 -388 -47 388
rect 47 -388 81 388
rect 175 -388 209 388
rect 303 -388 337 388
rect 431 -388 465 388
<< poly >>
rect -419 481 -349 497
rect -419 447 -403 481
rect -365 447 -349 481
rect -419 400 -349 447
rect -291 481 -221 497
rect -291 447 -275 481
rect -237 447 -221 481
rect -291 400 -221 447
rect -163 481 -93 497
rect -163 447 -147 481
rect -109 447 -93 481
rect -163 400 -93 447
rect -35 481 35 497
rect -35 447 -19 481
rect 19 447 35 481
rect -35 400 35 447
rect 93 481 163 497
rect 93 447 109 481
rect 147 447 163 481
rect 93 400 163 447
rect 221 481 291 497
rect 221 447 237 481
rect 275 447 291 481
rect 221 400 291 447
rect 349 481 419 497
rect 349 447 365 481
rect 403 447 419 481
rect 349 400 419 447
rect -419 -447 -349 -400
rect -419 -481 -403 -447
rect -365 -481 -349 -447
rect -419 -497 -349 -481
rect -291 -447 -221 -400
rect -291 -481 -275 -447
rect -237 -481 -221 -447
rect -291 -497 -221 -481
rect -163 -447 -93 -400
rect -163 -481 -147 -447
rect -109 -481 -93 -447
rect -163 -497 -93 -481
rect -35 -447 35 -400
rect -35 -481 -19 -447
rect 19 -481 35 -447
rect -35 -497 35 -481
rect 93 -447 163 -400
rect 93 -481 109 -447
rect 147 -481 163 -447
rect 93 -497 163 -481
rect 221 -447 291 -400
rect 221 -481 237 -447
rect 275 -481 291 -447
rect 221 -497 291 -481
rect 349 -447 419 -400
rect 349 -481 365 -447
rect 403 -481 419 -447
rect 349 -497 419 -481
<< polycont >>
rect -403 447 -365 481
rect -275 447 -237 481
rect -147 447 -109 481
rect -19 447 19 481
rect 109 447 147 481
rect 237 447 275 481
rect 365 447 403 481
rect -403 -481 -365 -447
rect -275 -481 -237 -447
rect -147 -481 -109 -447
rect -19 -481 19 -447
rect 109 -481 147 -447
rect 237 -481 275 -447
rect 365 -481 403 -447
<< locali >>
rect -419 447 -403 481
rect -365 447 -349 481
rect -291 447 -275 481
rect -237 447 -221 481
rect -163 447 -147 481
rect -109 447 -93 481
rect -35 447 -19 481
rect 19 447 35 481
rect 93 447 109 481
rect 147 447 163 481
rect 221 447 237 481
rect 275 447 291 481
rect 349 447 365 481
rect 403 447 419 481
rect -465 388 -431 404
rect -465 -404 -431 -388
rect -337 388 -303 404
rect -337 -404 -303 -388
rect -209 388 -175 404
rect -209 -404 -175 -388
rect -81 388 -47 404
rect -81 -404 -47 -388
rect 47 388 81 404
rect 47 -404 81 -388
rect 175 388 209 404
rect 175 -404 209 -388
rect 303 388 337 404
rect 303 -404 337 -388
rect 431 388 465 404
rect 431 -404 465 -388
rect -419 -481 -403 -447
rect -365 -481 -349 -447
rect -291 -481 -275 -447
rect -237 -481 -221 -447
rect -163 -481 -147 -447
rect -109 -481 -93 -447
rect -35 -481 -19 -447
rect 19 -481 35 -447
rect 93 -481 109 -447
rect 147 -481 163 -447
rect 221 -481 237 -447
rect 275 -481 291 -447
rect 349 -481 365 -447
rect 403 -481 419 -447
<< viali >>
rect -403 447 -365 481
rect -275 447 -237 481
rect -147 447 -109 481
rect -19 447 19 481
rect 109 447 147 481
rect 237 447 275 481
rect 365 447 403 481
rect -465 -388 -431 388
rect -337 -388 -303 388
rect -209 -388 -175 388
rect -81 -388 -47 388
rect 47 -388 81 388
rect 175 -388 209 388
rect 303 -388 337 388
rect 431 -388 465 388
rect -403 -481 -365 -447
rect -275 -481 -237 -447
rect -147 -481 -109 -447
rect -19 -481 19 -447
rect 109 -481 147 -447
rect 237 -481 275 -447
rect 365 -481 403 -447
<< metal1 >>
rect -415 481 -353 487
rect -415 447 -403 481
rect -365 447 -353 481
rect -415 441 -353 447
rect -287 481 -225 487
rect -287 447 -275 481
rect -237 447 -225 481
rect -287 441 -225 447
rect -159 481 -97 487
rect -159 447 -147 481
rect -109 447 -97 481
rect -159 441 -97 447
rect -31 481 31 487
rect -31 447 -19 481
rect 19 447 31 481
rect -31 441 31 447
rect 97 481 159 487
rect 97 447 109 481
rect 147 447 159 481
rect 97 441 159 447
rect 225 481 287 487
rect 225 447 237 481
rect 275 447 287 481
rect 225 441 287 447
rect 353 481 415 487
rect 353 447 365 481
rect 403 447 415 481
rect 353 441 415 447
rect -471 388 -425 400
rect -471 -388 -465 388
rect -431 -388 -425 388
rect -471 -400 -425 -388
rect -343 388 -297 400
rect -343 -388 -337 388
rect -303 -388 -297 388
rect -343 -400 -297 -388
rect -215 388 -169 400
rect -215 -388 -209 388
rect -175 -388 -169 388
rect -215 -400 -169 -388
rect -87 388 -41 400
rect -87 -388 -81 388
rect -47 -388 -41 388
rect -87 -400 -41 -388
rect 41 388 87 400
rect 41 -388 47 388
rect 81 -388 87 388
rect 41 -400 87 -388
rect 169 388 215 400
rect 169 -388 175 388
rect 209 -388 215 388
rect 169 -400 215 -388
rect 297 388 343 400
rect 297 -388 303 388
rect 337 -388 343 388
rect 297 -400 343 -388
rect 425 388 471 400
rect 425 -388 431 388
rect 465 -388 471 388
rect 425 -400 471 -388
rect -415 -447 -353 -441
rect -415 -481 -403 -447
rect -365 -481 -353 -447
rect -415 -487 -353 -481
rect -287 -447 -225 -441
rect -287 -481 -275 -447
rect -237 -481 -225 -447
rect -287 -487 -225 -481
rect -159 -447 -97 -441
rect -159 -481 -147 -447
rect -109 -481 -97 -447
rect -159 -487 -97 -481
rect -31 -447 31 -441
rect -31 -481 -19 -447
rect 19 -481 31 -447
rect -31 -487 31 -481
rect 97 -447 159 -441
rect 97 -481 109 -447
rect 147 -481 159 -447
rect 97 -487 159 -481
rect 225 -447 287 -441
rect 225 -481 237 -447
rect 275 -481 287 -447
rect 225 -487 287 -481
rect 353 -447 415 -441
rect 353 -481 365 -447
rect 403 -481 415 -447
rect 353 -487 415 -481
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 4 l 0.35 m 1 nf 7 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
