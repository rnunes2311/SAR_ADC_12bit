* SPICE3 file created from SAR_ADC_12bit_flat.ext - technology: sky130A

.subckt SAR_ADC_12bit VDD VCM VSS VREF VIN_P VIN_N RST_Z CLK_DATA DATA[5] DATA[4] DATA[3] DATA[2] DATA[1] DATA[0] START EN_OFFSET_CAL CLK VREF_GND
+ SINGLE_ENDED
X0 a_13076_44458# a_13259_45724# a_13296_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2 VSS a_12427_45724# a_10490_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VDD a_2324_44458# a_949_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=361.2627 ps=3.22652k w=0.87 l=2.89
X5 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X6 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X7 VDD a_2903_42308# a_3080_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8 VDD a_12861_44030# a_17829_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VSS a_1209_43370# a_n1557_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_16237_45028# a_16147_45260# a_16019_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_2075_43172# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VDD a_n755_45592# a_1176_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X13 a_6756_44260# a_5937_45572# a_6453_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X14 a_15868_43402# a_15681_43442# a_15781_43660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X15 a_n1533_42852# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X16 a_8103_44636# a_8375_44464# a_8333_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 VSS a_16327_47482# a_16377_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X18 a_2437_43646# a_n443_46116# a_2437_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_5088_37509# VSS VDAC_Ni VDD sky130_fd_pr__pfet_01v8_hvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X20 a_n2810_45028# a_n2840_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X21 a_2113_38308# VDAC_Ni a_2112_39137# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X22 VDD a_3626_43646# a_19647_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X23 VSS a_10334_44484# a_10440_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X24 a_1576_42282# a_1755_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X25 a_10933_46660# a_10554_47026# a_10861_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X26 a_14021_43940# a_13483_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X27 a_16867_43762# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X28 VREF a_21076_30879# C8_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X29 VSS a_n2946_37690# a_n3565_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 a_n913_45002# a_1307_43914# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 a_n2840_43370# a_n2661_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X32 a_3457_43396# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X33 a_14180_46482# a_14035_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X34 VSS a_18989_43940# a_19006_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X35 VSS a_9672_43914# a_2107_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X36 a_n1059_45260# a_17499_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X37 VSS a_10695_43548# a_10057_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X38 a_n2104_42282# a_n1925_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X39 a_20749_43396# a_12549_44172# a_743_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X40 VDD a_3877_44458# a_2382_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X41 a_n1699_44726# a_n1917_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X42 VSS a_n4334_39616# a_n4064_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X43 a_9241_45822# a_5066_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X44 VDD a_12883_44458# a_n2293_43922# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X45 a_11909_44484# a_3232_43370# a_11827_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X46 a_835_46155# a_584_46384# a_376_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X47 VSS a_1666_39043# a_1169_39043# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X48 a_5210_46155# a_5164_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X49 VDD a_n3690_39392# a_n3420_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X50 VDD a_167_45260# a_1609_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X51 VSS a_526_44458# a_3363_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X52 a_19268_43646# a_19319_43548# a_19095_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X53 VSS a_22959_44484# a_19237_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X54 a_n2216_39072# a_n2312_39304# a_n2302_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X55 a_19987_42826# a_10193_42453# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X56 a_6151_47436# a_14311_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X57 a_8145_46902# a_7927_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X58 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X59 a_14275_46494# a_13925_46122# a_14180_46482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X60 a_20512_43084# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X61 a_14539_43914# a_17701_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X62 a_6298_44484# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X63 a_644_44056# a_626_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X64 a_10949_43914# a_12429_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.28 ps=2.56 w=1 l=0.15
X65 VSS a_n2302_39866# a_n4209_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X66 VSS a_21811_47423# a_20916_46384# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X67 VDD a_3699_46634# a_3686_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X68 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X69 a_8035_47026# a_7411_46660# a_7927_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X70 a_5691_45260# a_5111_44636# a_5837_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X71 VDD a_1307_43914# a_1241_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X72 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X73 a_18249_42858# a_18083_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X74 VDD a_104_43370# a_n971_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X75 VDD a_n2833_47464# CLK_DATA VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X76 a_3363_44484# a_1823_45246# a_3232_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X77 a_n1331_43914# a_n1549_44318# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X78 VCM a_4958_30871# C9_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X79 VSS a_n3565_39590# a_n3607_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X80 VSS a_12281_43396# a_12563_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X81 VSS a_18780_47178# a_13661_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X82 a_n4318_39768# a_n2840_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X83 DATA[5] a_11459_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X84 a_7230_45938# a_6472_45840# a_6667_45809# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X85 VDD a_8049_45260# a_22959_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X86 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X87 a_8746_45002# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X88 a_15004_44636# a_11691_44458# a_15146_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X89 a_16223_45938# a_15599_45572# a_16115_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X90 a_n984_44318# a_n1899_43946# a_n1331_43914# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X91 a_n809_44244# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X92 a_n4064_39616# a_n4334_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X93 a_17124_42282# a_17303_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X94 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X95 VSS a_3065_45002# a_2680_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X96 a_5193_42852# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X97 VDD a_6969_46634# a_6999_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X98 VDD a_10623_46897# a_10554_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X99 a_16137_43396# a_15781_43660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X100 VDD a_n2472_46634# a_n2442_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X101 VDD a_4185_45028# a_22959_45036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X102 a_15225_45822# a_15037_45618# a_15143_45578# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X103 VSS a_3537_45260# a_4640_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X104 a_n2012_43396# a_n2129_43609# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X105 VDD a_n13_43084# a_n1853_43023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X106 a_5068_46348# a_n1151_42308# a_5210_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X107 a_873_42968# a_685_42968# a_791_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X108 a_17730_32519# a_22591_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X109 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X110 VDD a_22485_44484# a_20974_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X111 a_n1021_46688# a_n1151_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X112 VSS a_11599_46634# a_11735_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X113 a_13163_45724# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.14075 ps=1.325 w=0.42 l=0.15
X114 C9_P_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X115 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X116 a_n2012_44484# a_n2129_44697# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X117 a_13940_44484# a_13556_45296# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X118 VSS a_1414_42308# a_1525_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X119 a_8487_44056# a_4223_44672# a_8415_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X120 a_18194_35068# a_n1794_35242# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X121 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X122 a_16434_46660# a_16388_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X123 a_22613_38993# a_22527_39145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X124 a_3315_47570# a_n1151_42308# a_2952_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X125 a_2680_45002# a_1823_45246# a_2903_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X126 a_1307_43914# a_2779_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X127 a_22731_47423# SMPL_ON_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X128 VDD a_1307_43914# a_3681_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X129 a_n863_45724# a_1667_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X130 VDD a_11459_47204# DATA[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X131 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X132 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X133 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=218.18214 ps=2.11206k w=0.55 l=0.59
X134 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X135 a_n4209_38216# a_n2302_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X136 VSS a_n1794_35242# a_18194_35068# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X137 a_10467_46802# a_11599_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X138 VDD a_13747_46662# a_19862_44208# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X139 a_n2946_39866# a_n2956_39768# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X140 a_n1013_45572# a_n1079_45724# a_n1099_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.182 ps=1.86 w=0.65 l=0.15
X141 VSS a_15279_43071# a_14579_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X142 DATA[3] a_7227_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X143 VSS a_8049_45260# a_22959_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X144 a_7584_44260# a_7542_44172# a_7281_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X145 a_n97_42460# a_19700_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X146 VDD a_19647_42308# a_13258_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X147 a_3754_39466# a_7754_39300# VSS sky130_fd_pr__res_high_po_0p35 l=18
X148 VSS a_2952_47436# a_2747_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X149 VDD a_16751_45260# a_6171_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X150 a_18326_43940# a_18079_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X151 a_9248_44260# a_8270_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X152 a_3503_45724# a_3775_45552# a_3733_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X153 a_n2017_45002# a_19987_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X154 a_288_46660# a_171_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X155 a_10037_46155# a_9804_47204# a_9823_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X156 a_20075_46420# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X157 VDD a_196_42282# a_n3674_37592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X158 VSS a_14513_46634# a_14447_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X159 a_n4064_39072# a_n4334_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X160 a_1149_42558# a_961_42354# a_1067_42314# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X161 a_13569_47204# a_13381_47204# a_13487_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X162 VDD a_14840_46494# a_15015_46420# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X163 C6_P_btm a_n3565_39304# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=0.35
X164 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X165 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X166 a_14537_43396# a_14358_43442# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X167 VDD a_14955_47212# a_10227_46804# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X168 VDD a_7754_40130# a_11206_38545# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X169 a_n3565_39590# a_n2946_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X170 a_n901_43156# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X171 a_17668_45572# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X172 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X173 a_15493_43396# a_14955_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X174 a_7309_43172# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X175 VDD a_1138_42852# a_1337_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X176 a_1427_43646# a_1568_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X177 a_18184_42460# a_15743_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X178 VDD a_13351_46090# a_10903_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X179 a_8379_46155# a_8128_46384# a_7920_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X180 VSS a_3483_46348# a_17325_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X181 VDD a_9290_44172# a_10949_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X182 VSS a_11823_42460# a_14358_43442# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X183 a_18310_42308# a_10193_42453# a_18220_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X184 VDD a_n2288_47178# a_n2312_40392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X185 a_17719_45144# a_16375_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X186 VDD a_5891_43370# a_5147_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X187 a_7287_43370# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X188 a_11173_44260# a_2063_45854# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X189 EN_VIN_BSTR_P VDD a_n1550_35608# VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.9
X190 a_11897_42308# a_11823_42460# a_11551_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X191 VDD a_12861_44030# a_13759_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X192 a_19466_46812# a_19778_44110# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X193 a_9049_44484# a_8701_44490# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X194 a_n3565_38502# a_n2946_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X195 VDD a_16588_47582# a_16763_47508# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X196 a_9396_43370# a_4883_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X197 C0_P_btm a_n784_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X198 a_n1736_42282# a_n1557_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X199 VDD a_14113_42308# a_16522_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X200 a_10651_43940# a_3090_45724# a_10555_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X201 VDD a_8667_46634# a_n237_47217# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X202 a_6123_31319# a_7227_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X203 a_7499_43078# a_10083_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X204 VSS a_n755_45592# a_1145_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X205 C7_P_btm a_5534_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X206 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X207 VSS a_n4064_37984# a_n2302_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X208 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X209 a_3581_42558# a_3539_42460# a_3497_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X210 a_n3674_38680# a_n2840_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X211 VSS a_5907_45546# a_5937_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X212 VDD a_22589_40055# a_22527_39145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X213 a_18783_43370# a_15743_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X214 VSS a_1799_45572# a_1983_46706# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X215 VDD a_22959_46660# a_21076_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X216 a_13467_32519# a_21487_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X217 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X218 a_2864_46660# a_2747_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X219 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X220 a_8199_44636# a_10355_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X221 a_14403_45348# a_13259_45724# a_14309_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X222 a_556_44484# a_742_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X223 VSS a_15433_44458# a_15367_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X224 a_n1794_35242# a_564_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X225 a_n2840_43370# a_n2661_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X226 VSS a_13747_46662# a_13693_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X227 a_18245_44484# a_17767_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X228 a_19741_43940# a_19862_44208# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X229 a_16855_43396# a_16409_43396# a_16759_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X230 a_n1696_35090# a_n1794_35242# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X231 a_13113_42826# a_12895_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X232 VSS a_22365_46825# a_20202_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X233 a_n1079_45724# a_n755_45592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X234 a_19386_47436# a_19321_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X235 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X236 VSS a_526_44458# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X237 a_n89_47570# a_n237_47217# a_n452_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X238 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X239 a_1176_45822# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X240 a_10341_43396# a_9803_43646# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X241 w_11334_34010# a_11530_34132# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=10.615 ps=76.96 w=3.75 l=15
X242 VDD a_n4209_38502# a_n4334_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X243 a_5111_42852# a_4905_42826# a_5193_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X244 a_13887_32519# a_22223_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X245 a_5437_45600# a_n881_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X246 a_18953_45572# a_18909_45814# a_18787_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X247 VDD a_4791_45118# a_6165_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X248 VDD a_3429_45260# a_3316_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.28 ps=2.56 w=1 l=0.15
X249 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X250 a_n3607_39616# a_n3674_39768# a_n3690_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X251 a_4842_47570# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X252 a_1337_46116# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X253 a_11136_45572# a_11322_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X254 a_n2661_42834# a_10809_44734# a_12189_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X255 VSS a_10249_46116# a_11186_47026# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X256 a_16655_46660# a_n743_46660# a_16292_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X257 a_n1991_46122# a_n2157_46122# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X258 VREF_GND a_n3420_39072# C6_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X259 a_n3565_37414# a_n2946_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X260 VDD a_1576_42282# a_1606_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X261 a_5159_47243# a_n443_46116# a_4700_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X262 VSS a_5891_43370# a_8375_44464# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X263 a_2075_43172# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X264 VDD a_13076_44458# a_12883_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X265 VSS a_14539_43914# a_14485_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X266 C0_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X267 a_15297_45822# a_11823_42460# a_15225_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X268 VDD a_1169_39043# comp_n VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X269 a_18479_47436# a_20075_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X270 a_1423_45028# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X271 a_2382_45260# a_3877_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X272 a_8103_44636# a_8199_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X273 a_n1899_43946# a_n2065_43946# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X274 a_6765_43638# a_6547_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X275 VSS a_22400_42852# a_22848_40945# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X276 a_n2293_43922# a_12741_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X277 a_n3565_38216# a_n2946_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X278 VDD a_n3690_39392# a_n3420_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X279 a_945_42968# a_n1059_45260# a_873_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X280 VDD a_3785_47178# a_3815_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X281 VDD a_14084_46812# a_14035_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X282 a_765_45546# a_12549_44172# a_17829_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X283 VDD a_20974_43370# a_20556_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X284 a_14275_46494# a_13759_46122# a_14180_46482# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X285 VSS a_15051_42282# a_11823_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X286 a_1609_45822# a_n443_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X287 a_17517_44484# a_16979_44734# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X288 VDD a_4915_47217# a_12891_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X289 a_20679_44626# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X290 VSS a_1423_45028# a_9838_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X291 a_13921_42308# a_13259_45724# a_13575_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X292 VCM a_n784_42308# C0_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X293 VSS a_11599_46634# a_13759_46122# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X294 a_14127_45572# a_11823_42460# a_14033_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X295 a_13569_43230# a_12379_42858# a_13460_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X296 a_5072_46660# a_4955_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X297 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X298 a_8037_42858# a_7871_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X299 VSS a_22591_46660# a_20820_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X300 VDD a_n2833_47464# CLK_DATA VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X301 a_3686_47026# a_2609_46660# a_3524_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X302 a_9672_43914# a_10057_43914# a_9801_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X303 VDD a_18429_43548# a_16823_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X304 a_17339_46660# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X305 VSS a_1606_42308# a_2351_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X306 a_16409_43396# a_16243_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X307 VSS a_9625_46129# a_10044_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X308 VDD a_n4209_37414# a_n4334_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X309 a_13468_44734# a_768_44030# a_13213_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X310 VSS a_n2302_39072# a_n4209_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X311 a_2124_47436# a_584_46384# a_2266_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X312 VDD a_n971_45724# a_2809_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X313 a_10809_44734# a_2063_45854# a_10809_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X314 a_7577_46660# a_7411_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X315 a_4921_42308# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X316 a_16023_47582# a_15507_47210# a_15928_47570# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X317 a_12791_45546# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X318 a_10193_42453# a_20712_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X319 VSS a_n881_46662# a_n659_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X320 a_6481_42558# a_n913_45002# a_1755_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X321 a_n2956_38680# a_n2472_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X322 a_14955_43940# a_14537_43396# a_15037_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X323 VREF_GND a_14097_32519# C4_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X324 VDD a_21188_45572# a_21363_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X325 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X326 a_15682_43940# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X327 a_18907_42674# a_18727_42674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X328 a_12545_42858# a_12379_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X329 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X330 C9_P_btm a_n4064_39616# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X331 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X332 a_13720_44458# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X333 a_15125_43396# a_15095_43370# a_15037_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X334 VREF a_20692_30879# C6_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=0.35
X335 a_2998_44172# a_584_46384# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X336 a_20974_43370# a_22485_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X337 a_18548_42308# a_18494_42460# a_18057_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X338 a_n875_44318# a_n2065_43946# a_n984_44318# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X339 w_11334_34010# a_18194_35068# EN_VIN_BSTR_N w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X340 a_n2293_42834# a_8049_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X341 VSS a_4743_44484# a_4791_45118# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X342 a_3626_43646# a_3232_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X343 VDD a_19998_35138# a_21753_35634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X344 VSS a_n2438_43548# a_n2433_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X345 a_n1076_43230# a_n2157_42858# a_n1423_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X346 VDD a_17973_43940# a_18079_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X347 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X348 VREF_GND a_17538_32519# C8_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X349 VDD a_22223_46124# a_20205_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X350 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X351 a_4704_46090# a_4883_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X352 a_5815_47464# a_6151_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X353 a_17478_45572# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X354 DATA[3] a_7227_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X355 a_18194_35068# a_n1794_35242# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X356 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X357 a_17034_45572# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X358 VSS a_n3420_39616# a_n2946_39866# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X359 a_133_42852# a_n97_42460# a_n13_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X360 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X361 a_n1925_46634# a_8162_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X362 a_21350_47026# a_20273_46660# a_21188_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X363 VDD a_2713_42308# a_2903_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X364 a_n3674_39304# a_n2840_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X365 a_13565_43940# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X366 a_n4315_30879# a_n2302_40160# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X367 VDD a_1823_45246# a_2202_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X368 VSS a_n3690_38304# a_n3420_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X369 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X370 a_2211_45572# a_2063_45854# a_1848_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X371 VSS a_16112_44458# a_14673_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X372 VSS a_3316_45546# a_3260_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X373 VDD a_n443_46116# a_2896_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X374 a_n310_47570# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X375 a_21177_47436# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X376 VSS a_9290_44172# a_13943_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X377 a_n3674_37592# a_196_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X378 a_18780_47178# a_18597_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X379 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X380 VSS a_8791_42308# a_5934_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X381 a_421_43172# a_n97_42460# a_n13_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X382 VDD a_17339_46660# a_18051_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X383 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X384 VSS a_n2840_46090# a_n2956_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X385 a_n2661_43370# a_10907_45822# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X386 a_9396_43370# a_4883_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X387 VDD a_19333_46634# a_19123_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X388 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X389 a_5755_42852# a_n97_42460# a_5837_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X390 a_n4251_39392# a_n4318_39304# a_n4334_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X391 a_805_46414# a_472_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X392 VDD a_n1076_43230# a_n901_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X393 a_21845_43940# a_12549_44172# a_19692_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X394 VDD a_4520_42826# a_4093_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X395 a_12469_46902# a_12251_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X396 a_15415_45028# a_15227_44166# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X397 a_19479_31679# a_22223_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X398 a_7542_44172# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X399 a_3080_42308# a_2903_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X400 VSS a_22165_42308# a_22223_42860# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X401 VDD a_10249_46116# a_11186_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X402 a_3905_42558# a_2382_45260# a_3823_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X403 a_12347_46660# a_11901_46660# a_12251_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X404 VSS a_16137_43396# a_16414_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.089375 ps=0.925 w=0.65 l=0.15
X405 a_5066_45546# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X406 a_14581_44484# a_13249_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X407 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X408 a_2113_38308# a_1273_38525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X409 a_n473_42460# a_n755_45592# a_n327_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X410 VDD a_n1699_43638# a_n1809_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X411 a_13759_47204# a_13717_47436# a_13675_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X412 a_n3420_39616# a_n3690_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X413 C4_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X414 a_n967_46494# a_n2157_46122# a_n1076_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X415 a_2779_44458# a_1423_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X416 VDD a_19319_43548# a_19268_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.195 ps=1.39 w=1 l=0.15
X417 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X418 VDD a_9127_43156# a_5891_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X419 a_1123_46634# a_948_46660# a_1302_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X420 a_n755_45592# a_n809_44244# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X421 a_2952_47436# a_3160_47472# a_3094_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X422 a_5807_45002# a_16763_47508# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X423 a_3726_37500# a_3754_38470# VDAC_Ni VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X424 a_6293_42852# a_5755_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X425 a_8120_45572# a_8034_45724# a_n1925_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X426 a_11541_44484# a_11691_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X427 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X428 VSS a_10083_42826# a_7499_43078# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X429 a_5257_43370# a_5907_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X430 a_4880_45572# a_5066_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X431 VIN_P EN_VIN_BSTR_P C0_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X432 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X433 a_3497_42558# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X434 VSS a_1123_46634# a_584_46384# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X435 a_16223_45938# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X436 a_4883_46098# a_21363_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X437 a_2711_45572# a_768_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X438 VSS a_2553_47502# a_2487_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X439 VDD a_12469_46902# a_12359_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X440 a_6453_43914# a_6109_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X441 a_7765_42852# a_7227_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X442 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X443 a_17786_45822# a_15861_45028# a_17478_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X444 a_18450_45144# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X445 a_6765_43638# a_6547_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X446 a_n914_46116# a_n1991_46122# a_n1076_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X447 VSS a_n4334_40480# a_n4064_40160# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X448 a_12089_42308# a_11551_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X449 a_16547_43609# a_16414_43172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X450 a_3221_46660# a_3177_46902# a_3055_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X451 a_6667_45809# a_6472_45840# a_6977_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X452 a_n1190_43762# a_n2267_43396# a_n1352_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X453 a_6643_43396# a_6197_43396# a_6547_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X454 a_5837_45348# a_5807_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X455 a_5565_43396# a_4905_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X456 a_7418_45067# a_7229_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X457 a_1307_43914# a_2779_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X458 a_1793_42852# a_742_44458# a_1709_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X459 VDD a_10227_46804# a_10083_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X460 a_11301_43218# a_10922_42852# a_11229_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X461 VSS a_13291_42460# a_13249_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X462 a_18341_45572# a_18175_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X463 a_19113_45348# a_19321_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X464 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X465 a_8696_44636# a_16855_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X466 a_12189_44484# a_8975_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X467 a_n1736_46482# a_n1853_46287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X468 a_1239_47204# a_1209_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X469 VDD VDAC_Ni a_6886_37412# VSS sky130_fd_pr__nfet_03v3_nvt ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X470 a_n4064_37984# a_n4334_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X471 a_1606_42308# a_1576_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X472 VDD a_n443_42852# a_6481_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X473 VDD a_12005_46116# a_n1741_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X474 a_18315_45260# a_18587_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X475 VSS a_768_44030# a_3600_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X476 VIN_P EN_VIN_BSTR_P a_n1057_35174# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X477 VDD a_4958_30871# a_17531_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X478 a_16795_42852# a_n97_42460# a_16877_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X479 a_18900_46660# a_18834_46812# a_18285_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X480 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X481 a_17973_43940# a_17737_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X482 a_6419_46155# a_5257_43370# a_6347_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X483 a_18597_46090# a_19431_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X484 a_3737_43940# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X485 comp_n a_1169_39043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X486 VDD a_1823_45246# a_4419_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X487 a_22848_40945# COMP_P a_22589_40599# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X488 VDD a_4007_47204# DATA[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X489 VSS a_21496_47436# a_13507_46334# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X490 VSS a_10723_42308# a_5742_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X491 a_22737_36887# a_22527_39145# a_22629_37990# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X492 a_11823_42460# a_15051_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X493 VSS a_n4209_38216# a_n4251_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X494 a_12891_46348# a_4915_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X495 VSS a_20679_44626# a_20640_44752# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X496 a_21115_43940# a_20935_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X497 a_n1821_43396# a_n2267_43396# a_n1917_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X498 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X499 VDD a_10951_45334# a_10775_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X500 a_20850_46155# a_19692_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X501 VDD a_13661_43548# a_18587_45118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X502 a_11649_44734# a_3232_43370# a_n2661_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.174 ps=1.39 w=1 l=0.15
X503 a_20820_30879# a_22591_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X504 VSS a_21359_45002# a_21101_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X505 a_17364_32525# a_22959_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X506 a_18989_43940# a_18451_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X507 a_6197_43396# a_6031_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X508 VDD a_12891_46348# a_13213_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X509 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X510 VREF_GND a_13467_32519# C1_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X511 VDD a_584_46384# a_3540_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X512 a_8873_43396# a_5891_43370# a_8791_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X513 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X514 VSS a_n4334_39392# a_n4064_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X515 C9_P_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X516 a_10809_44484# a_10057_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X517 C6_N_btm a_5742_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X518 a_6545_47178# a_6419_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X519 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X520 a_6109_44484# a_5518_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X521 a_n4318_38216# a_n2472_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X522 VDD a_n901_46420# a_n443_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X523 a_13258_32519# a_19647_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X524 VDD a_11599_46634# a_18819_46122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X525 a_n1435_47204# a_n1605_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X526 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X527 a_15682_43940# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X528 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X529 a_14113_42308# a_13575_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X530 VSS a_4646_46812# a_4651_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X531 a_13381_47204# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X532 VSS a_n2472_46090# a_n2956_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X533 a_4958_30871# a_17124_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X534 VSS a_22223_42860# a_22400_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X535 C0_P_btm a_n3565_37414# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X536 VDD a_1208_46090# a_472_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X537 SMPL_ON_P a_n2002_35608# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X538 VSS a_18479_47436# a_19452_47524# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X539 VSS a_n2302_39072# a_n4209_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X540 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X541 a_n443_46116# a_n901_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X542 a_20623_45572# a_20107_45572# a_20528_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X543 a_12281_43396# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X544 C1_P_btm a_n4209_37414# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X545 VSS a_n3565_39304# a_n3607_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X546 a_15486_42560# a_15764_42576# a_15720_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X547 VSS a_n1613_43370# a_8649_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X548 a_15765_45572# a_15599_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X549 VSS a_n2946_39866# a_n3565_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X550 a_n1613_43370# a_5815_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X551 VSS a_14495_45572# a_n881_46662# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X552 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X553 a_10617_44484# a_10440_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X554 VDD a_5111_44636# a_8487_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X555 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X556 VCM a_5932_42308# C3_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X557 a_20708_46348# a_15227_44166# a_20850_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X558 a_n2267_44484# a_n2433_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X559 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X560 a_1115_44172# a_453_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X561 VSS COMP_P a_n1329_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X562 VSS a_1847_42826# a_2905_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X563 VSS a_15861_45028# a_17023_45118# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X564 a_16292_46812# a_5807_45002# a_16434_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X565 a_17325_44484# a_15227_44166# a_16979_44734# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X566 a_n4064_39072# a_n4334_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X567 a_15803_42450# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X568 a_5534_30871# a_12563_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X569 VSS a_3381_47502# a_3315_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X570 VDD a_9863_46634# a_2063_45854# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X571 VDD a_n2840_43370# a_n4318_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X572 VSS a_584_46384# a_3457_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X573 VIN_N EN_VIN_BSTR_N C3_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X574 a_3863_42891# a_3681_42891# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X575 VDD a_9049_44484# a_9313_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X576 VDD a_376_46348# a_171_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X577 a_11541_44484# a_11453_44696# a_n2661_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X578 VDD a_1431_47204# DATA[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X579 a_19553_46090# a_19335_46494# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X580 a_n1613_43370# a_5815_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X581 a_18727_42674# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X582 a_n1925_42282# a_4185_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X583 VDD a_n2302_37984# a_n4209_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X584 VSS a_17591_47464# a_16327_47482# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X585 VSS a_n3690_38304# a_n3420_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X586 VDD a_19164_43230# a_19339_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X587 a_2479_44172# a_2905_42968# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X588 VSS a_4361_42308# a_21855_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X589 a_n1741_47186# a_12891_46348# a_12839_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X590 VDD a_8103_44636# a_7640_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X591 a_8192_45572# a_8162_45546# a_8120_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X592 a_5009_45028# a_3090_45724# a_4927_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X593 a_12549_44172# a_20567_45036# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X594 VSS a_n2840_42282# a_n3674_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X595 a_5129_47502# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X596 a_14840_46494# a_13759_46122# a_14493_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X597 VSS a_2324_44458# a_949_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X598 VSS a_n913_45002# a_2713_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X599 VDD a_n863_45724# a_1221_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X600 a_8601_46660# a_7411_46660# a_8492_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X601 a_2307_45899# a_n237_47217# a_1848_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X602 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X603 VDD a_n4209_39304# a_n4334_39392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X604 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X605 a_n2946_39072# a_n2956_39304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X606 a_15861_45028# a_15595_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X607 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X608 VSS a_n1613_43370# a_3221_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X609 a_1756_43548# a_768_44030# a_1987_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X610 a_3754_39134# a_7754_39300# VSS sky130_fd_pr__res_high_po_0p35 l=18
X611 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X612 a_n4318_40392# a_n2840_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X613 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X614 VSS a_18143_47464# a_12861_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X615 a_19332_42282# a_19511_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X616 VSS a_17583_46090# a_13259_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X617 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X618 a_20623_43914# a_19321_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X619 VSS a_17499_43370# a_n1059_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X620 VSS a_7754_38470# a_6886_37412# VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X621 a_n3420_39616# a_n3690_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X622 a_4185_45348# a_3065_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X623 a_n2661_46634# a_13017_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X624 VDD a_19321_45002# a_20567_45036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X625 VDD a_6545_47178# a_6575_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X626 VDD a_18285_46348# a_18051_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.16 ps=1.32 w=1 l=0.15
X627 a_2864_46660# a_2747_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X628 VSS a_n809_44244# a_n755_45592# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X629 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X630 VDD a_1307_43914# a_2253_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X631 a_13351_46090# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X632 a_18374_44850# a_18248_44752# a_17970_44736# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X633 a_n913_45002# a_1307_43914# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X634 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X635 a_13657_42308# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X636 a_375_42282# a_413_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X637 a_3090_45724# a_19321_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X638 a_10334_44484# a_10157_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X639 VSS a_10903_43370# a_10057_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X640 a_5700_37509# VSS VDAC_Pi VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X641 a_2113_38308# a_2113_38308# a_2113_38308# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=3.02 ps=24.88 w=1 l=0.15
X642 VSS a_n2438_43548# a_n133_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X643 a_584_46384# a_1123_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X644 VSS a_22959_46124# a_20692_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X645 a_n3674_39768# a_n2472_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X646 VREF a_n4209_39304# C7_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X647 VSS a_20107_42308# a_7174_31319# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X648 a_n4209_39590# a_n2302_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X649 a_526_44458# a_3147_46376# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X650 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X651 a_20301_43646# a_19692_46634# a_20556_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X652 VDD a_n901_46420# a_n914_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X653 a_n971_45724# a_104_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X654 a_20447_31679# a_22959_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X655 VSS a_13348_45260# a_13159_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X656 a_n4334_38304# a_n4318_38216# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X657 VSS a_n881_46662# a_6517_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X658 a_8685_42308# a_8515_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X659 VSS a_6491_46660# a_6851_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X660 a_768_44030# a_13487_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X661 VDD a_14493_46090# a_14383_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X662 a_n327_42308# a_n357_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X663 a_22485_44484# a_22315_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X664 a_15673_47210# a_15507_47210# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X665 SMPL_ON_P a_n2002_35608# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X666 a_8605_42826# a_8387_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X667 a_1709_42852# a_n863_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X668 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X669 VDD a_n1736_42282# a_n4318_37592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X670 VREF a_19721_31679# C2_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X671 VSS a_895_43940# a_2537_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X672 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X673 a_17609_46634# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X674 VDD a_11599_46634# a_18175_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X675 a_8945_43396# a_3537_45260# a_8873_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X676 a_13249_42308# a_10903_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X677 a_601_46902# a_383_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X678 a_4640_45348# a_4574_45260# a_4558_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X679 a_n467_45028# a_n745_45366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X680 a_1208_46090# a_765_45546# a_1337_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X681 VSS a_n1550_35608# a_n2002_35608# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X682 a_3820_44260# a_2382_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X683 VSS a_n863_45724# a_2905_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X684 VSS a_16721_46634# a_16655_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X685 C5_P_btm a_n4064_38528# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X686 a_21588_30879# a_22223_47212# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X687 a_16877_42852# a_16823_43084# a_16795_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X688 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X689 VSS a_17715_44484# a_17737_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X690 a_16241_47178# a_16023_47582# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X691 a_12359_47026# a_11735_46660# a_12251_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X692 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X693 a_5883_43914# a_8333_44056# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X694 a_16759_43396# a_16409_43396# a_16664_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X695 VDD a_n3565_39590# a_n3690_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X696 a_17665_42852# a_17595_43084# a_14539_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X697 VSS a_n2438_43548# a_n2157_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X698 VDD a_4007_47204# DATA[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X699 a_1990_45572# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X700 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X701 a_5072_46660# a_4955_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X702 a_22889_38993# a_22400_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X703 VDD a_3357_43084# a_22591_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X704 VSS a_3815_47204# a_4007_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X705 a_1666_39587# a_1666_39043# a_2112_39137# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X706 a_15803_42450# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X707 a_20528_46660# a_20411_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X708 a_n3607_39392# a_n3674_39304# a_n3690_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X709 VDD a_n4064_39616# a_n2216_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X710 a_21421_42336# a_16327_47482# a_21335_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X711 a_6655_43762# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X712 a_14371_46494# a_13925_46122# a_14275_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X713 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X714 VDD a_3503_45724# a_3218_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X715 VDD a_n2840_43914# a_n4318_39768# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X716 a_15037_43940# a_13556_45296# a_14955_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X717 VSS a_n901_43156# a_n443_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X718 VDD a_10467_46802# a_10428_46928# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X719 a_15060_45348# a_13661_43548# a_14976_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X720 a_9895_44260# a_9290_44172# a_9801_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X721 VDD a_6171_42473# a_5379_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X722 a_5009_45028# a_5147_45002# a_5093_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X723 a_13904_45546# a_10903_43370# a_14127_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X724 a_3537_45260# a_7287_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X725 a_19900_46494# a_18985_46122# a_19553_46090# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X726 VDD a_8696_44636# a_17478_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X727 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X728 a_3935_42891# a_3905_42865# a_3863_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X729 DATA[0] a_327_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X730 VSS a_n881_46662# a_11117_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X731 C3_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X732 VSS a_n4334_39616# a_n4064_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X733 DATA[2] a_4007_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X734 a_15682_46116# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X735 a_1057_46660# a_n133_46660# a_948_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X736 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X737 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X738 VSS a_2982_43646# a_21487_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X739 a_21363_45546# a_21188_45572# a_21542_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X740 VSS a_11823_42460# a_11322_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X741 a_18204_44850# a_17767_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X742 a_n447_43370# a_n2497_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X743 a_17324_43396# a_16409_43396# a_16977_43638# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X744 VSS a_n4064_38528# a_n2302_38778# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X745 a_n443_42852# a_n901_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X746 a_15095_43370# a_15567_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X747 a_10150_46912# a_10428_46928# a_10384_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X748 VSS a_n2472_42282# a_n4318_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X749 a_8492_46660# a_7577_46660# a_8145_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X750 a_5649_42852# a_5111_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X751 VDD a_18287_44626# a_18248_44752# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X752 a_20894_47436# a_20990_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X753 a_19636_46660# a_19594_46812# a_19333_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X754 a_10249_46116# a_9823_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X755 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X756 a_10227_46804# a_14955_47212# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X757 a_739_46482# a_n743_46660# a_376_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X758 VSS a_10775_45002# a_10180_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X759 a_2896_43646# a_2479_44172# a_2982_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X760 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X761 VSS a_n2002_35608# SMPL_ON_P VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X762 a_12791_45546# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X763 VSS a_5807_45002# a_11691_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X764 VDD a_n1794_35242# a_n1696_35090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X765 VSS a_3357_43084# a_22591_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X766 VSS a_2382_45260# a_2304_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X767 a_n4315_30879# a_n2302_40160# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X768 VDD a_n901_46420# a_n443_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X769 a_6298_44484# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X770 a_949_44458# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X771 VDD a_2277_45546# a_2307_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X772 a_10053_45546# a_8746_45002# a_10306_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X773 a_n2956_39768# a_n2840_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X774 VDD a_4361_42308# a_21855_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X775 VDD a_17591_47464# a_16327_47482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X776 VSS a_6945_45028# a_22223_46124# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X777 VDD a_5257_43370# a_5263_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X778 a_n3565_39590# a_n2946_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X779 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X780 VDAC_Ni VSS a_5088_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X781 a_18494_42460# a_18907_42674# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X782 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X783 a_n1151_42308# a_n1329_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X784 a_16763_47508# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X785 a_21259_43561# a_4190_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X786 a_8349_46414# a_8016_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X787 VDD a_1431_47204# DATA[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X788 a_17970_44736# a_18287_44626# a_18245_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X789 a_1123_46634# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X790 a_n237_47217# a_8667_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X791 a_5837_42852# a_3537_45260# a_5755_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X792 VSS a_19692_46634# a_19636_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X793 a_8697_45572# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X794 a_1145_45348# a_n863_45724# a_626_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X795 SMPL_ON_N a_21753_35634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X796 VSS a_5934_30871# a_8515_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X797 VSS a_1239_47204# a_1431_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X798 VSS a_17591_47464# a_16327_47482# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X799 a_11173_44260# a_10729_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X800 VDD a_n4334_38304# a_n4064_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X801 a_22165_42308# a_21887_42336# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X802 a_5244_44056# a_5147_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X803 VSS a_n4064_37440# a_n2302_37690# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X804 VDD a_8952_43230# a_9127_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X805 a_n2956_37592# a_n2472_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X806 VSS a_2127_44172# a_n2661_45010# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X807 VSS a_15493_43940# a_22959_43948# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X808 a_n3565_38502# a_n2946_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X809 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X810 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X811 a_19339_43156# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X812 VDD a_n1920_47178# a_n2312_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X813 VDD a_n1177_44458# a_n1190_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X814 VDD a_16292_46812# a_15811_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X815 a_5164_46348# a_4927_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X816 a_9482_43914# a_9838_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X817 a_20835_44721# a_20679_44626# a_20980_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X818 VSS a_5937_45572# a_8781_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X819 a_19998_35138# VDD EN_VIN_BSTR_N VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.9
X820 a_5837_42852# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X821 a_10037_47542# a_n881_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X822 a_7221_43396# a_6031_43396# a_7112_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X823 VSS a_5937_45572# a_8560_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X824 C7_N_btm a_20820_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X825 VSS a_15559_46634# a_13059_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X826 a_5385_46902# a_5167_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X827 VDD a_10334_44484# a_10440_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X828 a_19597_46482# a_19553_46090# a_19431_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X829 VDD a_n2302_37984# a_n4209_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X830 a_18051_46116# a_18189_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X831 a_15493_43940# a_14955_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X832 a_16414_43172# a_n1059_45260# a_16328_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X833 a_21297_46660# a_20107_46660# a_21188_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X834 a_11813_46116# a_11387_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X835 VSS a_1666_39587# a_1169_39587# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X836 VSS SMPL_ON_P a_n1605_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X837 DATA[4] a_9067_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X838 a_5894_47026# a_4817_46660# a_5732_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X839 VDD a_4699_43561# a_3539_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X840 VSS a_n3420_39072# a_n2946_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X841 VDD a_n97_42460# a_16245_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X842 VDD a_13163_45724# a_11962_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X843 a_15433_44458# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X844 VDD a_16327_47482# a_20980_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X845 a_18114_32519# a_22223_45036# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X846 a_n452_44636# a_n1151_42308# a_n310_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X847 VDD a_22959_43396# a_17364_32525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X848 a_n4064_37984# a_n4334_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X849 VDD a_1307_43914# a_4149_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X850 VSS a_n357_42282# a_7573_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X851 VDD a_9863_47436# a_9804_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X852 a_3754_39134# a_7754_38968# VSS sky130_fd_pr__res_high_po_0p35 l=18
X853 a_4649_43172# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X854 a_526_44458# a_3147_46376# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X855 VSS a_1848_45724# a_1799_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X856 a_22485_38105# a_22775_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X857 a_20885_45572# a_20841_45814# a_20719_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X858 a_10554_47026# a_10428_46928# a_10150_46912# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X859 a_n746_45260# a_n1177_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X860 a_7_44811# a_n1151_42308# a_n452_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X861 VDD a_2324_44458# a_15682_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X862 VDD a_10355_46116# a_8199_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X863 a_4181_43396# a_4093_43548# a_n2661_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X864 VDD a_2437_43646# a_22223_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X865 a_21005_45260# a_21101_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X866 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X867 a_n3565_37414# a_n2946_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X868 a_3754_38802# a_7754_38968# VSS sky130_fd_pr__res_high_po_0p35 l=18
X869 a_2075_43172# a_1307_43914# a_n913_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X870 VSS a_17499_43370# a_n1059_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X871 VSS a_12861_44030# a_17339_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X872 VDD a_n2840_45002# a_n2810_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X873 a_10057_43914# a_10807_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X874 a_5343_44458# a_7963_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X875 a_n1423_42826# a_n1641_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X876 a_526_44458# a_3147_46376# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X877 VDD a_11827_44484# a_22223_45036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X878 VDD a_n2472_43914# a_n3674_39768# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X879 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X880 a_6945_45028# a_5937_45572# a_6945_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X881 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X882 a_20301_43646# a_13661_43548# a_743_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X883 VDD a_n3690_39616# a_n3420_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X884 a_n2216_39866# a_n2442_46660# a_n2302_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X885 VDD a_22000_46634# a_15227_44166# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X886 VSS a_2889_44172# a_413_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X887 VSS a_n97_42460# a_n144_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X888 a_n3674_38216# a_n2104_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X889 a_16321_45348# a_1307_43914# a_16019_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183625 ps=1.215 w=0.65 l=0.15
X890 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X891 VDD a_9290_44172# a_13070_42354# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X892 a_133_42852# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X893 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X894 a_n3420_39072# a_n3690_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X895 a_n2860_38778# a_n2956_38680# a_n2946_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X896 a_22485_38105# a_22775_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X897 a_6517_45366# a_5937_45572# a_6431_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X898 a_10555_44260# a_10729_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X899 VDD a_5111_44636# a_5837_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X900 a_14401_32519# a_22223_43948# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X901 VSS a_9290_44172# a_13070_42354# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X902 VSS a_5068_46348# a_4955_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X903 VDD a_9290_44172# a_10586_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X904 a_16751_45260# a_8696_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X905 a_1666_39587# a_1666_39043# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X906 a_n913_45002# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X907 VSS a_11599_46634# a_15507_47210# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X908 VSS a_768_44030# a_644_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X909 a_12465_44636# a_5807_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X910 VDD a_n357_42282# a_16877_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X911 a_5193_43172# a_3905_42865# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X912 VSS a_18783_43370# a_18525_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X913 a_3540_43646# a_1414_42308# a_3626_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X914 a_21363_45546# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X915 VSS a_n3690_38528# a_n3420_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X916 a_5421_42558# a_5379_42460# a_5337_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X917 VDD a_12861_44030# a_17609_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X918 a_n2956_38216# a_n2472_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X919 a_13885_46660# a_13607_46688# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X920 VCM a_4958_30871# C9_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X921 a_2232_45348# a_1609_45822# a_n2293_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X922 a_5691_45260# a_6171_45002# a_5837_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X923 a_9801_44260# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X924 VCM a_3080_42308# C2_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X925 a_327_44734# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X926 VSS a_7499_43078# a_8746_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X927 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X928 a_15743_43084# a_19339_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X929 VSS a_22591_43396# a_14209_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X930 VSS a_2437_43646# a_22223_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X931 a_6547_43396# a_6197_43396# a_6452_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X932 a_20556_43646# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X933 a_1987_43646# a_742_44458# a_1891_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X934 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X935 a_648_43396# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X936 VDD a_n23_47502# a_7_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X937 a_17609_46634# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X938 a_3602_45348# a_3537_45260# a_3495_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X939 VDD CLK a_8953_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X940 VDD a_2982_43646# a_21487_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X941 a_13661_43548# a_18780_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X942 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X943 a_9313_44734# a_3232_43370# a_9159_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X944 C6_P_btm a_5742_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X945 a_11323_42473# a_5742_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X946 a_14383_46116# a_13759_46122# a_14275_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X947 a_2813_43396# a_2479_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X948 a_16721_46634# a_16388_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X949 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X950 VDD a_526_44458# a_9885_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X951 VSS a_22537_40625# a_22737_36887# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X952 VREF a_20820_30879# C7_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X953 VDD a_15681_43442# a_15781_43660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X954 a_6125_45348# a_3232_43370# a_5691_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X955 VSS a_n1794_35242# a_18194_35068# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X956 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X957 a_10907_45822# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X958 a_14955_43396# a_9145_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X959 a_8128_46384# a_7903_47542# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X960 a_3429_45260# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X961 VDD a_15227_44166# a_17969_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06405 ps=0.725 w=0.42 l=0.15
X962 DATA[0] a_327_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X963 a_n2860_37690# a_n2956_37592# a_n2946_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X964 a_15682_46116# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X965 VSS a_7287_43370# a_3537_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X966 C4_P_btm a_n3420_38528# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X967 a_18599_43230# a_18083_42858# a_18504_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X968 DATA[2] a_4007_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X969 a_18057_42282# a_18494_42460# a_18214_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X970 a_11117_47542# a_4915_47217# a_11031_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X971 a_7112_43396# a_6197_43396# a_6765_43638# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X972 a_584_46384# a_1123_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X973 VSS a_n3690_37440# a_n3420_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X974 VSS a_n901_43156# a_n443_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X975 a_19240_46482# a_19123_46287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X976 VCM a_5742_30871# C6_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X977 VSS a_10193_42453# a_10149_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X978 VDD a_10193_42453# a_10210_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X979 VSS a_2324_44458# a_15682_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X980 VSS a_n967_45348# a_n961_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X981 a_564_42282# a_743_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X982 a_21195_42852# a_20922_43172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X983 VDD a_6575_47204# a_9067_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X984 a_22612_30879# a_22959_47212# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X985 a_21188_46660# a_20273_46660# a_20841_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X986 a_13749_43396# a_13661_43548# a_13667_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X987 VSS a_n2840_45546# a_n2810_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X988 a_13490_45394# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X989 a_n2840_43914# a_n2661_43922# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X990 a_n822_43940# a_n1899_43946# a_n984_44318# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X991 a_21613_42308# a_21335_42336# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X992 a_7112_43396# a_6031_43396# a_6765_43638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X993 a_14537_43396# a_13059_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X994 VDAC_Pi a_3754_38470# a_4338_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X995 a_n4064_39616# a_n4334_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X996 a_n23_47502# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X997 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X998 a_14543_43071# a_5534_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X999 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1000 VDD a_19900_46494# a_20075_46420# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1001 VDD a_7227_45028# a_7230_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1002 VSS a_16327_47482# a_19597_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1003 a_9823_46155# a_n743_46660# a_9751_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1004 VDD a_22959_43948# a_17538_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1005 a_18214_42558# a_16137_43396# a_18057_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1006 a_n3690_38304# a_n3674_38216# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1007 a_15009_46634# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1008 a_17591_47464# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X1009 VSS a_10227_46804# a_15521_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1010 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1011 a_22485_44484# a_22315_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1012 a_n1644_44306# a_n1761_44111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1013 VDD RST_Z a_8530_39574# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1014 VDD a_n1329_42308# a_n1151_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1015 VSS a_13507_46334# a_18184_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1016 a_n630_44306# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1017 a_18783_43370# a_15743_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1018 a_n4064_38528# a_n4334_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1019 a_8325_42308# a_n913_45002# a_8337_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1020 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X1021 a_21973_42336# a_20202_43084# a_21887_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1022 VSS a_n1613_43370# a_645_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1023 a_10341_42308# a_9803_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1024 a_n1920_47178# a_n1741_47186# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1025 VSS a_16327_47482# a_20885_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1026 VSS a_10807_43548# a_11173_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1027 VSS a_5257_43370# a_3905_42865# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1028 a_9127_43156# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1029 VDD a_n2472_45002# a_n2956_37592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1030 VSS a_n2946_39072# a_n3565_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1031 a_13259_45724# a_17583_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1032 VSS a_10586_45546# a_10544_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X1033 a_16751_45260# a_17023_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1034 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1035 VSS a_n4209_38502# a_n4251_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X1036 VSS a_7227_42308# a_6123_31319# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1037 VSS a_10083_42826# a_7499_43078# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1038 a_n2840_42826# a_n2661_42834# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1039 a_1302_46660# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1040 a_5907_45546# a_6194_45824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1041 a_13059_46348# a_15559_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1042 a_n2302_37984# a_n2810_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1043 VREF_GND a_14209_32519# C5_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1044 a_3065_45002# a_3318_42354# a_3581_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X1045 a_16023_47582# a_15673_47210# a_15928_47570# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1046 VSS a_n881_46662# a_n935_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1047 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1048 C6_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1049 VDD a_21487_43396# a_13467_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1050 a_2553_47502# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X1051 VDD a_n443_42852# a_997_45618# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X1052 a_8568_45546# a_8199_44636# a_8791_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1053 a_4338_37500# a_3754_38470# VDAC_Pi VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1054 a_13635_43156# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1055 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1056 VDD a_564_42282# a_n1794_35242# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1057 a_n473_42460# a_n971_45724# a_n327_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X1058 a_16335_44484# a_13661_43548# a_16241_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1059 VDD a_15861_45028# a_17023_45118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1060 a_5205_44734# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1061 a_7499_43078# a_10083_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=2.61 w=1 l=0.15
X1062 VSS a_1123_46634# a_1057_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1063 w_1575_34946# a_n1696_35090# EN_VIN_BSTR_P w_1575_34946# sky130_fd_pr__pfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1064 a_5700_37509# VSS VDAC_Pi VDD sky130_fd_pr__pfet_01v8_hvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1065 a_n4064_37440# a_n4334_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1066 VSS a_13259_45724# a_18315_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1067 a_22737_37285# a_22527_39145# a_22629_38406# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1068 a_n1453_44318# a_n1899_43946# a_n1549_44318# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1069 VSS a_22400_42852# a_22848_40081# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1070 VSS a_22223_43396# a_13887_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1071 a_11682_45822# a_11322_45546# a_11525_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1072 VDD a_22591_45572# a_19963_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1073 a_5934_30871# a_8791_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1074 a_18429_43548# a_18525_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X1075 a_509_45822# a_n1099_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X1076 a_20980_44850# a_20766_44850# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1077 a_4190_30871# a_19332_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1078 a_3381_47502# a_2905_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1079 VDD a_3537_45260# a_4649_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1080 a_6682_46660# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X1081 a_20273_45572# a_20107_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1082 VDD a_11963_45334# a_11787_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X1083 VDD a_1423_45028# a_9838_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1084 a_19256_45572# a_18175_45572# a_18909_45814# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1085 a_n755_45592# a_n809_44244# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1086 VSS a_3699_46634# a_3633_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1087 VSS a_5937_45572# a_9159_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1088 a_14226_46987# a_14180_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X1089 VSS a_n2438_43548# a_n2157_46122# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1090 VSS a_8953_45546# a_9241_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1091 a_n2840_45002# a_n2661_45010# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1092 a_n722_43218# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1093 a_12005_46436# a_2063_45854# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1094 a_9885_43396# a_8270_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1095 VSS a_n4209_37414# a_n4251_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X1096 VDD a_n3690_39616# a_n3420_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X1097 a_18817_42826# a_18599_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1098 EN_VIN_BSTR_P a_n1696_35090# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1099 VDD a_167_45260# a_1423_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1100 VDAC_Pi VSS a_5700_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1101 VSS a_4704_46090# a_1823_45246# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1102 a_16886_45144# a_8696_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X1103 a_11688_45572# a_11652_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X1104 a_8953_45002# CLK VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1105 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1106 a_4520_42826# a_1823_45246# a_4743_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1107 a_949_44458# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1108 a_n3420_39072# a_n3690_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1109 VSS a_22889_38993# a_22944_39857# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1110 VDD a_n2104_42282# a_n3674_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1111 VDD RST_Z a_14311_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1112 a_19721_31679# a_22959_45036# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1113 a_458_43396# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X1114 VSS a_n1696_35090# a_n1057_35174# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1115 a_19339_43156# a_19164_43230# a_19518_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1116 a_11453_44696# a_17719_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1117 VDD a_n3420_37984# a_n2860_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X1118 a_13711_45394# a_12891_46348# a_13348_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X1119 a_16664_43396# a_16547_43609# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1120 a_1138_42852# a_791_42968# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X1121 a_21259_43561# a_4190_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1122 a_10586_45546# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1123 VSS a_11599_46634# a_15599_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1124 VSS a_n3690_38528# a_n3420_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1125 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1126 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X1127 a_196_42282# a_375_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1128 VSS a_n881_46662# a_7989_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1129 a_7832_46660# a_7715_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1130 VDD a_n2109_45247# en_comp VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1131 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1132 a_15928_47570# a_15811_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1133 a_3633_46660# a_2443_46660# a_3524_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1134 VSS a_n2472_45546# a_n2956_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1135 a_2127_44172# a_2675_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X1136 a_9885_43646# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X1137 a_n2472_43914# a_n2293_43922# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1138 VDD a_12991_46634# a_12978_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1139 VDD a_1667_45002# a_n863_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1140 a_n4209_39304# a_n2302_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1141 a_14084_46812# a_n1151_42308# a_14226_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X1142 a_5837_45028# a_3232_43370# a_5691_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X1143 VDD a_21195_42852# a_21671_42860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1144 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1145 a_12427_45724# a_12791_45546# a_12749_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1146 VSS a_n913_45002# a_4921_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1147 a_14209_32519# a_22591_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1148 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1149 a_12553_44484# a_12465_44636# a_n2661_43922# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1150 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1151 a_5829_43940# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1152 a_16237_45028# a_n743_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X1153 VDD a_22959_45036# a_19721_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1154 a_14761_44260# a_14673_44172# a_n2293_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1155 VSS a_n1613_43370# a_5429_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1156 CAL_P a_22485_38105# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1157 VSS a_21363_46634# a_21297_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1158 VDD a_n452_45724# a_n1853_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1159 VDD a_584_46384# a_2998_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1160 VSS a_4699_43561# a_3539_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1161 VDD a_15959_42545# a_15890_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1162 VSS a_10227_46804# a_13157_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1163 a_n4209_38502# a_n2302_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X1164 VSS a_n2946_39866# a_n3565_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1165 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1166 a_17538_32519# a_22959_43948# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1167 a_n144_43396# a_n971_45724# a_n447_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X1168 a_16680_45572# a_15599_45572# a_16333_45814# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1169 VSS a_5937_45572# a_6101_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X1170 a_9672_43914# a_8199_44636# a_9895_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1171 a_15231_43396# a_9145_43396# a_15125_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1172 a_8387_43230# a_7871_42858# a_8292_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1173 VDD a_22731_47423# a_13717_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1174 VDD a_9290_44172# a_13667_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X1175 a_n3420_37984# a_n3690_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X1176 VDD a_10903_43370# a_13163_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.06615 ps=0.735 w=0.42 l=0.15
X1177 VDD a_17767_44458# a_17715_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X1178 VDD a_7845_44172# a_7542_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.28 ps=2.56 w=1 l=0.15
X1179 a_n2840_44458# a_n2661_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1180 a_22400_42852# a_22223_42860# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1181 VDD a_n863_45724# a_945_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X1182 VSS a_9482_43914# a_10157_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1183 VDD a_12549_44172# a_10949_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.195 ps=1.39 w=1 l=0.15
X1184 a_4933_42558# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1185 a_19333_46634# a_19466_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1186 a_13565_44260# a_12891_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1187 VSS a_n3690_37440# a_n3420_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1188 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1189 a_n2293_46098# a_5663_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X1190 VSS a_11453_44696# a_22959_47212# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1191 VSS a_12563_42308# a_5534_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1192 a_n2472_42826# a_n2293_42834# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1193 a_7920_46348# a_8128_46384# a_8062_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1194 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1195 a_n13_43084# a_n443_42852# a_133_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1196 a_2698_46116# a_2521_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1197 a_15785_43172# a_15743_43084# a_15095_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X1198 a_8654_47026# a_7577_46660# a_8492_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1199 VDD a_21363_46634# a_21350_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1200 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1201 VDD a_n809_44244# a_n822_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1202 a_766_43646# a_626_44172# a_458_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X1203 a_n784_42308# a_n961_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1204 a_12895_43230# a_12379_42858# a_12800_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1205 VSS a_805_46414# a_739_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1206 VSS a_8191_45002# a_8137_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1207 a_15959_42545# a_15803_42450# a_16104_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1208 a_5210_46482# a_5164_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X1209 a_11341_43940# a_3232_43370# a_11173_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.19825 ps=1.26 w=0.65 l=0.15
X1210 VDD a_7705_45326# a_7735_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1211 a_13720_44458# a_13661_43548# a_13940_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1212 a_2162_46660# a_2107_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X1213 VSS a_n4334_39392# a_n4064_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1214 a_n1423_42826# a_n1641_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1215 a_n2956_39304# a_n2840_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1216 VDD a_11415_45002# a_n2661_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1217 a_15037_43940# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X1218 VDD a_1606_42308# a_2351_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1219 a_2277_45546# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1220 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1221 a_6903_46660# a_6755_46942# a_6540_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X1222 VDD a_14180_45002# a_13017_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1223 a_3232_43370# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1224 VDD a_n2302_40160# a_n4315_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1225 VDD a_8199_44636# a_8191_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X1226 a_n4209_37414# a_n2302_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X1227 a_1576_42282# a_1755_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1228 a_7573_43172# a_7499_43078# a_7227_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1229 VSS a_21855_43396# a_13678_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1230 VDD a_18989_43940# a_19006_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1231 VSS a_6540_46812# a_6491_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1232 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1233 VDD a_22223_45572# a_19479_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1234 VIN_N EN_VIN_BSTR_N C0_dummy_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1235 VSS a_2903_42308# a_3080_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1236 VSS a_n863_45724# a_n906_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X1237 a_n2840_44458# a_n2661_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1238 a_22629_37990# a_22581_37893# CAL_P VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1239 a_3823_42558# a_3065_45002# a_3905_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1240 VSS a_2779_44458# a_1307_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X1241 VSS a_5263_45724# a_5204_45822# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1242 VDD a_2124_47436# a_1209_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1243 a_12925_46660# a_11735_46660# a_12816_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1244 VSS a_2957_45546# a_2905_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1245 a_376_46348# a_n743_46660# a_518_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X1246 a_11415_45002# a_4915_47217# a_14581_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1247 VDD a_7754_40130# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.5
X1248 a_n2104_42282# a_n1925_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1249 a_n2472_45002# a_n2293_45010# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1250 a_21398_44850# a_20679_44626# a_20835_44721# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1251 VDD a_16333_45814# a_16223_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1252 a_16241_44484# a_2711_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1253 a_3905_42865# a_5257_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1254 VSS a_8685_43396# a_15231_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1255 VSS a_10623_46897# a_10554_47026# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1256 a_13485_45572# a_12549_44172# a_13385_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X1257 C3_P_btm a_n4209_38216# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1258 VSS a_22959_45572# a_20447_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1259 a_22848_39857# a_22485_38105# a_22581_37893# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1260 VDD a_19987_42826# a_n2017_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.135 ps=1.27 w=1 l=0.15
X1261 a_9028_43914# a_9482_43914# a_9420_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X1262 VSS a_17973_43940# a_18079_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X1263 a_n2860_39072# a_n2956_39304# a_n2946_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X1264 a_9290_44172# a_13635_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1265 a_3059_42968# a_742_44458# a_2987_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1266 a_n452_44636# a_n467_45028# a_n310_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X1267 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1268 VDD a_768_44030# a_2711_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1269 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1270 VDD a_12281_43396# a_12563_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1271 VDD a_12741_44636# a_22959_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1272 a_8333_44734# a_3537_45260# a_8238_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X1273 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1274 a_17124_42282# a_17303_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1275 a_12156_46660# a_11813_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1276 VDD a_10809_44734# a_22959_46124# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1277 VSS a_1115_44172# a_n2293_45010# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X1278 a_5013_44260# a_1307_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1279 VDD a_n447_43370# a_n2129_43609# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1280 a_3357_43084# a_5257_43370# a_5565_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1281 a_1568_43370# a_1847_42826# a_1793_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1282 a_n967_43230# a_n2157_42858# a_n1076_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1283 a_11682_45822# a_10586_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X1284 a_18315_45260# a_15227_44166# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X1285 a_n2012_44484# a_n2129_44697# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1286 a_14543_43071# a_5534_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1287 a_16147_45260# a_17478_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1288 a_22848_40081# en_comp a_22589_40055# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1289 a_19963_31679# a_22591_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1290 a_n967_45348# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1291 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1292 VDD a_11599_46634# a_20107_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1293 VSS a_7276_45260# a_7227_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1294 a_1241_44260# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.102375 ps=0.965 w=0.65 l=0.15
X1295 VDD a_n809_44244# a_n755_45592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1296 VSS a_n815_47178# a_n785_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1297 a_n4334_40480# a_n4318_40392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1298 a_3175_45822# a_3090_45724# a_2957_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X1299 a_14621_43646# a_14579_43548# a_14537_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1300 VDD a_n2946_37984# a_n3565_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1301 VREF a_20205_31679# C4_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1302 VSS a_15227_44166# a_18900_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X1303 a_n310_44811# a_n356_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X1304 VDD a_16977_43638# a_16867_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1305 VDD a_15227_44166# a_17749_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X1306 a_3147_46376# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X1307 a_12638_46436# a_12594_46348# a_12379_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1308 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1309 VSS a_2324_44458# a_6298_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1310 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1311 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1312 a_21071_46482# a_15227_44166# a_20708_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X1313 a_n1059_45260# a_17499_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1314 VDD a_1273_38525# a_2684_37794# VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1315 a_961_42354# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1316 a_9127_43156# a_8952_43230# a_9306_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1317 VSS a_12741_44636# a_22959_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1318 VSS a_8349_46414# a_8283_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1319 VSS a_11787_45002# a_11652_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X1320 a_4223_44672# a_3537_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1321 a_509_45822# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1322 a_16119_47582# a_15673_47210# a_16023_47582# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1323 a_6452_43396# a_6293_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1324 VSS CLK a_8953_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1325 a_6194_45824# a_6472_45840# a_6428_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1326 a_3754_38802# a_7754_38636# VSS sky130_fd_pr__res_high_po_0p35 l=18
X1327 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1328 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1329 VDD a_n881_46662# a_11031_47542# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1330 VSS a_1209_47178# a_1239_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1331 a_n217_35174# a_n1696_35090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1332 a_15559_46634# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X1333 a_12429_44172# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1334 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1335 a_11229_43218# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1336 a_16020_45572# a_15903_45785# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1337 C3_P_btm a_5932_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1338 a_10149_42308# a_9290_44172# a_9803_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1339 VSS a_20708_46348# a_20411_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1340 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1341 C9_N_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1342 a_10793_43218# a_10083_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1343 a_n863_45724# a_1667_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1344 a_13635_43156# a_13460_43230# a_13814_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1345 a_12379_46436# a_12594_46348# a_12638_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1346 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1347 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1348 a_1209_43370# a_1049_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1349 a_2982_43646# a_3232_43370# a_2813_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1350 a_n443_46116# a_n901_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1351 a_21542_45572# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1352 VSS a_19647_42308# a_13258_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1353 a_18985_46122# a_18819_46122# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1354 a_12839_46116# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1355 VDD a_n2438_43548# a_2443_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1356 VDD a_9028_43914# a_8975_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1357 VDD a_17124_42282# a_4958_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1358 VSS a_10053_45546# a_9625_46129# VSS sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X1359 a_17639_46660# a_17609_46634# a_765_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1360 VSS a_380_45546# a_n356_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X1361 VSS a_n2002_35608# SMPL_ON_P VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1362 VSS a_20193_45348# a_21973_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1363 VSS a_196_42282# a_n3674_37592# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1364 VDD a_n1794_35242# a_n1696_35090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1365 VDD a_5257_43370# a_5826_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X1366 a_9803_42558# a_n97_42460# a_9885_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1367 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1368 VSS a_10227_46804# a_10553_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1369 VSS a_18597_46090# a_16375_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1370 VSS a_n913_45002# a_12281_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1371 a_12816_46660# a_11901_46660# a_12469_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1372 a_n3565_39590# a_n2946_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1373 a_20205_45028# a_18184_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1374 a_n3420_37984# a_n3690_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1375 VDD a_13259_45724# a_13667_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1376 a_n1736_42282# a_n1557_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1377 a_13747_46662# a_19386_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1378 VSS a_4791_45118# a_6165_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X1379 a_261_44278# a_n863_45724# a_175_44278# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1380 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1381 a_8325_42308# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1382 a_10623_46897# a_10467_46802# a_10768_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1383 a_17957_46116# a_765_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.208 ps=1.94 w=0.65 l=0.15
X1384 a_2675_43914# a_2998_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1385 a_18695_43230# a_18249_42858# a_18599_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1386 a_17613_45144# a_8696_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1387 a_n4318_39304# a_n2840_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1388 a_18799_45938# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1389 VSS a_19862_44208# a_20922_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.089375 ps=0.925 w=0.65 l=0.15
X1390 a_6151_47436# a_14311_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1391 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1392 VSS a_5129_47502# a_5063_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1393 VSS a_167_45260# a_2521_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1394 a_3733_45822# a_n755_45592# a_3638_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X1395 a_16333_45814# a_16115_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1396 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1397 a_1337_46116# a_1176_45822# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X1398 a_13163_45724# a_13527_45546# a_13485_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1399 a_8605_42826# a_8387_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1400 VDD a_4419_46090# a_n1925_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1401 a_n4209_38216# a_n2302_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1402 a_20712_42282# a_n357_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1403 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1404 a_1241_43940# a_1467_44172# a_1443_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1405 a_9145_43396# a_8791_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1406 VDD a_n961_42308# a_n784_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1407 a_7227_42852# a_n97_42460# a_7309_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1408 a_14976_45348# a_13059_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X1409 a_9863_47436# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X1410 a_743_42282# a_19692_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1411 a_4915_47217# a_12991_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1412 VSS a_12891_46348# a_12638_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1413 a_n3674_38680# a_n2840_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1414 VCM a_4958_30871# C9_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1415 VSS a_3539_42460# a_3065_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1416 a_17801_45144# a_17613_45144# a_17719_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X1417 VDD a_n4209_39590# a_n4334_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X1418 a_18787_45572# a_18341_45572# a_18691_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1419 a_10922_42852# a_10796_42968# a_10518_42984# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1420 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1421 a_3754_39964# a_7754_40130# VSS sky130_fd_pr__res_high_po_0p35 l=18
X1422 VDD a_n4334_40480# a_n4064_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1423 VDD a_526_44458# a_3232_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1424 a_n1794_35242# a_564_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1425 a_167_45260# a_2202_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1426 VDD a_11967_42832# a_20512_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1427 VDD a_16019_45002# a_15903_45785# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1428 a_2896_43646# a_n443_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1429 VSS a_9067_47204# DATA[4] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1430 a_n2312_38680# a_n2104_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1431 a_12005_46116# a_10903_43370# a_12005_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1432 a_n2288_47178# a_n2109_47186# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1433 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1434 a_14097_32519# a_22959_42860# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1435 a_6999_46987# a_3877_44458# a_6540_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1436 a_8199_44636# a_10355_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X1437 a_3429_45260# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1438 a_n217_35174# VDD EN_VIN_BSTR_P VSS sky130_fd_pr__nfet_05v0_nvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.9
X1439 C8_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1440 a_4338_37500# VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.589 ps=4.42 w=1.9 l=0.15
X1441 a_9293_42558# a_9223_42460# a_8953_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X1442 VDD a_n452_47436# a_n815_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1443 VDD a_n2302_40160# a_n4315_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1444 a_14309_45348# a_2711_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1445 a_13807_45067# a_13556_45296# a_13348_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1446 a_2981_46116# a_2804_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1447 a_1176_45822# a_997_45618# a_1260_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X1448 a_4185_45028# a_3877_44458# a_4185_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1449 VDD a_13159_45002# a_n2661_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1450 VSS a_20269_44172# a_19319_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1451 a_n1655_43396# a_n1699_43638# a_n1821_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1452 a_16104_42674# a_15890_42674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1453 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1454 a_22731_47423# SMPL_ON_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1455 a_n722_46482# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1456 VSS a_n443_42852# a_997_45618# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1457 a_6945_45348# a_5205_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1458 a_21513_45002# a_21363_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1459 a_4791_45118# a_4743_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X1460 VSS a_1576_42282# a_1606_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1461 a_n1533_46116# a_n2157_46122# a_n1641_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1462 a_15227_44166# a_22000_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1463 a_n743_46660# a_n1021_46688# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1464 a_n4064_40160# a_n4334_40480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X1465 a_2075_43172# a_1307_43914# a_n913_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1466 VSS a_5205_44484# a_6756_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1467 VDD a_327_44734# a_375_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1468 VDD a_19321_45002# a_3090_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X1469 VSS a_3483_46348# a_13829_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X1470 VDD a_7754_40130# a_11206_38545# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X1471 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1472 VDD a_5937_45572# a_6671_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1473 VDD a_n863_45724# a_458_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X1474 VDD a_n4334_38304# a_n4064_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X1475 VDD a_526_44458# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1476 VDD a_1756_43548# a_1467_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.28 ps=2.56 w=1 l=0.15
X1477 VDD a_4791_45118# a_5066_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1478 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1479 a_20269_44172# a_20365_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X1480 VDD a_14976_45028# a_15227_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1481 VSS a_13904_45546# a_12594_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X1482 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1483 VSS a_8953_45546# a_8568_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X1484 VDAC_Pi a_3754_38470# a_4338_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1485 a_16112_44458# a_15227_44166# a_16335_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1486 VSS a_16327_47482# a_17021_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1487 a_n913_45002# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1488 VSS a_20974_43370# a_20749_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1489 a_16388_46812# a_17957_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1725 ps=1.345 w=1 l=0.15
X1490 VSS a_20159_44458# a_19321_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X1491 VDD a_9672_43914# a_2107_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1492 VSS a_22589_40599# a_22737_37285# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1493 a_n4318_37592# a_n1736_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1494 VSS a_6151_47436# a_8189_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1495 VDD a_12549_44172# a_17609_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1496 a_6229_45572# a_6194_45824# a_5907_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1497 VDD a_19700_43370# a_n97_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1498 a_6851_47204# a_6491_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1499 a_n2002_35608# a_n1550_35608# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1500 VDD a_19615_44636# a_18579_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X1501 a_8423_43396# a_n443_42852# a_8317_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1502 VDD a_7499_43078# a_8697_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1503 a_18799_45938# a_18175_45572# a_18691_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1504 a_1755_42282# a_n913_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1505 a_n1741_47186# a_12005_46116# a_12379_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X1506 VSS a_2324_44458# a_6298_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1507 VDD a_6765_43638# a_6655_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1508 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1509 a_n4209_39304# a_n2302_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X1510 VDD a_22223_47212# a_21588_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1511 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1512 a_685_42968# a_n443_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1513 a_10467_46802# a_11599_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1514 VDD a_n443_42852# a_15781_43660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X1515 a_17749_42852# a_17701_42308# a_17665_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1516 a_18599_43230# a_18249_42858# a_18504_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1517 CLK_DATA a_n2833_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X1518 VDD a_7920_46348# a_7715_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1519 a_3537_45260# a_7287_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1520 a_2809_45028# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X1521 a_7832_46660# a_7715_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1522 a_3873_46454# a_n881_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X1523 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1524 VSS a_4905_42826# a_4520_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X1525 a_6709_45028# a_6431_45366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1526 VSS a_20202_43084# a_21421_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1527 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1528 a_20623_43914# a_19321_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1529 a_20193_45348# a_18494_42460# a_20205_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1530 VSS a_9313_45822# a_11459_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X1531 a_n4318_39768# a_n2840_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1532 a_n443_42852# a_n901_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1533 a_6428_45938# a_5907_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1534 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1535 a_1273_38525# a_1107_38525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1536 a_n2104_46634# a_n1925_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1537 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1538 VSS a_7287_43370# a_3537_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1539 a_2987_42968# a_1847_42826# a_2905_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1540 a_11031_47542# a_4915_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1541 VSS a_12991_46634# a_12925_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1542 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1543 VDAC_Ni a_7754_38636# VSS sky130_fd_pr__res_high_po_0p35 l=18
X1544 VSS a_20894_47436# a_20843_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1545 a_13076_44458# a_9482_43914# a_13468_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X1546 a_10752_42852# a_10083_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1547 a_n1809_43762# a_n2433_43396# a_n1917_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1548 a_17970_44736# a_18248_44752# a_18204_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1549 a_5663_43940# a_5883_43914# a_5841_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X1550 a_n2302_38778# a_n2312_38680# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1551 a_16588_47582# a_15507_47210# a_16241_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1552 VSS a_4099_45572# a_3483_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1553 VSS a_14539_43914# a_16112_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X1554 a_16867_43762# a_16243_43396# a_16759_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1555 VDD a_1107_38525# a_1273_38525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1556 a_n745_45366# a_n746_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1557 a_10518_42984# a_10835_43094# a_10793_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1558 C2_P_btm a_n3420_37984# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1559 VIN_P EN_VIN_BSTR_P C5_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1560 a_n37_45144# a_n443_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1561 a_18287_44626# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1562 a_20159_44458# a_20362_44736# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1563 VSS a_11341_43940# a_22223_43948# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1564 VSS a_8530_39574# a_3754_38470# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1565 DATA[5] a_11459_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1566 a_6969_46634# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1567 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1568 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1569 a_18861_43218# a_18817_42826# a_18695_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1570 a_11322_45546# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1571 a_n3674_37592# a_196_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1572 a_n1809_43762# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1573 a_n1696_35090# a_n1794_35242# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1574 a_4419_46090# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X1575 VDD a_11189_46129# a_11133_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X1576 VDD a_7227_47204# DATA[3] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1577 a_n1076_46494# a_n1991_46122# a_n1423_46090# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1578 VSS a_7640_43914# a_7584_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1579 a_15959_42545# a_15764_42576# a_16269_42308# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1580 a_16375_45002# a_18597_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1581 VDD a_n1699_44726# a_n1809_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1582 a_4235_43370# a_3935_42891# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X1583 a_21177_47436# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X1584 a_7418_45394# a_7229_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X1585 a_22000_46634# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1586 VDD a_7542_44172# a_7499_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1587 SMPL_ON_N a_21753_35634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1588 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1589 a_11309_47204# a_11031_47542# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1590 VDD a_1307_43914# a_3353_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1591 a_3905_42308# a_2382_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1592 a_8483_43230# a_8037_42858# a_8387_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1593 a_n2104_46634# a_n1925_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1594 a_453_43940# a_175_44278# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1595 a_7281_43914# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1596 a_9028_43914# a_9290_44172# a_9248_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1597 VDD a_n2302_38778# a_n4209_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1598 VDD a_4700_47436# a_3785_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1599 a_18909_45814# a_18691_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1600 a_15521_42308# a_15486_42560# a_15051_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1601 a_11551_42558# a_n97_42460# a_11633_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1602 VSS a_11459_47204# DATA[5] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1603 VDD a_15227_44166# a_15415_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X1604 VSS a_16327_47482# a_20397_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1605 a_n809_44244# a_n984_44318# a_n630_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1606 VDD a_8270_45546# a_9165_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1607 VDD a_948_46660# a_1123_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1608 VDD a_15009_46634# a_14180_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1609 a_20766_44850# a_20679_44626# a_20362_44736# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1610 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1611 a_13385_45572# a_10903_43370# a_13297_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X1612 VDD a_13777_45326# a_13807_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1613 VSS a_21753_35634# SMPL_ON_N VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1614 VSS a_n755_45592# a_n39_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1615 a_14976_45028# a_14797_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X1616 VSS a_22589_40599# a_22537_40625# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1617 a_6886_37412# VDAC_Pi VDD VSS sky130_fd_pr__nfet_03v3_nvt ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X1618 a_6419_46482# a_6165_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X1619 VSS a_768_44030# a_5244_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1620 a_n2302_37690# a_n2810_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1621 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1622 VSS a_n2946_39072# a_n3565_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1623 VDD a_8199_44636# a_8336_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X1624 a_20623_45572# a_20273_45572# a_20528_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1625 VSS a_9396_43370# a_5111_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1626 a_n2312_39304# a_n1920_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1627 a_20009_46494# a_18819_46122# a_19900_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1628 a_n1190_44850# a_n2267_44484# a_n1352_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1629 a_7309_42852# a_5891_43370# a_7227_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1630 a_743_42282# a_13661_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1631 VSS a_n4064_40160# a_n2302_40160# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X1632 a_22397_42558# a_n913_45002# a_17303_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1633 a_12991_43230# a_12545_42858# a_12895_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1634 VSS a_3905_42865# a_5013_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1635 VDD a_21753_35634# SMPL_ON_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1636 a_22765_42852# a_15743_43084# a_18184_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1637 a_7705_45326# a_7229_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1638 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1639 VSS a_10405_44172# a_8016_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1640 a_3065_45002# a_1823_45246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X1641 a_742_44458# a_n443_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1642 a_310_45028# a_n37_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1643 VDD a_3232_43370# a_2982_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1644 VDD a_526_44458# a_3905_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1645 VSS a_18184_42460# a_20256_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.11375 ps=1 w=0.65 l=0.15
X1646 VDD a_16241_47178# a_16131_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1647 a_19466_46812# a_13747_46662# a_19929_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1648 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1649 a_20850_46482# a_19692_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X1650 VSS a_768_44030# a_9028_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X1651 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1652 a_12089_42308# a_11551_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1653 a_11173_43940# a_2063_45854# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1654 a_3457_43396# a_1414_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1655 VDD a_5907_46634# a_5894_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1656 a_8034_45724# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1657 a_5841_46660# a_4651_46660# a_5732_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1658 a_22000_46634# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1659 VSS a_3699_46348# a_3160_47472# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1660 VSS a_22223_45036# a_18114_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1661 a_2437_43396# a_1568_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1662 VDD a_n2104_46634# a_n2312_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1663 a_2448_45028# a_2382_45260# a_n2293_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X1664 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1665 a_21167_46155# a_20916_46384# a_20708_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1666 a_22725_37990# a_22589_40055# a_22629_37990# VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1667 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1668 a_5205_44484# a_5343_44458# a_5289_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1669 a_7499_43078# a_10083_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1670 a_948_46660# a_33_46660# a_601_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1671 VSS a_21005_45260# a_19778_44110# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1672 VDD a_n2302_37690# a_n4209_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1673 VSS a_13487_47204# a_768_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X1674 a_9241_46436# a_n237_47217# a_8049_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1675 a_15015_46420# a_14840_46494# a_15194_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1676 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1677 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1678 VDD a_20567_45036# a_12549_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1679 a_21398_44850# a_20640_44752# a_20835_44721# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1680 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1681 a_1823_45246# a_4704_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1682 a_5527_46155# a_5204_45822# a_5068_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1683 a_1606_42308# a_1576_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1684 VSS a_4235_43370# a_4181_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1685 VDD a_18783_43370# a_18525_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X1686 a_n881_46662# a_14495_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X1687 a_21188_45572# a_20107_45572# a_20841_45814# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1688 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1689 a_n1821_44484# a_n2267_44484# a_n1917_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1690 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1691 a_22944_39857# a_22613_38993# a_22848_39857# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1692 VCM a_5534_30871# C7_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X1693 VSS a_8270_45546# a_8192_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X1694 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1695 a_5891_43370# a_9127_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1696 VDD a_n863_45724# a_3059_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1697 VDD a_17609_46634# a_765_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1698 VSS a_n755_45592# a_3503_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1699 a_19237_31679# a_22959_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1700 a_12156_46660# a_11813_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1701 a_n4334_38528# a_n4318_38680# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1702 a_n901_43156# a_n1076_43230# a_n722_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1703 a_n2810_45028# a_n2840_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1704 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1705 a_16333_45814# a_16115_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1706 a_16795_42852# a_n97_42460# a_16877_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1707 a_n913_45002# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1708 VDD a_21188_46660# a_21363_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1709 a_6905_45572# a_6151_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1710 a_14180_45002# a_13059_46348# a_14403_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1711 a_16405_45348# a_16375_45002# a_16321_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1712 VDD a_5934_30871# a_8515_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1713 w_1575_34946# a_n1057_35174# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=10.615 ps=76.96 w=3.75 l=15
X1714 VREF a_19963_31679# C3_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1715 VDD a_3422_30871# a_22315_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1716 a_2123_42473# a_n784_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1717 VSS a_n1613_43370# a_n1287_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1718 VSS a_22223_43948# a_14401_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1719 a_19518_43218# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1720 VSS a_20075_46420# a_20009_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1721 VSS a_16922_45042# a_16751_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1722 VDD a_3232_43370# a_11341_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.3925 ps=1.785 w=1 l=0.15
X1723 a_1049_43396# a_458_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1724 VDD a_1169_39587# COMP_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1725 VDD a_526_44458# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1726 VDD a_n237_47217# a_8270_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1727 a_1848_45724# a_n237_47217# a_1990_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1728 VDD a_14539_43914# a_12465_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1729 VDD a_n881_46662# a_7903_47542# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1730 VDD a_1666_39043# a_1169_39043# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1731 VDD a_n1423_46090# a_n1533_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1732 VDD a_5111_44636# a_5421_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X1733 a_20623_46660# a_20107_46660# a_20528_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1734 a_11778_45572# a_10193_42453# a_11688_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X1735 a_6347_46155# a_6165_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1736 a_4700_47436# a_n443_46116# a_4842_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1737 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1738 VDD a_21359_45002# a_21101_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X1739 C4_P_btm a_n3565_38502# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1740 a_14113_42308# a_13575_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1741 VDD a_5755_42308# a_5932_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1742 a_10695_43548# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1743 a_4958_30871# a_17124_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1744 a_17333_42852# a_16795_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1745 VSS a_19339_43156# a_19273_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1746 a_8387_43230# a_8037_42858# a_8292_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1747 VDD a_n2840_44458# a_n4318_40392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1748 VDD a_15004_44636# a_14815_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1749 VSS a_16327_47482# a_18861_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1750 VSS a_1823_45246# a_3602_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X1751 VDD a_18780_47178# a_13661_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1752 a_n4334_37440# a_n4318_37592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1753 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1754 a_2455_43940# a_895_43940# a_2253_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1755 a_2680_45002# a_3065_45002# a_2809_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1756 a_13667_43396# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X1757 a_21381_43940# a_21115_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1758 a_380_45546# a_765_45546# a_509_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1759 a_15781_43660# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X1760 a_16019_45002# a_16147_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.183625 pd=1.215 as=0.160875 ps=1.145 w=0.65 l=0.15
X1761 VDD a_3537_45260# a_4558_45348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X1762 a_12741_44636# a_6755_46942# a_16789_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1763 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1764 a_5534_30871# a_12563_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1765 VSS a_2324_44458# a_15682_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1766 VDD en_comp a_1107_38525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1767 VDD a_n473_42460# a_n1761_44111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X1768 VSS a_7754_38470# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0 ps=0 w=2 l=0.15
X1769 a_20836_43172# a_20193_45348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1770 a_12895_43230# a_12545_42858# a_12800_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1771 VSS a_n2833_47464# CLK_DATA VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1772 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X1773 VDD a_1123_46634# a_584_46384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1774 a_726_44056# a_626_44172# a_644_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1775 a_6655_43762# a_6031_43396# a_6547_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1776 DATA[5] a_11459_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X1777 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1778 a_2889_44172# a_1414_42308# a_3052_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1779 VDD a_3232_43370# a_3626_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1780 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1781 a_5343_44458# a_7963_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1782 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1783 a_3483_46348# a_4099_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1784 a_9313_44734# a_5883_43914# a_9241_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1785 a_2809_45028# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1786 VDD a_6171_45002# a_11827_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1787 VDD a_9625_46129# a_9569_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X1788 a_15567_42826# a_15227_44166# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1789 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X1790 a_2113_38308# a_2113_38308# a_2113_38308# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1791 a_7_45899# a_n443_46116# a_n452_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1792 a_n2810_45572# a_n2840_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1793 a_5732_46660# a_4817_46660# a_5385_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1794 a_5708_44484# a_3483_46348# a_5608_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X1795 VDD a_13259_45724# a_22397_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1796 a_11823_42460# a_15051_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=2.61 w=1 l=0.15
X1797 VDD a_13507_46334# a_22765_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1798 a_13678_32519# a_21855_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1799 a_5365_45348# a_5111_44636# a_4927_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1800 a_17021_43396# a_16977_43638# a_16855_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1801 VDD a_7227_47204# DATA[3] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1802 VREF_GND a_n4064_39616# C9_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1803 a_7989_47542# a_n237_47217# a_7903_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1804 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1805 a_19332_42282# a_19511_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1806 VSS a_6851_47204# a_7227_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X1807 a_13607_46688# a_6755_46942# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1808 a_4880_45572# a_526_44458# a_4808_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X1809 EN_VIN_BSTR_N a_18194_35068# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1810 a_20922_43172# a_10193_42453# a_20836_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X1811 a_12978_47026# a_11901_46660# a_12816_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1812 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1813 VDD a_13720_44458# a_12607_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1814 VDD a_2952_47436# a_2747_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1815 a_5147_45002# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1816 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1817 VDD a_14513_46634# a_14543_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1818 VDD a_21259_43561# a_16922_45042# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1819 VDD a_n4334_38528# a_n4064_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1820 VSS a_11459_47204# DATA[5] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1821 VDD a_21137_46414# a_21167_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1822 C9_N_btm a_17730_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1823 a_3905_42558# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X1824 VSS a_22959_47212# a_22612_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1825 a_383_46660# a_33_46660# a_288_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1826 VSS a_6755_46942# a_13556_45296# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1827 a_n4209_38216# a_n2302_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X1828 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1829 a_17061_44734# a_11691_44458# a_16979_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1830 a_4149_42891# a_2382_45260# a_3935_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X1831 DATA[3] a_7227_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1832 VDD a_n755_45592# a_3318_42354# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X1833 VDD a_n443_46116# a_1427_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1834 VDD a_5497_46414# a_5527_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1835 a_5937_45572# a_5907_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1836 a_11323_42473# a_5742_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1837 VSS a_4921_42308# a_5755_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1838 a_21076_30879# a_22959_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1839 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1840 VDD a_n2302_38778# a_n4209_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1841 a_n3565_39304# a_n2946_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1842 a_3699_46634# a_3524_46660# a_3878_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1843 VDD a_17583_46090# a_13259_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1844 VSS a_3600_43914# a_3499_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X1845 VSS a_n755_45592# a_3318_42354# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1846 a_5111_44636# a_9396_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1847 a_17595_43084# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1848 a_13829_44260# a_13059_46348# a_13483_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1849 a_18341_45572# a_18175_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1850 a_9290_44172# a_13635_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1851 a_12991_46634# a_12816_46660# a_13170_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1852 VSS a_2277_45546# a_2211_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1853 a_18429_43548# a_18525_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X1854 VSS a_6453_43914# a_n2661_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1855 a_6773_42558# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1856 a_2253_44260# a_n443_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.102375 ps=0.965 w=0.65 l=0.15
X1857 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1858 a_9885_42558# a_7499_43078# a_9803_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1859 a_16414_43172# a_16137_43396# a_16245_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X1860 a_21811_47423# SINGLE_ENDED VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1861 a_2304_45348# a_n863_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X1862 a_3726_37500# a_6886_37412# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=0.15
X1863 a_13351_46090# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X1864 a_n4064_38528# a_n4334_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X1865 a_n1435_47204# a_n1605_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1866 a_n935_46688# a_n1151_42308# a_n1021_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1867 VSS a_12549_44172# a_17639_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.099125 ps=0.955 w=0.65 l=0.15
X1868 a_6977_45572# a_6598_45938# a_6905_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1869 VSS a_n23_44458# a_n89_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1870 VSS a_n1177_43370# a_n1243_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1871 VDD a_13460_43230# a_13635_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1872 VSS a_n913_45002# a_n967_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1873 VDD a_11525_45546# a_11189_46129# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X1874 VDD a_n755_45592# a_626_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1875 a_n1287_44306# a_n1331_43914# a_n1453_44318# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1876 VDD a_10227_46804# a_10768_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1877 a_n755_45592# a_n809_44244# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1878 a_895_43940# a_644_44056# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X1879 a_n699_43396# a_n1177_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1880 a_11136_42852# a_10922_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1881 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1882 VDD a_8568_45546# a_8162_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1883 VDD a_n4334_37440# a_n4064_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1884 a_11551_42558# a_n97_42460# a_11633_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1885 a_6293_42852# a_5755_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1886 a_n2840_42826# a_n2661_42834# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1887 a_16131_47204# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1888 a_14033_45572# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1889 a_5289_44734# a_4223_44672# a_5205_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1890 VSS a_n1736_42282# a_n4318_37592# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1891 VDD a_10083_42826# a_7499_43078# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1892 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1893 a_768_44030# a_13487_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1894 VDD a_11415_45002# a_22591_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1895 VSS a_5147_45002# a_5708_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X1896 VIN_N EN_VIN_BSTR_N C8_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1897 VDD a_13259_45724# a_14309_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1898 VSS a_6886_37412# a_4338_37500# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=0.15
X1899 a_10053_45546# a_10490_45724# a_10210_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X1900 a_n4064_40160# a_n4334_40480# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1901 VDD a_19332_42282# a_4190_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1902 a_n998_43396# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1903 a_3090_45724# a_18911_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1468 ps=1.34 w=1 l=0.15
X1904 VSS a_18287_44626# a_18248_44752# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1905 a_6671_43940# a_6109_44484# a_6453_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X1906 a_n1352_43396# a_n2433_43396# a_n1699_43638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1907 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1908 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1909 VDD a_n2302_37690# a_n4209_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1910 VDD a_n2946_37984# a_n3565_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1911 a_16131_47204# a_15507_47210# a_16023_47582# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1912 a_n23_44458# a_n356_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1913 VSS a_2779_44458# a_1307_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1914 a_11750_44172# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1915 a_7845_44172# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1916 VIN_N EN_VIN_BSTR_N C1_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1917 VSS a_6123_31319# a_7963_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1918 a_5907_46634# a_5732_46660# a_6086_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1919 a_8560_45348# a_8746_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X1920 a_19095_43396# a_13661_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X1921 a_21363_46634# a_21188_46660# a_21542_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1922 VSS a_n4315_30879# a_n4251_40480# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X1923 VSS a_n4064_39616# a_n2302_39866# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X1924 a_14180_46482# a_14035_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1925 a_n4064_37440# a_n4334_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X1926 a_18315_45260# a_18587_45118# a_18545_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1927 a_8349_46414# a_8016_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X1928 a_2537_44260# a_2479_44172# a_2127_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X1929 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1930 VSS a_3499_42826# a_3445_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1931 VDD a_3815_47204# a_4007_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1932 a_9306_43218# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1933 VDD a_6667_45809# a_6598_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1934 a_7230_45938# a_6511_45714# a_6667_45809# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1935 VDD a_2779_44458# a_1307_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X1936 a_8685_43396# a_8147_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X1937 VDD a_22400_42852# a_22589_40599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1938 VDD a_1273_38525# a_1666_39043# VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1939 VSS VSS a_3726_37500# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.589 pd=4.42 as=0.3135 ps=2.23 w=1.9 l=0.15
X1940 COMP_P a_1169_39587# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1941 a_8270_45546# a_n237_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1942 a_15765_45572# a_15599_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1943 a_3992_43940# a_768_44030# a_3737_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X1944 a_3815_47204# a_3785_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1945 a_2063_45854# a_9863_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1946 VSS a_11415_45002# a_22591_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1947 a_6755_46942# a_15015_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1948 VDD a_19431_45546# a_19418_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1949 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1950 VSS a_14021_43940# a_22959_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1951 a_19328_44172# a_19478_44306# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1386 ps=1.08 w=0.42 l=0.15
X1952 VSS a_10227_46804# a_14537_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1953 a_21073_44484# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1954 VDD a_768_44030# a_726_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X1955 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1956 VDD a_13059_46348# a_15297_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X1957 VSS a_12465_44636# a_22223_47212# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1958 VDD a_n1352_43396# a_n1177_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1959 VSS a_n863_45724# a_1067_42314# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1960 a_19164_43230# a_18083_42858# a_18817_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1961 a_383_46660# a_n133_46660# a_288_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1962 a_3524_46660# a_2443_46660# a_3177_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1963 a_13814_43218# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1964 VSS a_9127_43156# a_9061_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1965 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1966 VDD a_9482_43914# a_10157_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1967 VSS a_12607_44458# a_12553_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1968 a_n1057_35174# EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1969 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1970 VSS a_10903_43370# a_11963_45334# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1971 VSS a_17499_43370# a_17433_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1972 C1_P_btm a_1606_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1973 VDD a_12427_45724# a_10490_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X1974 a_13213_44734# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1975 VSS a_14815_43914# a_14761_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1976 a_12513_46660# a_12469_46902# a_12347_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1977 VDD a_n2302_39072# a_n4209_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1978 VSS a_11323_42473# a_10807_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1979 a_18989_43940# a_18451_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1980 VDD a_1209_43370# a_n1557_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1981 VSS a_8667_46634# a_8601_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1982 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1983 a_2889_44172# a_2998_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X1984 VSS a_7281_43914# a_7229_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1985 VSS a_21195_42852# a_21671_42860# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1986 a_n2956_38680# a_n2472_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1987 VSS a_n699_43396# a_4743_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X1988 VDD a_n443_46116# a_2437_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1989 a_n3565_39590# a_n2946_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X1990 a_10553_43218# a_10518_42984# a_10083_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1991 a_16789_44484# a_14537_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1992 VSS a_13635_43156# a_13569_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1993 a_18834_46812# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1994 a_10405_44172# a_7499_43078# a_10555_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X1995 a_n1151_42308# a_n1329_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X1996 VSS a_n2833_47464# CLK_DATA VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X1997 VSS a_18315_45260# a_18189_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X1998 a_n1917_43396# a_n2433_43396# a_n2012_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1999 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2000 a_n1441_43940# a_n2065_43946# a_n1549_44318# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2001 VDD a_17499_43370# a_17486_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2002 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2003 VDD a_22223_42860# a_22400_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2004 VDD a_3524_46660# a_3699_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2005 a_n1059_45260# a_17499_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2006 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2007 a_21753_35634# a_19998_35138# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2008 VSS a_12861_44030# a_17639_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2009 a_10765_43646# a_10695_43548# a_10057_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X2010 VDD a_12549_44172# a_20556_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2011 a_15890_42674# a_15803_42450# a_15486_42560# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X2012 VDD a_5815_47464# a_n1613_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2013 a_17433_43396# a_16243_43396# a_17324_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2014 VCM a_4958_30871# C9_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2015 a_11827_44484# a_3232_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2016 a_1847_42826# a_2351_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2017 VSS a_6151_47436# a_14955_47212# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2018 a_20205_31679# a_22223_46124# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2019 VSS a_15227_44166# a_15785_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2020 VDD a_1239_47204# a_1431_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2021 VDD a_8667_46634# a_8654_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2022 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2023 a_n452_45724# a_n443_46116# a_n310_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2024 a_700_44734# a_n746_45260# a_327_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X2025 a_19862_44208# a_13747_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2026 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2027 a_10775_45002# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X2028 a_3232_43370# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2029 VDD a_22959_44484# a_19237_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2030 a_1115_44172# a_453_43940# a_1443_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2031 a_484_44484# a_n863_45724# a_327_44734# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X2032 a_n3690_38528# a_n3674_38680# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2033 VDD a_14543_43071# a_13291_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2034 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2035 a_20512_43084# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2036 VSS a_12549_44172# a_21205_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2037 a_20256_43172# a_20202_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.203125 ps=1.275 w=0.65 l=0.15
X2038 a_6761_42308# a_n913_45002# a_6773_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2039 a_6298_44484# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2040 a_n2840_42282# a_n2661_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2041 a_n2661_46098# a_1983_46706# a_2162_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2042 a_5429_46660# a_5385_46902# a_5263_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2043 VSS a_15368_46634# a_15312_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2044 VDD a_8685_43396# a_14955_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X2045 VDD a_16855_45546# a_16842_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2046 VSS a_5815_47464# a_n1613_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2047 a_11315_46155# a_11133_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2048 a_16522_42674# a_15803_42450# a_15959_42545# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X2049 a_1221_42558# a_1184_42692# a_1149_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X2050 a_20885_46660# a_20841_46902# a_20719_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2051 a_20719_45572# a_20273_45572# a_20623_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2052 a_1756_43548# a_1307_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X2053 a_14456_42282# a_14635_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2054 a_n2472_42826# a_n2293_42834# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2055 a_7276_45260# a_6709_45028# a_7418_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2056 VDD a_1823_45246# a_3232_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2057 a_n4315_30879# a_n2302_40160# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2058 a_3260_45572# a_3218_45724# a_2957_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X2059 a_n2497_47436# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2060 VSS a_3422_30871# a_22315_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2061 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2062 VDD a_10341_42308# a_11554_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2063 a_11280_45822# a_2063_45854# a_10907_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X2064 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2065 a_603_45572# a_310_45028# a_509_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X2066 a_15002_46116# a_13925_46122# a_14840_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2067 a_8746_45002# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2068 a_n906_45572# a_n971_45724# a_n1013_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X2069 a_11064_45572# a_10903_43370# a_10907_45822# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X2070 a_21205_44306# a_20935_43940# a_21115_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X2071 a_2479_44172# a_2905_42968# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X2072 a_12861_44030# a_18143_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2073 DATA[3] a_7227_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X2074 VDD a_n2840_46090# a_n2956_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2075 VDD a_6945_45028# a_22223_46124# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2076 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2077 a_13556_45296# a_6755_46942# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2078 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2079 VCM a_7174_31319# C0_dummy_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2080 VDD a_8199_44636# a_9377_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X2081 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X2082 a_n4334_39392# a_n4318_39304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2083 a_12710_44260# a_10903_43370# a_12603_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X2084 a_13777_45326# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2085 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2086 a_16522_42674# a_15764_42576# a_15959_42545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X2087 a_14205_43396# a_13667_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X2088 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2089 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2090 VDD a_5732_46660# a_5907_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2091 a_6419_46155# a_5807_45002# a_6419_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2092 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X2093 a_n2860_39866# a_n2956_39768# a_n2946_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X2094 VDD a_13556_45296# a_13857_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2095 a_18533_44260# a_18326_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2096 a_n901_46420# a_n1076_46494# a_n722_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2097 a_5066_45546# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2098 w_1575_34946# a_n1057_35174# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=0 ps=0 w=3.75 l=15
X2099 a_18194_35068# a_n1794_35242# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2100 a_12861_44030# a_18143_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2101 VSS a_11599_46634# a_18175_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2102 VSS a_13635_43156# a_9290_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2103 VSS a_11599_46634# a_18819_46122# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2104 a_n3690_37440# a_n3674_37592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2105 VSS a_n3690_39616# a_n3420_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2106 a_n2442_46660# a_n2472_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2107 VSS a_n1435_47204# a_13487_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X2108 VDD a_3147_46376# a_526_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X2109 a_8317_43396# a_n755_45592# a_8229_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2110 a_n3674_38216# a_n2104_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2111 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2112 VDD a_n1794_35242# a_18194_35068# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2113 a_n2312_40392# a_n2288_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2114 VDD a_n1079_45724# a_n1099_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.28 ps=2.56 w=1 l=0.15
X2115 VSS a_22591_44484# a_17730_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2116 a_n914_42852# a_n1991_42858# a_n1076_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2117 a_n97_42460# a_19700_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2118 VDD a_n809_44244# a_n755_45592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2119 a_3877_44458# a_3699_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2120 VDD a_22537_40625# a_22725_37990# VDD sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2121 a_n913_45002# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2122 a_15368_46634# a_15143_45578# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X2123 a_11206_38545# CAL_N a_4338_37500# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2124 a_4905_42826# a_5379_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2125 VSS a_10467_46802# a_10428_46928# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2126 VSS a_3147_46376# a_526_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X2127 a_9313_45822# a_9049_44484# a_9159_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2128 a_21145_44484# a_20766_44850# a_21073_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X2129 VDD a_n4334_40480# a_n4064_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2130 VSS a_2680_45002# a_2274_45254# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X2131 VDD a_2324_44458# a_15682_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2132 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2133 a_22613_38993# a_22527_39145# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2134 a_10768_47026# a_10554_47026# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X2135 VSS a_21671_42860# a_3422_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2136 a_n785_47204# a_n815_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2137 a_5837_45028# a_5807_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X2138 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2139 C0_dummy_P_btm a_7174_31319# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2140 a_14537_43396# a_14358_43442# a_14621_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X2141 a_n3565_38216# a_n2946_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2142 a_n1736_43218# a_n1853_43023# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2143 a_6640_46482# a_5257_43370# a_6419_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X2144 VDD a_3090_45724# a_17786_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X2145 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2146 a_15493_43396# a_14955_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X2147 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2148 a_16877_42852# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X2149 a_9823_46482# a_9569_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X2150 VDD a_14021_43940# a_22959_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2151 VDD a_n3420_38528# a_n2860_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X2152 VSS a_10227_46804# a_12513_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2153 VDD a_3483_46348# a_17061_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2154 VSS a_17339_46660# a_19095_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2155 a_3699_46348# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X2156 VSS a_10533_42308# a_10723_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2157 VSS a_3537_45260# a_4223_44672# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2158 a_18214_42558# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X2159 VSS a_14537_43396# a_14180_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X2160 a_16501_45348# a_10193_42453# a_16405_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2161 VSS a_15743_43084# a_15567_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2162 VSS a_21259_43561# a_16922_45042# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2163 VSS a_n2840_46634# a_n2956_39768# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2164 a_9049_44484# a_8701_44490# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X2165 VDD a_2382_45260# a_3737_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2166 VDD a_n967_45348# a_n961_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2167 a_19615_44636# a_12861_44030# a_19789_44512# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2168 a_22589_40599# COMP_P VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2169 a_1273_38525# a_1107_38525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2170 VSS a_1169_39043# comp_n VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2171 a_9863_46634# a_10150_46912# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X2172 VDD a_n881_46662# a_n745_45366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2173 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2174 VDD a_21496_47436# a_13507_46334# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X2175 a_n2109_45247# a_n2017_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2176 VSS a_n143_45144# a_n37_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2177 a_19418_45938# a_18341_45572# a_19256_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2178 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2179 VDD a_n2438_43548# a_n2433_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2180 VDD a_5907_45546# a_5937_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X2181 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2182 C5_P_btm a_n4209_38502# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2183 VSS a_n452_44636# a_n2129_44697# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X2184 a_n2472_42282# a_n2293_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2185 a_n4318_38680# a_n2472_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2186 a_5608_44484# a_5111_44636# a_5518_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X2187 VDD a_742_44458# a_700_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X2188 VDD a_n901_43156# a_n443_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2189 VSS a_768_44030# a_13720_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X2190 VSS a_7287_43370# a_7221_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2191 VDD a_327_47204# DATA[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2192 a_2609_46660# a_2443_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2193 a_n89_44484# a_n467_45028# a_n452_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X2194 VDD a_9290_44172# a_9801_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X2195 VSS a_n1613_43370# a_6809_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2196 a_n4064_39616# a_n4334_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2197 a_556_44484# a_526_44458# a_484_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X2198 VDD a_n4334_39392# a_n4064_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2199 VSS a_4007_47204# DATA[2] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2200 VDD a_2324_44458# a_15682_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2201 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2202 a_2112_39137# a_1273_38525# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2203 VSS a_19328_44172# a_19279_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.169 ps=1.82 w=0.65 l=0.15
X2204 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X2205 a_n1696_35090# a_n1794_35242# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2206 VDD a_n3420_37440# a_n2860_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X2207 a_n3420_38528# a_n3690_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X2208 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2209 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2210 a_10554_47026# a_10467_46802# a_10150_46912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X2211 a_11387_46155# a_n1151_42308# a_11315_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2212 a_10341_43396# a_9803_43646# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2213 a_13887_32519# a_22223_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2214 VSS a_10227_46804# a_20885_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2215 C0_P_btm a_n3420_37440# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2216 VIN_P EN_VIN_BSTR_P C2_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2217 VSS a_16137_43396# a_18548_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X2218 a_n452_45724# a_n743_46660# a_n310_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2219 a_11682_45822# a_11652_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X2220 a_n443_42852# a_n901_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2221 VDD a_n2472_46090# a_n2956_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2222 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X2223 VDD a_11322_45546# a_11280_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X2224 VSS a_13747_46662# a_14495_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X2225 VDD a_10809_44734# a_n2661_42834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2226 SMPL_ON_P a_n2002_35608# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2227 C0_dummy_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2228 VSS a_n4209_39590# a_n4251_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X2229 VSS a_n1329_42308# a_n1151_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2230 a_3381_47502# a_2905_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2231 VDD a_18479_47436# a_13747_46662# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X2232 VSS a_n746_45260# a_261_44278# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2233 VDD a_n2302_39072# a_n4209_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2234 a_5649_42852# a_5111_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2235 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2236 a_11136_45572# a_3483_46348# a_11064_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X2237 VSS a_13249_42308# a_13904_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X2238 a_17486_43762# a_16409_43396# a_17324_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2239 VSS a_n913_45002# a_8325_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2240 VSS a_1307_43914# a_2675_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2241 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2242 a_3699_46634# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2243 VSS a_13259_45724# a_14797_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X2244 VSS a_2324_44458# a_949_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2245 a_20841_45814# a_20623_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2246 VIN_N EN_VIN_BSTR_N C9_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X2247 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2248 a_17639_46660# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2249 a_10341_42308# a_9803_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X2250 a_16327_47482# a_17591_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2251 VSS a_2324_44458# a_15682_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2252 a_1260_45572# a_n755_45592# a_1176_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X2253 a_20397_44484# a_20362_44736# a_20159_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X2254 a_12991_46634# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2255 a_518_46155# a_472_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2256 a_n4064_39072# a_n4334_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X2257 VDD a_20841_45814# a_20731_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2258 a_9751_46155# a_9569_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2259 a_1443_43940# a_1414_42308# a_1241_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2260 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=0.35
X2261 DATA[1] a_1431_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2262 VDD a_11823_42460# a_14033_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X2263 VSS a_n2840_42826# a_n3674_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2264 VSS a_3537_45260# a_5365_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X2265 a_3065_45002# a_3318_42354# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X2266 a_n310_45899# a_n356_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2267 C8_P_btm a_n3420_39616# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2268 a_16327_47482# a_17591_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2269 VDD a_22591_46660# a_20820_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2270 a_n3420_37440# a_n3690_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X2271 a_8337_42558# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2272 VDD a_4646_46812# a_7411_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2273 a_11186_47026# a_10428_46928# a_10623_46897# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X2274 a_20273_46660# a_20107_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2275 VSS a_3877_44458# a_2382_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2276 VDD a_n1331_43914# a_n1441_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2277 w_11334_34010# a_18194_35068# EN_VIN_BSTR_N w_11334_34010# sky130_fd_pr__pfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2278 VDD a_10835_43094# a_10796_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2279 VSS a_5066_45546# a_9159_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2280 VSS a_12883_44458# a_12829_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2281 a_11341_43940# a_10729_43914# a_11257_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3925 pd=1.785 as=0.135 ps=1.27 w=1 l=0.15
X2282 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2283 VSS a_564_42282# a_n1794_35242# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2284 a_12549_44172# a_20567_45036# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2285 VDD a_14456_42282# a_5342_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2286 a_645_46660# a_601_46902# a_479_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2287 VDD a_2063_45854# a_10809_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2288 VDD a_2127_44172# a_n2661_45010# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.26 ps=2.52 w=1 l=0.15
X2289 VDD a_10227_46804# a_16104_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X2290 a_12861_44030# a_18143_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2291 a_14513_46634# a_14180_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2292 a_n2840_46090# a_n2661_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2293 a_5088_37509# VSS VDAC_Ni VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2294 a_21137_46414# a_19692_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2295 a_1609_45822# a_167_45260# a_1609_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2296 VREF_GND a_17730_32519# C9_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2297 a_14635_42282# a_n913_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2298 a_10544_45572# a_10490_45724# a_10053_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X2299 a_10555_44260# a_10949_43914# a_10405_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.13325 ps=1.06 w=0.65 l=0.15
X2300 C2_P_btm a_n3565_38216# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2301 VSS a_1431_47204# DATA[1] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2302 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2303 a_8952_43230# a_7871_42858# a_8605_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2304 a_3067_47026# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2305 a_9377_42558# a_8685_42308# a_9293_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2306 a_4190_30871# a_19332_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2307 VDD a_9067_47204# DATA[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2308 a_15861_45028# a_15595_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2309 a_15194_46482# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2310 a_6469_45572# a_5907_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X2311 a_13720_44458# a_9482_43914# a_14112_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2312 a_15493_43940# a_14955_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2313 a_n1352_43396# a_n2267_43396# a_n1699_43638# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2314 a_16245_42852# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X2315 VSS a_n357_42282# a_6101_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2316 a_20692_30879# a_22959_46124# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2317 VSS a_n2302_37984# a_n4209_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2318 a_3177_46902# a_2959_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2319 a_5907_46634# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2320 a_5497_46414# a_5164_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2321 VSS a_104_43370# a_n971_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2322 VREF_GND a_13258_32519# C0_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2323 VDD a_4743_44484# a_4791_45118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2324 a_19700_43370# a_18579_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2325 a_12861_44030# a_18143_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X2326 a_21363_46634# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2327 VSS a_n443_42852# a_15940_43402# VSS sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X2328 a_12427_45724# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.14075 ps=1.325 w=0.42 l=0.15
X2329 VSS a_n3690_39616# a_n3420_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X2330 a_5891_43370# a_9127_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2331 a_n1920_47178# a_n1741_47186# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2332 a_10903_43370# a_13351_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2333 a_n955_45028# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2334 VDD a_n357_42282# a_7309_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2335 VDD a_3147_46376# a_526_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2336 a_18596_45572# a_18479_45785# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2337 a_4185_45028# a_3065_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2338 a_6575_47204# a_6545_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2339 a_16137_43396# a_15781_43660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X2340 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2341 VSS a_22775_42308# a_22485_38105# VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2342 VSS a_n2472_46634# a_n2442_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2343 a_4649_42852# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2344 VSS a_2711_45572# a_20107_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2345 VSS a_n2104_42282# a_n3674_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2346 VSS a_15015_46420# a_14949_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2347 VSS a_5691_45260# a_n2109_47186# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2348 a_18194_35068# a_n1794_35242# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2349 a_17583_46090# a_17715_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X2350 a_17730_32519# a_22591_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2351 a_3600_43914# a_1307_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X2352 a_13925_46122# a_13759_46122# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2353 VDD a_n901_43156# a_n914_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2354 a_8191_45002# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X2355 VDD a_22959_46124# a_20692_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2356 a_n310_44484# a_n356_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X2357 a_21125_42558# a_18597_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2358 VDD a_1169_39587# COMP_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2359 a_5932_42308# a_5755_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2360 VSS a_14543_43071# a_13291_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2361 VDD a_1307_43914# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2362 VSS a_3147_46376# a_526_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2363 VDD a_n2946_38778# a_n3565_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2364 VDD a_16112_44458# a_14673_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X2365 a_n1641_46494# a_n1991_46122# a_n1736_46482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2366 a_3175_45822# a_3316_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2367 VSS a_16763_47508# a_5807_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2368 VREF a_20447_31679# C5_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2369 a_14226_46660# a_14180_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X2370 VDD a_13348_45260# a_13159_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X2371 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2372 VDD a_6491_46660# a_6851_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2373 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2374 a_n4209_39590# a_n2302_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X2375 a_6511_45714# a_4646_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2376 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2377 VDD a_22775_42308# a_22485_38105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2378 a_3422_30871# a_21671_42860# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2379 VSS a_16763_47508# a_16697_47582# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2380 VDD a_2889_44172# a_413_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.34 ps=2.68 w=1 l=0.15
X2381 SMPL_ON_P a_n2002_35608# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2382 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2383 VSS a_n443_42852# a_1755_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2384 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2385 a_10405_44172# a_10729_43914# a_10651_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X2386 a_n2840_45546# a_n2661_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2387 a_14401_32519# a_22223_43948# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2388 VREF a_21076_30879# C8_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2389 a_4558_45348# a_4574_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2390 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2391 a_5193_42852# a_3905_42865# a_5111_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2392 a_18143_47464# a_18479_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X2393 a_10533_42308# a_n913_45002# a_10545_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2394 VDD a_16721_46634# a_16751_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2395 a_18909_45814# a_18691_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2396 VDD a_n1550_35608# a_n2002_35608# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2397 a_n2840_45002# a_n2661_45010# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2398 a_948_46660# a_n133_46660# a_601_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2399 a_3699_46348# a_3877_44458# a_3873_46454# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2400 a_117_45144# a_n443_42852# a_45_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X2401 a_11415_45002# a_13249_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2402 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2403 a_15681_43442# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2404 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2405 a_n4209_38502# a_n2302_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X2406 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2407 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=10
X2408 VDD a_n1059_45260# a_18727_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X2409 VSS a_5013_44260# a_5663_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2410 a_9801_43940# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2411 VSS a_10193_42453# a_18797_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2412 a_n4251_38304# a_n4318_38216# a_n4334_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X2413 a_2779_44458# a_1423_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2414 a_19789_44512# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X2415 VDD a_1107_38525# a_1273_38525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2416 comp_n a_1169_39043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2417 VDD a_18057_42282# a_n356_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X2418 a_13113_42826# a_12895_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2419 a_16197_42308# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X2420 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2421 VDD a_8034_45724# a_n1925_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X2422 VDD a_11691_44458# a_11649_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2423 VSS a_22581_37893# a_22537_39537# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2424 a_n3690_39392# a_n3674_39304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2425 a_15761_42308# a_15051_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X2426 a_16680_45572# a_15765_45572# a_16333_45814# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2427 VSS a_1568_43370# a_1512_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2428 VDD a_5066_45546# a_5024_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X2429 VSS a_n809_44244# a_n875_44318# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2430 VDD a_n2946_37690# a_n3565_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2431 a_n2267_43396# a_n2433_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2432 a_10518_42984# a_10796_42968# a_10752_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X2433 VDD a_1123_46634# a_584_46384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2434 a_8189_46660# a_8145_46902# a_8023_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2435 VDD a_13661_43548# a_14976_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X2436 a_11691_44458# a_5807_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2437 VSS a_n4064_39072# a_n2302_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X2438 a_20062_46116# a_18985_46122# a_19900_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2439 a_20269_44172# a_20365_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X2440 VSS a_5891_43370# a_5837_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2441 VSS a_n2472_42826# a_n4318_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2442 VSS a_7754_38470# a_7754_38470# VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2443 a_18707_42852# a_18083_42858# a_18599_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2444 VDD a_327_47204# DATA[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2445 a_12638_46436# a_13059_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2446 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2447 a_n784_42308# a_n961_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2448 a_13157_43218# a_13113_42826# a_12991_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2449 VSS a_4007_47204# DATA[2] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2450 VDD a_15015_46420# a_15002_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2451 VDD a_16327_47482# a_20159_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2452 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2453 VSS a_n785_47204# a_327_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X2454 a_18834_46812# a_13661_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X2455 a_n2840_45546# a_n2661_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2456 VSS a_21177_47436# a_20990_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2457 VSS a_7499_43078# a_11816_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X2458 a_n3420_38528# a_n3690_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2459 a_6761_42308# a_3537_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2460 a_10623_46897# a_10428_46928# a_10933_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X2461 a_5263_45724# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X2462 VDD a_11823_42460# a_11322_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2463 VSS a_5111_44636# a_8018_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X2464 a_7903_47542# a_n237_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2465 VSS a_8667_46634# a_n237_47217# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2466 a_3357_43084# a_4905_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2467 a_n2472_46090# a_n2293_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2468 VREF a_19237_31679# C0_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2469 VCM a_5742_30871# C6_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2470 VSS a_22589_40055# a_22527_39145# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2471 VDD a_n901_43156# a_n443_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2472 VSS a_22959_46660# a_21076_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2473 a_10249_46116# a_9823_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X2474 VDD a_10775_45002# a_10180_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X2475 CAL_N a_22485_38105# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2476 a_2684_37794# VDAC_Pi a_2113_38308# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2477 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2478 a_8696_44636# a_16855_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X2479 a_n4209_37414# a_n2302_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X2480 a_13467_32519# a_21487_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2481 a_6633_46155# a_5807_45002# a_6419_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X2482 a_n2661_42834# a_8975_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2483 a_n1243_43396# a_n2433_43396# a_n1352_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2484 VDD a_n2002_35608# SMPL_ON_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2485 a_7274_43762# a_6197_43396# a_7112_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2486 a_10922_42852# a_10835_43094# a_10518_42984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X2487 DATA[0] a_327_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2488 VDD a_5807_45002# a_11691_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2489 a_n1917_43396# a_n2267_43396# a_n2012_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2490 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2491 a_n4209_38502# a_n2302_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2492 VSS RST_Z a_14311_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2493 a_16327_47482# a_17591_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2494 a_18285_46348# a_18834_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2495 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2496 a_18597_46090# a_19431_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X2497 VSS a_18443_44721# a_18374_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X2498 VSS a_8199_44636# a_10951_45334# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2499 a_1176_45572# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X2500 a_7735_45067# a_6709_45028# a_7276_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X2501 C8_P_btm a_5342_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2502 DATA[4] a_9067_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2503 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=0.35
X2504 a_n3565_39304# a_n2946_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X2505 VSS a_n2109_45247# en_comp VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2506 a_n1076_43230# a_n1991_42858# a_n1423_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2507 DATA[1] a_1431_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2508 a_13348_45260# a_13556_45296# a_13490_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2509 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2510 a_n2302_40160# a_n2312_40392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2511 VSS a_21356_42826# a_n357_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2512 VDD a_11453_44696# a_22959_47212# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2513 VSS a_15037_45618# a_15143_45578# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2514 VSS a_8696_44636# a_8701_44490# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2515 a_3878_46660# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2516 a_2277_45546# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2517 a_626_44172# a_n863_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2518 a_18479_45785# a_19268_43646# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.3275 ps=1.655 w=1 l=0.15
X2519 SMPL_ON_N a_21753_35634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2520 a_16327_47482# a_17591_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X2521 a_20273_45572# a_20107_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2522 a_10555_44260# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X2523 a_n3420_37440# a_n3690_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2524 VSS a_n443_42852# a_742_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2525 VSS a_n901_43156# a_n967_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2526 a_20820_30879# a_22591_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2527 VSS a_13076_44458# a_12883_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X2528 a_685_42968# a_n443_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2529 a_17364_32525# a_22959_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2530 a_13170_46660# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2531 a_11633_42558# a_9290_44172# a_11551_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2532 VDD a_4791_45118# a_6633_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X2533 a_20731_45938# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2534 a_19700_43370# a_18579_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2535 VDD a_11599_46634# a_20107_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2536 a_16751_45260# a_17023_45118# a_16981_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2537 a_2382_45260# a_3877_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2538 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2539 VSS a_13487_47204# a_768_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2540 a_12829_44484# a_12741_44636# a_n2293_43922# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2541 a_11257_43940# a_10807_43548# a_11173_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2542 VCM a_6123_31319# C4_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2543 VSS a_14084_46812# a_14035_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X2544 VDD a_5937_45572# a_8034_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2545 a_5342_30871# a_14456_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2546 a_17639_46660# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
X2547 a_10809_44734# a_10057_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2548 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2549 VDD a_11823_42460# a_14853_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2550 a_20749_43396# a_20974_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2551 VDD a_11967_42832# a_16243_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2552 a_19511_42282# a_n913_45002# a_21125_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2553 VSS a_1431_47204# DATA[1] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2554 a_1609_45572# a_n443_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2555 a_17517_44484# a_16979_44734# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X2556 a_20075_46420# a_19900_46494# a_20254_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2557 a_n4209_37414# a_n2302_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2558 VDD a_10083_42826# a_7499_43078# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2559 a_16020_45572# a_15903_45785# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2560 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2561 a_20731_45938# a_20107_45572# a_20623_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2562 a_22629_38406# a_22581_37893# CAL_N VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2563 a_n1057_35174# a_n1696_35090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2564 VDD a_n3420_39072# a_n2860_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X2565 VSS a_22731_47423# a_13717_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2566 a_16855_45546# a_16680_45572# a_17034_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2567 a_18114_32519# a_22223_45036# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2568 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2569 a_17339_46660# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2570 a_n2472_45546# a_n2293_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2571 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2572 VSS a_18429_43548# a_16823_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2573 VSS a_n4334_38304# a_n4064_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2574 VSS a_8325_42308# a_8791_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2575 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2576 VDD a_n4334_38528# a_n4064_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2577 VSS a_768_44030# a_13076_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X2578 VSS a_12861_44030# a_19692_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2579 VDD a_14495_45572# a_n881_46662# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2580 a_18596_45572# a_18479_45785# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2581 a_n2472_45002# a_n2293_45010# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2582 VDD a_n881_46662# a_6431_45366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2583 a_5326_44056# a_5147_45002# a_5244_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2584 VSS a_22959_42860# a_14097_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2585 a_3445_43172# a_3357_43084# a_n2293_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2586 a_13003_42852# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2587 VSS a_9127_43156# a_5891_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2588 a_3503_45724# a_3775_45552# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2589 C6_N_btm a_14401_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2590 a_19929_45028# a_19778_44110# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2591 a_3540_43646# a_584_46384# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2592 VSS a_n2302_37984# a_n4209_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2593 DATA[4] a_9067_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2594 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2595 VDD a_167_45260# a_117_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X2596 a_6086_46660# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2597 a_3147_46376# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2598 a_n1533_46116# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2599 VSS a_n3565_38216# a_n3607_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X2600 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2601 a_5337_42558# a_5267_42460# a_4905_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X2602 a_21542_46660# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2603 a_10216_45572# a_10180_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X2604 a_4699_43561# a_3080_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2605 a_3626_43646# a_3232_43370# a_3457_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2606 a_n4064_37984# a_n4334_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X2607 VDD a_21613_42308# a_22775_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2608 a_16269_42308# a_15890_42674# a_16197_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X2609 a_1067_42314# a_1184_42692# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2610 VDD a_5937_45572# a_6945_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2611 COMP_P a_1169_39587# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2612 a_21356_42826# a_21381_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2613 VDD CLK a_8953_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2614 VDD a_2324_44458# a_949_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2615 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2616 VDD a_1307_43914# a_16237_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2617 a_n1549_44318# a_n2065_43946# a_n1644_44306# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2618 VSS a_19862_44208# a_19808_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2619 VDD a_5891_43370# a_8791_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2620 VSS a_n3690_39392# a_n3420_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2621 a_20256_43172# a_18494_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X2622 a_7927_46660# a_7411_46660# a_7832_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2623 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2624 VREF_GND a_13887_32519# C3_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2625 a_n3420_39072# a_n3690_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X2626 a_n2472_45546# a_n2293_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2627 a_17668_45572# a_n881_46662# a_17568_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X2628 C9_P_btm a_n4064_39616# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2629 a_4649_42852# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2630 a_6540_46812# a_3877_44458# a_6682_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2631 VDD a_6511_45714# a_6472_45840# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2632 VSS a_15493_43396# a_19478_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2633 a_16664_43396# a_16547_43609# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2634 VDD a_5068_46348# a_4955_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X2635 a_9159_44484# a_5883_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X2636 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2637 VSS a_10341_43396# a_22591_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2638 VDD a_n4334_37440# a_n4064_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2639 VSS a_17124_42282# a_4958_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2640 a_n1545_46494# a_n1991_46122# a_n1641_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2641 C8_P_btm a_n3565_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2642 a_5267_42460# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X2643 a_1138_42852# a_791_42968# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X2644 a_n4318_40392# a_n2840_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2645 a_n1644_44306# a_n1761_44111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2646 VDD a_7754_40130# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.5
X2647 VDD a_1609_45822# a_n2293_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X2648 a_5267_42460# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X2649 VREF_GND a_17364_32525# C7_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X2650 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2651 a_2127_44172# a_2675_43914# a_2455_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2652 a_11787_45002# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X2653 a_19250_35138# a_18194_35068# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2654 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2655 VDD a_17499_43370# a_n1059_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2656 VSS a_19333_46634# a_19123_46287# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X2657 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2658 a_n2946_37984# a_n2956_38216# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2659 a_3316_45546# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X2660 VSS a_13777_45326# a_13711_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2661 a_20712_42282# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2662 a_19479_31679# a_22223_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2663 a_20573_43172# a_20512_43084# a_20256_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.118625 ps=1.015 w=0.65 l=0.15
X2664 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2665 a_n2293_46634# a_14673_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2666 a_n1177_43370# a_n1352_43396# a_n998_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2667 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2668 VSS a_526_44458# a_5457_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2669 a_33_46660# a_n133_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2670 a_584_46384# a_1123_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2671 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2672 VDD a_10903_43370# a_10849_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X2673 VDD a_7754_40130# a_7754_40130# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X2674 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2675 a_8495_42852# a_7871_42858# a_8387_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2676 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2677 a_5495_43940# a_5244_44056# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X2678 a_16842_45938# a_15765_45572# a_16680_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2679 VDD a_167_45260# a_2521_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X2680 VDD a_2779_44458# a_1307_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2681 VSS a_n961_42308# a_n784_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2682 VSS a_13259_45724# a_17303_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2683 VDD a_5937_45572# a_5829_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X2684 a_17538_32519# a_22959_43948# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2685 a_21496_47436# a_4883_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2686 a_11816_44260# a_11750_44172# a_10729_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2687 a_9801_43940# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2688 a_5742_30871# a_10723_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2689 VDD a_15051_42282# a_11823_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2690 a_2123_42473# a_n784_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2691 a_13565_43940# a_12891_46348# a_13483_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2692 a_7227_42852# a_n97_42460# a_7309_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2693 a_5257_43370# a_5907_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2694 VDD a_13747_46662# a_13607_46688# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2695 a_1667_45002# a_1823_45246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X2696 a_n1655_44484# a_n1699_44726# a_n1821_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2697 a_n2293_46098# a_5663_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X2698 a_13003_42852# a_12379_42858# a_12895_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2699 a_2711_45572# a_768_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2700 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2701 DATA[0] a_327_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X2702 a_16763_47508# a_16588_47582# a_16942_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2703 a_4883_46098# a_21363_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2704 VSS a_16751_45260# a_6171_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X2705 VDD a_20835_44721# a_20766_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X2706 a_11750_44172# a_10903_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X2707 VSS a_15861_45028# a_17668_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X2708 a_7845_44172# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X2709 a_15597_42852# a_15743_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2710 a_n4064_39072# a_n4334_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2711 VSS a_9223_42460# a_8953_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X2712 VDD a_11967_42832# a_18083_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2713 a_13487_47204# a_13381_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.16535 ps=1.82 w=0.65 l=0.15
X2714 a_13297_45572# a_13259_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1034 ps=1 w=0.42 l=0.15
X2715 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2716 C2_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2717 C10_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2718 VDD a_n3565_38216# a_n3690_38304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X2719 a_6101_43172# a_5891_43370# a_5755_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2720 a_11901_46660# a_11735_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2721 a_16979_44734# a_14539_43914# a_17061_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2722 VSS a_14955_47212# a_10227_46804# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2723 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2724 a_18443_44721# a_18248_44752# a_18753_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X2725 VDD a_18909_45814# a_18799_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2726 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2727 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2728 a_1431_46436# a_1138_42852# a_1337_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X2729 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2730 VDD a_n4064_37984# a_n2216_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X2731 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2732 a_18443_44721# a_18287_44626# a_18588_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X2733 VDD a_768_44030# a_5326_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X2734 VSS a_n4209_39304# a_n4251_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X2735 a_n357_42282# a_21356_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2736 VSS a_n2288_47178# a_n2312_40392# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2737 a_491_47026# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2738 a_n901_46420# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2739 VSS a_3483_46348# a_15301_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2740 VCM a_1606_42308# C1_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2741 VDD a_20712_42282# a_10193_42453# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2742 VSS a_13635_43156# a_9290_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2743 a_5068_46348# a_5204_45822# a_5210_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2744 a_14033_45822# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2745 VSS a_11599_46634# a_20107_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2746 a_3537_45260# a_7287_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2747 w_1575_34946# EN_VIN_BSTR_P VDD w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2748 VSS a_6761_42308# a_7227_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2749 VDD a_13661_43548# a_15595_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2750 a_9803_42558# a_n97_42460# a_9885_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2751 VDD a_10227_46804# a_11136_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X2752 a_n1177_43370# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2753 VREF_GND a_n3420_39616# C8_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2754 VDD a_n2946_39072# a_n3565_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2755 a_601_46902# a_383_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2756 a_5024_45822# a_n443_46116# a_4419_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X2757 VDAC_Ni a_3754_38470# a_3726_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2758 a_17701_42308# a_17531_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2759 VSS a_12861_44030# a_13487_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X2760 w_11334_34010# a_11530_34132# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=0 ps=0 w=3.75 l=15
X2761 a_4808_45572# a_1823_45246# a_4419_46090# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X2762 a_6598_45938# a_6472_45840# a_6194_45824# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X2763 a_n229_43646# a_n2497_47436# a_n447_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2764 a_n3607_38304# a_n3674_38216# a_n3690_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X2765 VSS a_6969_46634# a_6903_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2766 a_18214_42558# a_18184_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X2767 a_491_47026# a_n133_46660# a_383_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2768 VSS a_4883_46098# a_10355_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X2769 VDD a_16327_47482# a_18588_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X2770 VDD a_4646_46812# a_6031_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2771 VSS a_n1613_43370# a_n1655_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2772 a_6812_45938# a_6598_45938# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X2773 a_8147_43396# a_n443_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X2774 VDAC_Ni VSS a_5088_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2775 a_12427_45724# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.1281 ps=1.03 w=0.42 l=0.15
X2776 C9_N_btm a_17730_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2777 VDD a_19594_46812# a_19551_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2778 a_n4318_37592# a_n1736_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2779 a_9290_44172# a_13635_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2780 VSS a_2698_46116# a_2804_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2781 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2782 a_1414_42308# a_1067_42314# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X2783 VSS a_5649_42852# a_22223_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2784 VDD a_13259_45724# a_14797_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2785 a_n2288_47178# a_n2109_47186# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2786 a_4817_46660# a_4651_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2787 a_8062_46155# a_8016_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2788 a_949_44458# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2789 a_13296_44484# a_12891_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X2790 VDD a_20623_43914# a_20365_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X2791 a_11601_46155# a_11309_47204# a_11387_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X2792 a_10210_45822# a_8746_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X2793 a_18287_44626# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2794 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2795 VSS a_11189_46129# a_11133_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X2796 a_n3565_38216# a_n2946_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X2797 a_6431_45366# a_5937_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2798 a_6109_44484# a_5518_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2799 a_14021_43940# a_13483_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X2800 a_17499_43370# a_17324_43396# a_17678_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2801 a_3495_45348# a_3429_45260# a_3316_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.182 ps=1.86 w=0.65 l=0.15
X2802 VDD a_1115_44172# a_n2293_45010# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.26 ps=2.52 w=1 l=0.15
X2803 VDD a_19787_47423# a_19594_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2804 a_18707_42852# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2805 a_19787_47423# START VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2806 a_8667_46634# a_8492_46660# a_8846_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2807 a_1208_46090# a_n881_46662# a_1431_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2808 a_5431_46482# a_n1151_42308# a_5068_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X2809 a_n1809_44850# a_n2433_44484# a_n1917_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2810 a_n2302_39866# a_n2442_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2811 VSS a_n2438_43548# a_2443_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2812 a_18797_44260# a_13661_43548# a_18451_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2813 a_19551_46910# a_19692_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2814 VDD a_8953_45546# a_8049_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2815 a_8697_45822# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2816 VDD a_10341_43396# a_22591_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2817 a_12005_46116# a_2063_45854# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2818 VSS a_12861_44030# a_18911_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.194 pd=1.95 as=0.1092 ps=1.36 w=0.42 l=0.15
X2819 a_1241_43940# a_584_46384# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1575 ps=1.315 w=1 l=0.15
X2820 VSS a_2123_42473# a_1184_42692# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2821 a_1273_38525# a_1107_38525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2822 a_16285_47570# a_16241_47178# a_16119_47582# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2823 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2824 a_1423_45028# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2825 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2826 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X2827 a_10617_44484# a_10440_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2828 C7_P_btm a_n4064_39072# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X2829 VSS a_1169_39043# comp_n VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2830 VSS a_961_42354# a_1067_42314# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2831 VDD a_4704_46090# a_1823_45246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2832 a_18479_47436# a_20075_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2833 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2834 VDD a_9313_45822# a_11459_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2835 a_n1809_44850# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2836 VSS a_n3690_39392# a_n3420_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X2837 a_19987_42826# a_10193_42453# a_20573_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X2838 VSS a_3785_47178# a_3815_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2839 VDD a_5891_43370# a_8375_44464# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2840 a_n3420_39072# a_n3690_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2841 VSS a_9863_46634# a_2063_45854# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X2842 a_7920_46348# a_n1151_42308# a_8062_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2843 VDD a_22889_38993# a_22581_37893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2844 a_19721_31679# a_22959_45036# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2845 a_19808_44306# a_19778_44110# a_19328_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2846 VDD a_10193_42453# a_11633_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2847 VDD a_15559_46634# a_13059_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2848 VDD a_11189_46129# a_11601_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X2849 a_5263_45724# a_5257_43370# a_5437_45600# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2850 a_12495_44260# a_12429_44172# a_10949_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.2275 ps=2 w=0.65 l=0.15
X2851 VSS a_n2840_43370# a_n4318_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2852 a_15037_43396# a_14205_43396# a_14955_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X2853 VSS a_4915_47217# a_12891_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2854 a_14084_46812# a_13885_46660# a_14226_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2855 a_6452_43396# a_6293_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2856 VSS a_1107_38525# a_1273_38525# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2857 a_7705_45326# a_7229_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2858 a_8953_45002# CLK VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2859 a_16981_45144# a_16922_45042# a_16886_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X2860 a_1115_44172# a_1307_43914# a_1241_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2861 a_19478_44306# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X2862 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2863 a_4223_44672# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2864 a_7174_31319# a_20107_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2865 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2866 VDD a_n2302_39866# a_n4209_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2867 VDD a_10227_46804# a_15051_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2868 CLK_DATA a_n2833_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2869 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2870 a_n2833_47464# a_n2497_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X2871 VSS a_8103_44636# a_7640_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X2872 a_15146_44811# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2873 a_n4209_39304# a_n2302_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2874 a_2903_45348# a_n971_45724# a_2809_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X2875 VSS a_3537_45260# a_8103_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2876 VSS a_21137_46414# a_21071_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2877 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2878 VSS a_1414_42308# a_2889_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2879 VDD a_1848_45724# a_1799_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X2880 VSS a_19279_43940# a_21398_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X2881 a_1666_39587# a_1273_38525# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2882 VSS a_n13_43084# a_n1853_43023# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2883 a_18479_45785# a_19268_43646# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2884 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2885 VSS a_22485_44484# a_20974_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2886 VSS a_n3420_37984# a_n2946_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X2887 a_5275_47026# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2888 a_5841_44260# a_5495_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X2889 C5_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2890 a_n2661_45546# a_4093_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2891 VSS a_n2302_38778# a_n4209_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2892 VSS a_5497_46414# a_5431_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2893 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2894 VDD a_19339_43156# a_19326_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2895 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2896 a_8137_45348# a_8049_45260# a_n2293_42834# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2897 VDD a_17499_43370# a_n1059_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2898 VDD a_6123_31319# a_7963_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2899 VDD a_12861_44030# a_17339_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2900 VSS a_19998_35138# a_21753_35634# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2901 a_10849_43646# a_10807_43548# a_10765_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2902 VSS a_13507_46334# a_18997_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2903 a_8560_45348# a_3483_46348# a_8488_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X2904 VDD a_n3690_38304# a_n3420_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2905 a_13249_42308# a_13070_42354# a_13333_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X2906 a_6969_46634# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2907 a_n2216_37984# a_n2810_45572# a_n2302_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X2908 VSS a_22223_46124# a_20205_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2909 a_6194_45824# a_6511_45714# a_6469_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X2910 a_17613_45144# a_8696_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2911 a_n229_43646# a_n97_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2912 VSS a_n1613_43370# a_n1379_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2913 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2914 VSS a_13747_46662# a_19862_44208# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2915 a_17303_42282# a_n913_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2916 a_8649_43218# a_8605_42826# a_8483_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2917 VSS a_n901_46420# a_n967_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2918 a_15004_44636# a_13556_45296# a_15146_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2919 a_11186_47026# a_10467_46802# a_10623_46897# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X2920 a_n1076_46494# a_n2157_46122# a_n1423_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2921 VSS a_526_44458# a_4169_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2922 a_n23_45546# a_n356_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2923 a_3353_43940# a_2998_44172# a_2675_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2924 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2925 a_18326_43940# a_18079_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2926 a_20922_43172# a_19862_44208# a_20753_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X2927 a_10334_44484# a_10157_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2928 VSS a_742_44458# a_1756_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2929 C5_P_btm a_5934_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2930 a_n2017_45002# a_19987_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.208 ps=1.94 w=0.65 l=0.15
X2931 a_n2956_38216# a_n2472_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2932 VDD a_10193_42453# a_13657_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2933 a_13885_46660# a_13607_46688# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2934 VDD a_8191_45002# a_n2293_42834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2935 VSS RST_Z a_7754_39964# VSS sky130_fd_pr__nfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.15
X2936 VSS a_4223_44672# a_n2497_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2937 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2938 a_4699_43561# a_3080_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2939 a_19511_42282# a_18597_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2940 a_n1991_46122# a_n2157_46122# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2941 a_n3420_37984# a_n3690_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X2942 VSS a_19692_46634# a_743_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2943 VDD a_22591_43396# a_14209_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2944 VDD a_7499_43078# a_8746_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2945 a_n971_45724# a_104_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2946 a_22889_38993# a_22400_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2947 VDD a_n4334_39392# a_n4064_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2948 a_20447_31679# a_22959_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2949 VDD a_15493_43940# a_22959_43948# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2950 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2951 VSS a_n2302_37690# a_n4209_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2952 a_18147_46436# a_17339_46660# a_17957_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2953 a_8336_45822# a_8270_45546# a_n1925_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X2954 VDD a_13527_45546# a_13163_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X2955 a_n4334_39616# a_n4318_39768# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2956 a_n2956_39304# a_n2840_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2957 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2958 VDD a_584_46384# a_766_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X2959 a_11361_45348# a_10907_45822# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2960 VDD a_11599_46634# a_11735_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2961 a_19431_45546# a_19256_45572# a_19610_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2962 VSS a_9290_44172# a_12710_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.118125 pd=1.04 as=0.08775 ps=0.92 w=0.65 l=0.15
X2963 VDD a_11323_42473# a_10807_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2964 a_2266_47243# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2965 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2966 a_2982_43646# a_2479_44172# a_2896_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2967 a_18280_46660# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2968 VDD a_8492_46660# a_8667_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2969 C1_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2970 VDD a_n1794_35242# a_18194_35068# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2971 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2972 VDD a_n1076_46494# a_n901_46420# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2973 a_n4251_38528# a_n4318_38680# a_n4334_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X2974 a_4361_42308# a_3823_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2975 VDD a_11967_42832# a_12379_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2976 VDD a_21811_47423# a_20916_46384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2977 VDD a_11599_46634# a_13759_46122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2978 a_18985_46122# a_18819_46122# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2979 VDD a_n971_45724# a_3775_45552# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2980 VDD a_5649_42852# a_22223_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2981 VSS a_5343_44458# a_8333_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2982 VDD a_7287_43370# a_3537_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2983 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2984 VSS a_3090_45724# a_10555_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X2985 a_20528_45572# a_19466_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2986 a_13487_47204# a_13717_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2987 VREF_GND a_13678_32519# C2_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2988 VDD a_22485_38105# a_22581_37893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2989 VDD a_20269_44172# a_19319_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X2990 a_5807_45002# a_16763_47508# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X2991 VSS a_16327_47482# a_16285_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2992 a_n23_44458# a_n356_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2993 VDD a_n1059_45260# a_8791_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2994 a_1847_42826# a_2351_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2995 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2996 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2997 VSS a_1169_39587# COMP_P VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2998 a_19553_46090# a_19335_46494# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2999 VDD a_n2840_45546# a_n2810_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3000 VSS a_3503_45724# a_3218_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X3001 a_15037_45618# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3002 a_14537_43646# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X3003 VDD a_1307_43914# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3004 a_6671_43940# a_5205_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3005 a_n1699_43638# a_n1917_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3006 C6_P_btm a_n3420_39072# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3007 VDD a_n2946_38778# a_n3565_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3008 VSS a_5111_44636# a_4905_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X3009 VDD a_9313_44734# a_22959_42860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3010 a_2124_47436# a_2063_45854# a_2266_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3011 VSS a_9625_46129# a_9569_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X3012 a_n4064_37984# a_n4334_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3013 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3014 VDD a_19279_43940# a_21398_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X3015 VDD a_3483_46348# a_13565_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3016 a_22725_38406# a_22589_40055# a_22629_38406# VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3017 a_6171_42473# a_5932_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3018 a_17568_45572# a_8696_44636# a_17478_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X3019 a_18588_44850# a_18374_44850# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X3020 a_18451_43940# a_18579_44172# a_18533_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3021 a_22485_38105# a_22775_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X3022 VSS a_5755_42308# a_5932_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3023 a_2959_46660# a_2609_46660# a_2864_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3024 a_21359_45002# a_21513_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3025 a_7_47243# a_n746_45260# a_n452_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3026 a_15227_46910# a_3090_45724# a_15009_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3027 a_14493_46090# a_14275_46494# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3028 a_19478_44306# a_15493_43396# a_19478_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X3029 a_7287_43370# a_7112_43396# a_7466_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3030 a_12251_46660# a_11901_46660# a_12156_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3031 a_8495_42852# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3032 a_n4251_37440# a_n4318_37592# a_n4334_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X3033 a_11633_42558# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X3034 VDD a_7276_45260# a_7227_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3035 VSS a_2479_44172# a_2813_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X3036 a_15279_43071# a_5342_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3037 VREF_GND a_14401_32519# C6_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3038 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3039 VDD a_n815_47178# a_n785_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3040 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3041 VSS a_n1794_35242# a_n1696_35090# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3042 a_1239_47204# a_1209_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3043 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3044 VDD a_3877_44458# a_3699_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3045 a_9313_45822# a_5937_45572# a_9241_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X3046 a_20841_45814# a_20623_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3047 VDD a_805_46414# a_835_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3048 a_12379_46436# a_12005_46116# a_n1741_47186# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3049 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3050 a_6298_44484# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3051 a_4338_37500# a_3754_38470# VDAC_Pi VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3052 a_961_42354# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3053 a_n2956_39768# a_n2840_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3054 a_n1741_47186# a_12594_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3055 VDD a_5257_43370# a_3905_42865# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3056 VSS en_comp a_1107_38525# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3057 VSS a_n473_42460# a_n1761_44111# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3058 a_13163_45724# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.1281 ps=1.03 w=0.42 l=0.15
X3059 VDD a_10227_46804# a_9863_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3060 a_10210_45822# a_10586_45546# a_10053_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3061 comp_n a_1169_39043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3062 VSS a_4185_45028# a_22959_45036# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3063 a_22485_38105# a_22775_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X3064 VDD a_n2438_43548# a_n2065_43946# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3065 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X3066 a_5457_43172# a_5111_44636# a_5111_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3067 VDD a_11787_45002# a_11652_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X3068 a_10695_43548# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X3069 VDD a_n2946_37690# a_n3565_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3070 a_13059_46348# a_15559_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3071 VDD a_n23_44458# a_7_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3072 a_12891_46348# a_4915_47217# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3073 a_8023_46660# a_7577_46660# a_7927_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3074 VSS a_10057_43914# a_9672_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X3075 a_n237_47217# a_8667_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X3076 a_n143_45144# a_n755_45592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3077 a_20637_44484# a_20159_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X3078 a_4520_42826# a_4905_42826# a_4649_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3079 VSS a_n971_45724# a_8423_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X3080 VSS RST_Z a_8530_39574# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3081 VSS a_n2946_37984# a_n3565_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3082 a_n1379_43218# a_n1423_42826# a_n1545_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3083 a_8697_45822# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3084 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3085 VDD a_n4334_39616# a_n4064_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3086 VSS a_3626_43646# a_19647_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3087 a_n443_42852# a_n901_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3088 VDD a_1209_47178# a_1239_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3089 a_3094_47243# a_2905_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3090 a_15051_42282# a_15486_42560# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X3091 a_n1641_46494# a_n2157_46122# a_n1736_46482# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3092 VDD a_13661_43548# a_16241_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X3093 a_11823_42460# a_15051_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3094 a_5167_46660# a_4817_46660# a_5072_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3095 VSS a_10835_43094# a_10796_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3096 VDD a_20708_46348# a_20411_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3097 VSS a_16327_47482# a_18005_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X3098 VSS a_16292_46812# a_15811_47375# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X3099 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3100 a_9482_43914# a_9838_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3101 a_20623_46660# a_20273_46660# a_20528_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3102 VDD a_12594_46348# a_n1741_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3103 a_18374_44850# a_18287_44626# a_17970_44736# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X3104 a_16750_47204# a_15673_47210# a_16588_47582# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3105 a_6545_47178# a_6419_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X3106 a_8783_44734# a_8696_44636# a_8701_44490# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3107 a_175_44278# a_n863_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3108 VDD a_22400_42852# a_22589_40055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3109 VDD a_22223_43396# a_13887_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3110 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3111 VSS a_n901_46420# a_n443_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3112 VDD a_18479_47436# a_20935_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X3113 VSS a_7754_38470# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0 ps=0 w=2 l=0.15
X3114 VSS a_5907_46634# a_5841_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3115 a_5745_43940# a_5883_43914# a_5829_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3116 VSS a_18194_35068# a_19250_35138# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3117 a_3754_38470# a_7754_38470# VSS sky130_fd_pr__res_high_po_0p35 l=18
X3118 a_1110_47026# a_33_46660# a_948_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3119 a_16434_46987# a_16388_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3120 VSS a_2324_44458# a_15682_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3121 VDD a_n2302_39866# a_n4209_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3122 a_13381_47204# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3123 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3124 a_2998_44172# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3125 a_20974_43370# a_22485_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3126 VDD a_4921_42308# a_5755_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3127 a_10991_42826# a_10835_43094# a_11136_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X3128 VDD a_6851_47204# a_7227_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3129 a_3052_44056# a_2998_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14575 ps=1.335 w=0.42 l=0.15
X3130 VDD a_n2002_35608# SMPL_ON_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3131 VSS a_n4334_38528# a_n4064_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3132 a_3177_46902# a_2959_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3133 VSS a_1208_46090# a_472_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X3134 a_9241_44734# a_5937_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3135 a_n1699_43638# a_n1917_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3136 a_22365_46825# EN_OFFSET_CAL VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3137 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3138 VSS a_13163_45724# a_11962_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3139 a_3055_46660# a_2609_46660# a_2959_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3140 a_19326_42852# a_18249_42858# a_19164_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3141 a_n443_46116# a_n901_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3142 a_9885_43646# a_8270_45546# a_9803_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3143 VDD a_18597_46090# a_16375_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3144 a_19431_45546# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3145 VSS a_22959_43396# a_17364_32525# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3146 VDD a_n3690_38304# a_n3420_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X3147 a_n4064_39616# a_n4334_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X3148 VSS a_n1177_44458# a_n1243_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3149 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3150 VSS a_n23_45546# a_n89_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X3151 a_n452_47436# a_n746_45260# a_n310_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3152 a_2952_47436# a_n1151_42308# a_3094_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3153 VDD a_12816_46660# a_12991_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3154 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3155 a_7499_43940# a_7640_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3156 w_11334_34010# a_11530_34132# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=1.0875 pd=8.08 as=0 ps=0 w=3.75 l=15
X3157 VSS a_n2302_38778# a_n4209_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3158 a_4235_43370# a_3935_42891# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X3159 a_5105_45348# a_4558_45348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X3160 a_18051_46116# a_765_45546# a_17957_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X3161 a_n1441_43940# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3162 a_15301_44260# a_15227_44166# a_14955_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3163 a_n746_45260# a_n1177_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X3164 VSS a_n3565_38502# a_n3607_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X3165 a_n2840_43914# a_n2661_43922# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3166 a_6809_43396# a_6765_43638# a_6643_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3167 VSS a_376_46348# a_171_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X3168 a_19443_46116# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3169 VSS a_13059_46348# a_15143_45578# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3170 VSS a_8199_44636# a_8701_44490# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3171 a_7499_43940# a_3090_45724# a_7281_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3172 a_9165_43940# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3173 a_453_43940# a_175_44278# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X3174 a_9885_42308# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3175 a_n3674_39304# a_n2840_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3176 a_2959_46660# a_2443_46660# a_2864_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3177 a_14543_46987# a_13885_46660# a_14084_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3178 VDD a_413_45260# a_22959_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3179 a_17969_45144# a_16375_45002# a_17896_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
X3180 a_n4064_38528# a_n4334_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X3181 a_16292_46812# a_n743_46660# a_16434_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3182 a_21188_46660# a_20107_46660# a_20841_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3183 a_12251_46660# a_11735_46660# a_12156_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3184 a_4365_46436# a_4185_45028# a_n1925_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3185 a_n998_44484# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3186 VDD a_3177_46902# a_3067_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3187 a_7577_46660# a_7411_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3188 VDD a_n2472_45546# a_n2956_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3189 a_14976_45028# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X3190 a_10835_43094# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3191 a_12638_46436# a_12891_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X3192 a_n1352_44484# a_n2433_44484# a_n1699_44726# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3193 a_n3420_37984# a_n3690_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3194 VSS a_13661_43548# a_743_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3195 a_12839_46116# a_12891_46348# a_n1741_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3196 VSS a_3090_45724# a_4927_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3197 VSS a_22000_46634# a_15227_44166# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3198 VSS a_n863_45724# a_791_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3199 a_14209_32519# a_22591_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3200 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3201 VSS a_n4334_37440# a_n4064_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3202 a_n1613_43370# a_5815_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3203 a_n2661_43922# a_12465_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3204 a_n2012_43396# a_n2129_43609# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3205 VSS a_11823_42460# a_14635_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3206 a_19692_46634# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3207 C8_P_btm a_n3565_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3208 VSS a_4520_42826# a_4093_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X3209 a_5013_44260# a_3905_42865# a_5025_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3210 a_8018_44260# a_7499_43078# a_7911_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X3211 VDD a_11823_42460# a_14358_43442# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X3212 a_167_45260# a_2202_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3213 a_20254_46482# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3214 VDD a_10405_44172# a_8016_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X3215 VIN_N EN_VIN_BSTR_N C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X3216 a_742_44458# a_n443_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3217 VSS a_19332_42282# a_4190_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3218 a_14840_46494# a_13925_46122# a_14493_46090# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3219 VSS a_1414_42308# a_3457_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X3220 a_20356_42852# a_18184_42460# a_20256_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.175 ps=1.35 w=1 l=0.15
X3221 a_19006_44850# a_18287_44626# a_18443_44721# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X3222 a_9420_43940# a_768_44030# a_9165_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X3223 VDD a_10903_43370# a_12005_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3224 a_n4209_38216# a_n2302_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3225 VSS a_12861_44030# a_18280_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3226 VSS a_13661_43548# a_15685_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X3227 C4_P_btm a_6123_31319# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X3228 a_13575_42558# a_n97_42460# a_13657_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3229 VSS a_n2302_37690# a_n4209_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3230 a_8667_46634# a_6151_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3231 a_n1613_43370# a_5815_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3232 VDD a_n971_45724# a_n229_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3233 a_n1533_42852# a_n2157_42858# a_n1641_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3234 a_21335_42336# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3235 VSS a_n3565_37414# a_n3607_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X3236 a_n2946_38778# a_n2956_38680# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3237 VSS a_9127_43156# a_5891_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3238 VSS a_13351_46090# a_10903_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X3239 a_14309_45028# a_2711_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X3240 VSS a_413_45260# a_22959_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3241 a_743_42282# a_12549_44172# a_20749_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3242 VDD a_3877_44458# a_4185_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3243 a_13105_45348# a_13017_45260# a_n2661_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3244 VSS a_6545_47178# a_6575_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3245 a_8229_43396# a_7499_43078# a_8147_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X3246 a_19551_46910# a_19466_46812# a_19333_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3247 a_18280_46660# a_12549_44172# a_17609_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X3248 VSS a_18285_46348# a_18243_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.104 ps=0.97 w=0.65 l=0.15
X3249 a_6945_45028# a_5205_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3250 a_3726_37500# a_3754_38470# VDAC_Ni VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3251 a_n4064_37440# a_n4334_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X3252 a_20708_46348# a_20916_46384# a_20850_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3253 a_5167_46660# a_4651_46660# a_5072_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3254 VDD a_n1352_44484# a_n1177_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3255 a_15685_45394# a_15415_45028# a_15595_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3256 VDD a_10193_42453# a_18214_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X3257 a_21350_45938# a_20273_45572# a_21188_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3258 a_7639_45394# a_n1151_42308# a_7276_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X3259 VSS a_526_44458# a_10149_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3260 a_7765_42852# a_7227_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X3261 a_501_45348# a_413_45260# a_375_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3262 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3263 COMP_P a_1169_39587# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3264 a_16547_43609# a_16414_43172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25675 ps=1.44 w=0.65 l=0.15
X3265 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3266 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3267 a_n3565_38502# a_n2946_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3268 a_5891_43370# a_9127_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3269 a_13857_44734# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3270 a_n2661_46098# a_2107_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X3271 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3272 VSS a_16327_47482# a_18953_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3273 VSS a_742_44458# a_1568_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3274 a_19273_43230# a_18083_42858# a_19164_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3275 a_6123_31319# a_7227_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3276 a_768_44030# a_13487_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X3277 a_584_46384# a_1123_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3278 VDD a_2711_45572# a_4099_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3279 a_12293_43646# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3280 C8_N_btm a_5342_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3281 a_8035_47026# a_6151_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3282 a_10306_45572# a_10193_42453# a_10216_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X3283 a_18545_45144# a_13259_45724# a_18450_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X3284 a_n1917_44484# a_n2433_44484# a_n2012_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3285 a_22629_37990# a_22537_39537# CAL_P VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3286 a_n1423_46090# a_n1641_46494# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3287 a_16977_43638# a_16759_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3288 VDD a_21855_43396# a_13678_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3289 VDD a_6540_46812# a_6491_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3290 VDD a_22223_43948# a_14401_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3291 VDD a_n863_45724# a_n1099_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3292 C10_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X3293 a_n2946_37690# a_n2956_37592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3294 a_5111_42852# a_4905_42826# a_5193_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3295 VDD a_5263_45724# a_5204_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X3296 a_n467_45028# a_n745_45366# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3297 VSS a_765_45546# a_1208_46090# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X3298 VDD a_15095_43370# a_14955_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X3299 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X3300 a_n2002_35608# a_n1550_35608# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3301 VSS a_n4334_38304# a_n4064_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X3302 VDD a_2957_45546# a_2905_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3303 a_8855_44734# a_4791_45118# a_8783_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3304 a_11963_45334# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X3305 a_n2661_44458# a_11453_44696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.182 ps=1.92 w=0.7 l=0.15
X3306 VDD a_4915_47217# a_11415_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3307 a_n1741_47186# a_12005_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3308 a_3600_43914# a_3537_45260# a_3820_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3309 a_21588_30879# a_22223_47212# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3310 a_1848_45724# a_2063_45854# a_1990_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3311 a_14537_46482# a_14493_46090# a_14371_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3312 a_10425_46660# a_9863_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X3313 a_16241_44734# a_2711_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X3314 a_3905_42865# a_5257_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3315 a_21811_47423# SINGLE_ENDED VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3316 a_19365_45572# a_18175_45572# a_19256_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3317 VDD a_22959_45572# a_20447_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3318 a_3090_45724# a_18911_45144# a_19113_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3319 DATA[2] a_4007_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3320 a_13777_45326# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X3321 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3322 VCM a_5934_30871# C5_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3323 a_n3690_39616# a_n3674_39768# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3324 a_17333_42852# a_16795_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3325 a_11525_45546# a_11962_45724# a_11682_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X3326 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3327 a_17595_43084# a_13259_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X3328 a_n13_43084# a_n755_45592# a_133_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X3329 a_11530_34132# EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3330 a_n3565_37414# a_n2946_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3331 a_n2840_42282# a_n2661_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3332 a_20193_45348# a_18184_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3333 a_20719_46660# a_20273_46660# a_20623_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3334 a_1756_43548# a_768_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3335 VSS a_n1613_43370# a_n1379_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3336 a_n2472_43914# a_n2293_43922# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3337 a_n2302_39072# a_n2312_39304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3338 a_14456_42282# a_14635_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3339 VDD a_20075_46420# a_20062_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3340 VSS a_2711_45572# a_4099_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3341 a_4927_45028# a_5147_45002# a_5105_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X3342 a_21381_43940# a_21115_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X3343 VSS a_10227_46804# a_10185_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X3344 a_n3607_38528# a_n3674_38680# a_n3690_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X3345 a_4169_42308# a_1823_45246# a_3823_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3346 CLK_DATA a_n2833_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X3347 VDD a_20894_47436# a_20843_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X3348 a_4704_46090# a_4883_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3349 VSS a_n913_45002# a_6761_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3350 VDD a_12465_44636# a_22223_47212# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3351 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3352 VDD a_15051_42282# a_11823_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3353 VDD a_20193_45348# a_20753_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3354 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3355 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X3356 VDD a_5257_43370# a_3357_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3357 VSS a_14113_42308# a_16522_42674# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X3358 a_22589_40055# en_comp VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3359 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3360 a_13460_43230# a_12379_42858# a_13113_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3361 a_19240_46482# a_19123_46287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3362 a_5829_43940# a_5495_43940# a_5745_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3363 a_10227_46804# a_14955_47212# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3364 VSS a_21487_43396# a_13467_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3365 VDD a_7287_43370# a_7274_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3366 VDD a_12861_44030# a_18911_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1468 pd=1.34 as=0.1092 ps=1.36 w=0.42 l=0.15
X3367 a_14955_43940# a_14537_43396# a_15037_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3368 a_15953_42852# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3369 a_9114_42852# a_8037_42858# a_8952_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3370 a_n4315_30879# a_n2302_40160# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X3371 VSS a_n901_46420# a_n443_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3372 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3373 VSS a_8199_44636# a_8953_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X3374 a_18780_47178# a_18597_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3375 VDD a_15227_44166# a_18285_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3376 a_16375_45002# a_18597_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3377 VDD a_2324_44458# a_6298_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3378 a_15279_43071# a_5342_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3379 a_10193_42453# a_20712_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3380 a_19335_46494# a_18985_46122# a_19240_46482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3381 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3382 a_5205_44484# a_5111_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3383 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3384 a_4842_47243# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3385 SMPL_ON_N a_21753_35634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3386 VSS a_685_42968# a_791_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3387 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3388 VSS a_22591_45572# a_19963_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3389 C8_N_btm a_21076_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3390 a_509_45572# a_n1099_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X3391 VSS a_11322_45546# a_12016_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X3392 a_n1059_45260# a_17499_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3393 a_20753_42852# a_10193_42453# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X3394 DATA[5] a_11459_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3395 a_16789_45572# a_15599_45572# a_16680_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3396 a_20362_44736# a_20640_44752# a_20596_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X3397 a_13622_42852# a_12545_42858# a_13460_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3398 a_n1991_42858# a_n2157_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3399 a_15143_45578# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3400 VSS a_n746_45260# a_556_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X3401 a_8701_44490# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3402 a_n3607_37440# a_n3674_37592# a_n3690_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X3403 a_10775_45002# a_10951_45334# a_10903_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X3404 VDD a_21753_35634# SMPL_ON_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3405 VSS a_7227_47204# DATA[3] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3406 VDD a_6151_47436# a_14955_47212# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3407 a_15673_47210# a_15507_47210# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3408 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3409 VDD a_22589_40599# a_22537_40625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3410 a_20679_44626# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3411 VDD a_n2946_39072# a_n3565_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3412 VDD a_10991_42826# a_10922_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X3413 a_5815_47464# a_6151_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X3414 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X3415 a_n2956_37592# a_n2472_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3416 a_13667_43396# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X3417 VSS a_n1920_47178# a_n2312_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3418 VDD a_n4064_40160# a_n2216_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X3419 a_5164_46348# a_4927_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X3420 a_949_44458# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3421 a_15940_43402# a_12549_44172# a_15868_43402# VSS sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X3422 VDD a_4646_46812# a_4651_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3423 a_1427_43646# a_1049_43396# a_1209_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3424 a_19164_43230# a_18249_42858# a_18817_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3425 VDD a_12861_44030# a_21845_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3426 a_2982_43646# a_3232_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X3427 VDD a_3600_43914# a_3499_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X3428 a_648_43396# a_526_44458# a_548_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X3429 a_16409_43396# a_16243_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3430 VSS a_2063_45854# a_11136_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X3431 VSS a_1823_45246# a_2202_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3432 a_10903_45394# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X3433 VDD a_n3420_39616# a_n2860_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X3434 a_18243_46436# a_18189_46348# a_18147_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.10725 ps=0.98 w=0.65 l=0.15
X3435 VSS a_n971_45724# a_3775_45552# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3436 a_9290_44172# a_13635_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3437 a_4700_47436# a_4915_47217# a_4842_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3438 VDD a_6453_43914# a_n2661_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3439 VSS a_n2438_43548# a_n2433_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3440 a_11813_46116# a_11387_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X3441 VDD a_380_45546# a_n356_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X3442 VDD a_10053_45546# a_9625_46129# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X3443 VDD a_12861_44030# a_19615_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3444 a_2253_43940# a_n443_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1575 ps=1.315 w=1 l=0.15
X3445 VDD a_13113_42826# a_13003_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3446 a_765_45546# a_17609_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X3447 a_3503_45724# a_1823_45246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X3448 VDD a_3699_46348# a_3160_47472# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X3449 VDD a_9625_46129# a_10037_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X3450 VDD a_22223_45036# a_18114_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3451 a_18997_42308# a_18727_42674# a_18907_42674# VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3452 a_5755_42852# a_n97_42460# a_5837_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3453 EN_VIN_BSTR_P a_n1696_35090# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3454 VDAC_Pi VSS a_5700_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3455 a_12281_43396# a_n913_45002# a_12293_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3456 VDD a_10533_42308# a_10723_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3457 VSS a_9863_47436# a_9804_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X3458 a_8049_45260# a_n237_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3459 a_11387_46482# a_11133_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X3460 VDD a_21005_45260# a_19778_44110# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X3461 VDD a_8791_42308# a_5934_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3462 VDD a_13487_47204# a_768_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3463 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X3464 a_895_43940# a_644_44056# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X3465 VSS a_n3420_38528# a_n2946_38778# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X3466 VDD a_4646_46812# a_7871_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3467 a_3067_47026# a_2443_46660# a_2959_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3468 a_19256_45572# a_18341_45572# a_18909_45814# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3469 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3470 C3_P_btm a_n4064_37984# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X3471 VSS a_2713_42308# a_2903_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3472 a_9863_47436# a_2063_45854# a_10037_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3473 a_15037_45618# a_13259_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3474 a_3726_37500# CAL_P a_11206_38545# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3475 a_10991_42826# a_10796_42968# a_11301_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X3476 a_2127_44172# a_1307_43914# a_2253_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X3477 a_1823_45246# a_4704_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3478 VDD a_n2438_43548# a_n2433_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3479 a_17678_43396# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3480 a_n452_47436# a_n237_47217# a_n310_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3481 VDD a_10903_43370# a_12427_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.06615 ps=0.735 w=0.42 l=0.15
X3482 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3483 a_3080_42308# a_2903_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3484 a_22581_37893# a_22613_38993# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X3485 a_18057_42282# a_n1059_45260# a_18310_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X3486 VSS a_n452_45724# a_n1853_46287# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X3487 a_n3674_39768# a_n2472_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3488 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3489 a_8846_46660# a_6151_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3490 a_1307_43914# a_2779_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3491 a_22365_46825# EN_OFFSET_CAL VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3492 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=10
X3493 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3494 a_1273_38525# a_1107_38525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3495 a_n89_45572# a_n743_46660# a_n452_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X3496 a_n2472_42282# a_n2293_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3497 VSS a_n2840_45002# a_n2810_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3498 a_11530_34132# a_18194_35068# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3499 a_15928_47570# a_15811_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3500 a_518_46482# a_472_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X3501 a_15463_44811# a_11691_44458# a_15004_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3502 VSS a_17767_44458# a_17715_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X3503 a_20556_43646# a_19692_46634# a_20301_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3504 a_n3420_39616# a_n3690_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X3505 a_14309_45028# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3506 a_16237_45028# a_16375_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3507 a_8791_43396# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3508 VDD a_22589_40599# a_22725_38406# VDD sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3509 VDD a_n4209_38216# a_n4334_38304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X3510 a_9061_43230# a_7871_42858# a_8952_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3511 a_1568_43370# a_n863_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3512 VDD a_n1423_42826# a_n1533_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3513 a_n1379_46482# a_n1423_46090# a_n1545_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3514 a_13575_42558# a_n97_42460# a_13657_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3515 a_6667_45809# a_6511_45714# a_6812_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X3516 a_3754_39964# a_7754_39964# VSS sky130_fd_pr__res_high_po_0p35 l=18
X3517 VSS a_9290_44172# a_10586_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3518 a_16115_45572# a_15765_45572# a_16020_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3519 VDD a_18911_45144# a_3090_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.165 ps=1.33 w=1 l=0.15
X3520 a_2725_42558# a_n755_45592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3521 a_18504_43218# a_17333_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3522 VDD a_3499_42826# a_n2293_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3523 a_16979_44734# a_14539_43914# a_17061_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3524 a_2253_43940# a_2479_44172# a_2455_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3525 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3526 VSS a_1307_43914# a_3681_42891# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X3527 a_n310_47243# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3528 a_5025_43940# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3529 VSS a_626_44172# a_648_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X3530 VSS a_n3420_37440# a_n2946_37690# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X3531 a_n3420_38528# a_n3690_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X3532 a_21356_42826# a_21381_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3533 a_16877_43172# a_16823_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3534 a_20841_46902# a_20623_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3535 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X3536 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3537 VSS a_6171_45002# a_6125_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3538 VSS a_17595_43084# a_14539_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X3539 a_21137_46414# a_19692_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X3540 a_5883_43914# a_8333_44056# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X3541 a_20766_44850# a_20640_44752# a_20362_44736# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X3542 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3543 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3544 a_805_46414# a_472_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3545 a_1176_45822# a_997_45618# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X3546 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3547 a_21887_42336# a_20202_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3548 VSS a_11967_42832# a_18083_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3549 DATA[2] a_4007_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X3550 VDD a_1823_45246# a_3316_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3551 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3552 a_21513_45002# a_21363_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X3553 a_8704_45028# a_5937_45572# a_8191_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X3554 a_3232_43370# a_1823_45246# a_3363_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3555 a_13333_42558# a_13291_42460# a_13249_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3556 a_13661_43548# a_18780_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3557 a_5497_46414# a_5164_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X3558 a_12749_45572# a_12549_44172# a_12649_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X3559 VSS a_n2840_43914# a_n4318_39768# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3560 a_15037_44260# a_13556_45296# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3561 VSS a_22223_45572# a_19479_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3562 w_1575_34946# a_n1057_35174# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=0 ps=0 w=3.75 l=15
X3563 VDD a_n2438_43548# a_n133_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3564 VDD a_n984_44318# a_n809_44244# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3565 VDD a_14815_43914# a_n2293_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3566 a_n1545_43230# a_n1991_42858# a_n1641_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3567 a_8128_46384# a_7903_47542# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3568 VDD a_7281_43914# a_7229_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3569 VDD a_13507_46334# a_18907_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3570 CLK_DATA a_n2833_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3571 a_479_46660# a_33_46660# a_383_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3572 VSS a_6667_45809# a_6598_45938# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X3573 VDD a_13904_45546# a_12594_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X3574 VDD a_n881_46662# a_n1021_46688# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3575 VDD a_2324_44458# a_15682_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3576 a_8568_45546# a_8953_45546# a_8697_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3577 a_17767_44458# a_17970_44736# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X3578 VREF a_19479_31679# C1_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X3579 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3580 VDD a_n755_45592# a_133_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X3581 a_16241_44734# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3582 a_10867_43940# a_7499_43078# a_10405_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
X3583 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3584 VDD a_10723_42308# a_5742_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3585 a_11823_42460# a_15051_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3586 a_20556_43646# a_20974_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3587 a_n3420_37440# a_n3690_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X3588 a_4574_45260# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X3589 a_13483_43940# a_13249_42308# a_13565_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3590 VDD a_20159_44458# a_19321_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X3591 a_n1352_44484# a_n2267_44484# a_n1699_44726# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3592 a_2583_47243# a_584_46384# a_2124_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3593 a_22612_30879# a_22959_47212# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3594 VDD a_8349_46414# a_8379_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3595 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3596 VSS a_768_44030# a_2711_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3597 a_n2216_40160# a_n2312_40392# a_n2302_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X3598 VSS a_14456_42282# a_5342_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3599 a_n984_44318# a_n2065_43946# a_n1331_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3600 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3601 a_11608_46482# a_n1151_42308# a_11387_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X3602 a_5093_45028# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3603 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3604 a_19862_44208# a_13747_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3605 VDD a_15227_44166# a_15597_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3606 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3607 a_19335_46494# a_18819_46122# a_19240_46482# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3608 VDD a_2324_44458# a_6298_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3609 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3610 a_8953_45546# a_8685_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3611 a_n4318_38216# a_n2472_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3612 a_18249_42858# a_18083_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3613 a_12816_46660# a_11735_46660# a_12469_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3614 a_19268_43646# a_13661_43548# a_19177_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.1525 ps=1.305 w=1 l=0.15
X3615 a_13258_32519# a_19647_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3616 a_20256_42852# a_20202_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3125 ps=1.625 w=1 l=0.15
X3617 VDD a_16680_45572# a_16855_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3618 VSS a_n447_43370# a_n2129_43609# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X3619 a_20528_45572# a_19466_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3620 a_11525_45546# a_10586_45546# a_11778_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X3621 VREF a_n3565_39590# C8_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3622 a_3537_45260# a_7287_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3623 VDD a_2711_45572# a_20107_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3624 a_16147_45260# a_17478_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3625 a_n2109_45247# a_n2017_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3626 a_19610_45572# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3627 a_19963_31679# a_22591_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3628 a_5837_43172# a_3537_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3629 a_n143_45144# a_n755_45592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3630 VDD a_18143_47464# a_12861_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X3631 VDD a_22959_47212# a_22612_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3632 a_n310_45572# a_n356_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X3633 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3634 VSS a_7227_47204# DATA[3] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3635 a_15015_46420# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3636 VSS a_7227_45028# a_7230_45938# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X3637 a_20596_44850# a_20159_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3638 a_2957_45546# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X3639 VSS a_14579_43548# a_14537_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3640 VDD a_n2946_39866# a_n3565_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3641 VDD a_11599_46634# a_15507_47210# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3642 VDD a_6151_47436# a_6812_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X3643 VSS a_5111_44636# a_8333_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3644 VDD a_7287_43370# a_3537_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X3645 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3646 VDD a_20679_44626# a_20640_44752# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3647 a_n3565_39304# a_n2946_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3648 VDD COMP_P a_n1329_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X3649 VSS a_19321_45002# a_20567_45036# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3650 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3651 a_14513_46634# a_14180_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X3652 a_10903_43370# a_13351_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3653 VSS a_n2472_45002# a_n2956_37592# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3654 a_10949_43914# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X3655 a_10149_43396# a_5111_44636# a_9803_43646# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3656 VSS a_19431_45546# a_19365_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3657 VSS a_16922_45042# a_17719_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X3658 a_16112_44458# a_14539_43914# a_16241_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3659 a_13943_43396# a_11823_42460# a_13837_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X3660 C8_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3661 VDD a_4099_45572# a_3483_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3662 a_6197_43396# a_6031_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3663 VSS a_18143_47464# a_12861_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X3664 a_n2840_46634# a_n2661_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3665 a_380_45546# a_n357_42282# a_603_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3666 a_18533_43940# a_18326_43940# a_18451_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3667 a_7309_42852# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X3668 VDD a_n863_45724# a_2448_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X3669 VSS a_1169_39587# COMP_P VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3670 a_5932_42308# a_5755_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3671 a_16328_43172# a_n97_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3672 VSS a_n2946_38778# a_n3565_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3673 a_17583_46090# a_17715_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X3674 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3675 VDD a_13635_43156# a_9290_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3676 VDD a_15433_44458# a_15463_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3677 a_n2267_43396# a_n2433_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3678 VDD a_n755_45592# a_8147_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X3679 VSS a_10991_42826# a_10922_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X3680 a_5732_46660# a_4651_46660# a_5385_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3681 a_19615_44636# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X3682 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X3683 VDD a_5129_47502# a_5159_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3684 a_n2840_46090# a_n2661_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3685 a_n967_45348# a_n913_45002# a_n955_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3686 a_19006_44850# a_18248_44752# a_18443_44721# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X3687 a_n4209_39590# a_n2302_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X3688 VDD a_18817_42826# a_18707_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3689 a_15559_46634# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X3690 a_9803_43646# a_8953_45546# a_9885_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3691 VDD a_3232_43370# a_9313_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X3692 VDD a_n2840_42282# a_n3674_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3693 a_13460_43230# a_12545_42858# a_13113_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3694 a_20362_44736# a_20679_44626# a_20637_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X3695 a_2713_42308# a_n913_45002# a_2725_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3696 a_768_44030# a_13487_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3697 a_16241_47178# a_16023_47582# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3698 a_14955_43396# a_14205_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X3699 VSS a_n913_45002# a_10533_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3700 a_7466_43396# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3701 a_n4064_40160# a_n4334_40480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3702 VDD a_6151_47436# a_5907_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3703 a_16697_47582# a_15507_47210# a_16588_47582# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3704 a_n2267_44484# a_n2433_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3705 a_15682_43940# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3706 a_13693_46688# a_6755_46942# a_13607_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3707 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3708 a_19250_35138# VDD EN_VIN_BSTR_N VSS sky130_fd_pr__nfet_05v0_nvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.9
X3709 VDAC_Ni a_3754_38470# a_3726_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3710 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3711 VDD a_19778_44110# a_19741_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3712 VSS a_n1794_35242# a_n1696_35090# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3713 a_2609_46660# a_2443_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3714 a_5708_44484# a_5257_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X3715 a_18143_47464# a_18479_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X3716 a_5263_46660# a_4817_46660# a_5167_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3717 VSS a_n2472_43914# a_n3674_39768# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3718 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3719 a_12016_45572# a_11962_45724# a_11525_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3720 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3721 VSS a_1107_38525# a_1273_38525# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3722 VSS a_18057_42282# a_n356_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X3723 VDD a_21671_42860# a_3422_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3724 VDD a_8746_45002# a_8704_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X3725 C9_N_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3726 a_3411_47243# a_3160_47472# a_2952_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3727 a_n2840_46634# a_n2661_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3728 VSS a_7705_45326# a_7639_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X3729 VSS a_167_45260# a_1423_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3730 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3731 VDD a_9396_43370# a_5111_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3732 a_743_42282# a_13661_43548# a_20301_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3733 a_n3420_39616# a_n3690_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3734 a_133_43172# a_n357_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X3735 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3736 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3737 VSS a_n2946_37690# a_n3565_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3738 VDD a_20512_43084# a_19987_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
X3739 a_1891_43646# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.14825 ps=1.34 w=0.42 l=0.15
X3740 VSS a_526_44458# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3741 a_14485_44260# a_5807_45002# a_12465_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3742 a_n4318_39304# a_n2840_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3743 VIN_P EN_VIN_BSTR_P C8_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3744 VSS a_n357_42282# a_17141_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3745 a_11453_44696# a_17719_45144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
X3746 VSS a_n1059_45260# a_8945_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3747 a_17701_42308# a_17531_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3748 a_13657_42558# a_11823_42460# a_13575_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3749 a_10545_42558# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3750 a_8292_43218# a_7765_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3751 a_16751_46987# a_5807_45002# a_16292_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3752 a_10586_45546# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3753 a_n1243_44484# a_n2433_44484# a_n1352_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3754 VSS a_16855_45546# a_16789_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3755 a_45_45144# a_n143_45144# a_n37_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3756 VDD a_3537_45260# a_4223_44672# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3757 a_3626_43646# a_1414_42308# a_3540_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3758 VSS a_n2946_37984# a_n3565_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3759 VDD a_20107_42308# a_7174_31319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3760 a_3815_47204# a_3785_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3761 a_n1917_44484# a_n2267_44484# a_n2012_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3762 VCM a_5342_30871# C8_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3763 a_15567_42826# a_15743_43084# a_15953_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3764 VSS a_10341_42308# a_11554_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X3765 VSS a_4791_45118# a_6640_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X3766 a_6755_46942# a_15015_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X3767 a_2437_43646# a_1568_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3768 VDAC_Pi a_7754_39632# VSS sky130_fd_pr__res_high_po_0p35 l=18
X3769 a_n3420_38528# a_n3690_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3770 a_n4209_39590# a_n2302_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3771 a_9823_46155# a_9804_47204# a_9823_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3772 a_1990_45899# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3773 a_15743_43084# a_19339_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X3774 a_5129_47502# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3775 VDD a_5385_46902# a_5275_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3776 a_9145_43396# a_8791_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X3777 VDD a_20841_46902# a_20731_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3778 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3779 VIN_P EN_VIN_BSTR_P C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3780 VDD a_n785_47204# a_327_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3781 a_7276_45260# a_n1151_42308# a_7418_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3782 a_8103_44636# a_8375_44464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3783 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3784 a_4915_47217# a_12991_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X3785 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3786 VDD a_8199_44636# a_8855_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X3787 VDD a_12549_44172# a_21115_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3788 VDD a_2553_47502# a_2583_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3789 a_n327_42558# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X3790 a_12800_43218# a_12089_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3791 VSS a_20623_43914# a_20365_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X3792 VSS a_n743_46660# a_16501_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X3793 VSS a_22959_45036# a_19721_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3794 VSS a_11967_42832# a_16243_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3795 VDD a_7754_40130# a_11206_38545# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3796 a_n4318_38680# a_n2472_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3797 a_3363_44484# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3798 a_13483_43940# a_13249_42308# a_13565_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3799 a_7754_40130# RST_Z VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3800 VDD a_4235_43370# a_n2661_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3801 a_n4209_38502# a_n2302_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3802 a_13249_42558# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X3803 a_18504_43218# a_17333_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3804 a_n39_42308# a_n97_42460# a_n473_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3805 a_10210_45822# a_10180_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X3806 VSS a_11967_42832# a_20512_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3807 VSS a_n443_46116# a_2813_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3808 VSS a_4646_46812# a_7411_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3809 a_20273_46660# a_20107_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3810 VDD a_11341_43940# a_22223_43948# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3811 a_n2312_38680# a_n2104_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3812 VDD a_12791_45546# a_12427_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X3813 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3814 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X3815 a_19237_31679# a_22959_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3816 VDD a_19328_44172# a_19279_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16675 pd=1.435 as=0.26 ps=2.52 w=1 l=0.15
X3817 VIN_N EN_VIN_BSTR_N a_11530_34132# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3818 VDD SMPL_ON_P a_n1605_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3819 VSS a_11967_42832# a_12379_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3820 VSS a_15227_44166# a_17719_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3821 VDD a_18315_45260# a_18189_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X3822 a_10951_45334# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X3823 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3824 VDD a_2123_42473# a_1184_42692# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3825 a_4791_45118# a_4743_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X3826 a_21753_35634# a_19998_35138# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3827 a_21195_42852# a_20922_43172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25675 ps=1.44 w=0.65 l=0.15
X3828 a_4156_43218# a_3905_42865# a_3935_42891# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X3829 a_15227_44166# a_22000_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3830 a_n3420_37440# a_n3690_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3831 a_n1899_43946# a_n2065_43946# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3832 VDD a_17591_47464# a_16327_47482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X3833 a_n743_46660# a_n1021_46688# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3834 a_n2293_45546# a_2274_45254# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X3835 a_11633_42308# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3836 a_15682_46116# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3837 a_20205_31679# a_22223_46124# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3838 a_n2472_46634# a_n2293_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3839 a_2698_46116# a_2521_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3840 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X3841 VDD a_10193_42453# a_11682_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X3842 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3843 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3844 VDD a_n3565_38502# a_n3690_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X3845 a_5342_30871# a_14456_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3846 VDD a_8325_42308# a_8791_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3847 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3848 a_548_43396# a_n863_45724# a_458_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X3849 VDD a_n4334_39616# a_n4064_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X3850 VSS a_1756_43548# a_1467_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.182 ps=1.86 w=0.65 l=0.15
X3851 a_288_46660# a_171_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3852 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3853 VDD a_17517_44484# a_22591_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3854 VSS a_n913_45002# a_19511_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3855 a_20894_47436# a_20990_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3856 a_15312_46660# a_14976_45028# a_15009_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X3857 a_n2472_46090# a_n2293_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3858 VDD a_n2438_43548# a_n2157_46122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3859 VSS a_22959_43948# a_17538_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3860 C9_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X3861 VDD a_n4064_38528# a_n2216_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X3862 a_8037_42858# a_7871_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3863 a_n1736_43218# a_n1853_43023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3864 a_n4209_37414# a_n2302_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3865 a_13527_45546# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3866 VDD a_n2472_42282# a_n4318_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3867 a_n2661_43370# a_11415_45002# a_11361_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3868 VSS a_1273_38525# a_2113_38308# VSS sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X3869 VDD a_22165_42308# a_22223_42860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3870 VDD a_n2840_42826# a_n3674_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3871 VSS a_14180_45002# a_13017_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X3872 a_15681_43442# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3873 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3874 C8_N_btm a_21076_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3875 VSS a_n2302_40160# a_n4315_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3876 a_8488_45348# a_8199_44636# a_8191_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X3877 a_16588_47582# a_15673_47210# a_16241_47178# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3878 a_18220_42308# a_18184_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X3879 a_n1423_46090# a_n1641_46494# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3880 EN_VIN_BSTR_N VDD a_19250_35138# VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.9
X3881 VSS a_n4334_38528# a_n4064_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X3882 VDD a_18143_47464# a_12861_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3883 a_17609_46634# a_12549_44172# a_18280_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3884 a_16115_45572# a_15599_45572# a_16020_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3885 VSS a_19700_43370# a_n97_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3886 VSS a_2124_47436# a_1209_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X3887 VREF_GND a_17730_32519# C9_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3888 a_15595_45028# a_15415_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X3889 VDD a_6755_46942# a_12741_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3890 VSS a_19615_44636# a_18579_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X3891 a_12545_42858# a_12379_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3892 a_16942_47570# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3893 a_8791_45572# a_7499_43078# a_8697_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3894 a_14853_42852# a_n913_45002# a_14635_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3895 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3896 a_8333_44056# a_4223_44672# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3897 VSS a_4958_30871# a_17531_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3898 a_6511_45714# a_4646_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3899 VDD a_10949_43914# a_10867_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X3900 a_17973_43940# a_17737_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X3901 a_18494_42460# a_18907_42674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X3902 a_17061_44734# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X3903 a_n2472_46634# a_n2293_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3904 C2_P_btm a_3080_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X3905 VSS a_5267_42460# a_4905_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X3906 VSS a_n2438_43548# a_n2065_43946# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3907 VDD a_7754_40130# a_3754_38470# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3908 a_22629_38406# a_22537_39537# CAL_N VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3909 VDD a_n357_42282# a_5837_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3910 a_9159_45572# a_5937_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X3911 a_3483_46348# a_4099_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3912 a_8238_44734# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X3913 VSS a_17517_44484# a_22591_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3914 VDD a_n3565_37414# a_n3690_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X3915 VDD a_3381_47502# a_3411_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3916 VSS a_21613_42308# a_22775_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X3917 COMP_P a_1169_39587# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3918 a_10150_46912# a_10467_46802# a_10425_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X3919 a_526_44458# a_3147_46376# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3920 a_n2810_45572# a_n2840_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3921 a_13675_47204# a_n1435_47204# a_13569_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X3922 VSS a_11827_44484# a_22223_45036# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3923 a_5518_44484# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X3924 VDD a_n4064_37440# a_n2216_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X3925 a_22165_42308# a_21887_42336# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X3926 a_n3565_38502# a_n2946_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X3927 a_5891_43370# a_9127_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3928 a_13678_32519# a_21855_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3929 a_n2312_40392# a_n2288_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3930 VDD a_8605_42826# a_8495_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3931 a_7499_43078# a_10083_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3932 VDD a_20193_45348# a_21887_42336# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3933 a_18691_45572# a_18341_45572# a_18596_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3934 a_13076_44458# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X3935 w_1575_34946# a_n1696_35090# EN_VIN_BSTR_P w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X3936 a_3600_43914# a_1307_43914# a_3992_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X3937 VSS a_n4334_37440# a_n4064_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X3938 a_4743_43172# a_3537_45260# a_4649_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3939 a_11387_46155# a_11309_47204# a_11387_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3940 a_n755_45592# a_n809_44244# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3941 a_15682_43940# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3942 VDD a_1666_39587# a_1169_39587# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3943 a_n1177_44458# a_n1352_44484# a_n998_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3944 a_11554_42852# a_10835_43094# a_10991_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X3945 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3946 VDD a_2680_45002# a_2274_45254# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X3947 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3948 VSS a_9313_44734# a_22959_42860# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3949 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3950 VDD a_n1177_43370# a_n1190_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3951 w_1575_34946# a_n1057_35174# w_1575_34946# w_1575_34946# sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=0 ps=0 w=3.75 l=15
X3952 VDD a_6755_46942# a_13556_45296# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3953 a_n785_47204# a_n815_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3954 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3955 VDD a_n971_45724# a_8147_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X3956 a_n1696_35090# a_n1794_35242# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3957 a_n4251_40480# a_n4318_40392# a_n4334_40480# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X3958 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3959 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3960 a_19900_46494# a_18819_46122# a_19553_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3961 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3962 a_12359_47026# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3963 a_12561_45572# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1034 ps=1 w=0.42 l=0.15
X3964 a_10083_42826# a_10518_42984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X3965 VSS a_10355_46116# a_8199_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3966 a_3422_30871# a_21671_42860# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3967 a_5937_45572# a_5907_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3968 a_21005_45260# a_21101_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X3969 VDD a_16327_47482# a_17767_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3970 a_12649_45572# a_10903_43370# a_12561_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X3971 VSS a_19321_45002# a_19113_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3972 a_5111_44636# a_9396_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3973 VSS a_18194_35068# a_11530_34132# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3974 a_12469_46902# a_12251_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3975 a_21297_45572# a_20107_45572# a_21188_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3976 a_376_46348# a_584_46384# a_518_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3977 a_15146_44484# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X3978 VIN_P EN_VIN_BSTR_P C6_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X3979 VDD a_n971_45724# a_n327_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X3980 a_n3565_37414# a_n2946_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X3981 a_14180_45002# a_14537_43396# a_14309_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3982 VDD a_10193_42453# a_16237_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3983 a_18681_44484# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X3984 VSS a_15009_46634# a_14180_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X3985 a_17829_46910# a_12549_44172# a_765_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1525 ps=1.305 w=1 l=0.15
X3986 a_2304_45348# a_2274_45254# a_2232_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X3987 VDD a_1169_39043# comp_n VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3988 a_6598_45938# a_6511_45714# a_6194_45824# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X3989 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3990 a_n3565_38216# a_n2946_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3991 a_5745_43940# a_5013_44260# a_5663_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3992 VDD a_10193_42453# a_18533_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3993 a_5742_30871# a_10723_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3994 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3995 a_19478_44056# a_3090_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.16675 ps=1.435 w=0.42 l=0.15
X3996 VSS a_15051_42282# a_11823_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3997 a_10185_46660# a_10150_46912# a_9863_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X3998 a_8192_45572# a_8199_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X3999 a_15890_42674# a_15764_42576# a_15486_42560# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X4000 a_10835_43094# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4001 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4002 a_n699_43396# a_n1177_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X4003 a_14033_45822# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X4004 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4005 a_6101_44260# a_1307_43914# a_5663_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4006 a_7927_46660# a_7577_46660# a_7832_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4007 a_21496_47436# a_4883_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X4008 a_16721_46634# a_16388_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4009 a_5826_44734# a_5147_45002# a_5518_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X4010 VDD a_16763_47508# a_16750_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4011 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4012 VDD a_n746_45260# a_175_44278# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X4013 a_n443_46116# a_n901_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4014 a_2813_43396# a_3232_43370# a_2982_43646# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4015 a_6171_42473# a_5932_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4016 VDD a_601_46902# a_491_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X4017 VSS a_4646_46812# a_6031_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4018 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4019 VDD a_1123_46634# a_1110_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4020 VSS a_13059_46348# a_12638_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X4021 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4022 a_11787_45002# a_11963_45334# a_11915_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X4023 VSS a_584_46384# a_2998_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4024 a_8292_43218# a_7765_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4025 VDD a_n2472_42826# a_n4318_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4026 a_1667_45002# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X4027 VDD a_n3690_38528# a_n3420_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4028 a_20731_47026# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X4029 a_8062_46482# a_8016_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4030 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4031 a_n2216_38778# a_n2312_38680# a_n2302_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X4032 VSS a_11599_46634# a_20107_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4033 a_13925_46122# a_13759_46122# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4034 VSS CLK a_8953_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4035 VSS a_n2104_46634# a_n2312_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4036 a_5385_46902# a_5167_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4037 a_n1177_44458# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4038 VDD a_7499_43078# a_10729_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X4039 a_9803_43646# a_8953_45546# a_9885_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4040 VDD a_19256_45572# a_19431_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4041 a_7911_44260# a_7845_44172# a_7542_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.182 ps=1.86 w=0.65 l=0.15
X4042 VDD a_5111_44636# a_7542_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X4043 VDD a_6761_42308# a_7227_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X4044 VDD a_19553_46090# a_19443_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X4045 a_n1641_43230# a_n2157_42858# a_n1736_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4046 a_5205_44484# a_5343_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4047 a_22400_42852# a_22223_42860# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4048 a_12603_44260# a_12549_44172# a_12495_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.12675 ps=1.04 w=0.65 l=0.15
X4049 a_3638_45822# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X4050 a_17324_43396# a_16243_43396# a_16977_43638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X4051 a_19452_47524# a_19386_47436# a_13747_46662# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4052 a_5275_47026# a_4651_46660# a_5167_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4053 VSS a_327_47204# DATA[0] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4054 a_11915_45394# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X4055 a_14447_46660# a_n1151_42308# a_14084_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4056 a_20731_47026# a_20107_46660# a_20623_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4057 VSS a_n1613_43370# a_n1655_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4058 a_12800_43218# a_12089_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4059 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4060 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4061 VSS a_20712_42282# a_10193_42453# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4062 a_15720_42674# a_15051_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4063 VSS a_n443_42852# a_421_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X4064 a_14493_46090# a_14275_46494# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4065 VDD a_11599_46634# a_15599_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4066 a_n659_45366# a_n746_45260# a_n745_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4067 a_15682_46116# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X4068 a_n881_46662# a_14495_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X4069 a_8685_43396# a_8147_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X4070 C7_P_btm a_n4209_39304# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4071 a_765_45546# a_17609_46634# a_17639_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4072 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X4073 a_11554_42852# a_10796_42968# a_10991_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X4074 a_19386_47436# a_19321_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4075 a_8492_46660# a_7411_46660# a_8145_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X4076 a_2063_45854# a_9863_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4077 VDD a_15803_42450# a_15764_42576# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4078 a_1337_46436# a_1176_45822# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4079 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4080 VSS a_4419_46090# a_4365_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4081 a_n1549_44318# a_n1899_43946# a_n1644_44306# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4082 VDD a_9067_47204# DATA[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4083 VSS a_6575_47204# a_9067_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X4084 a_n1331_43914# a_n1549_44318# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4085 VDD a_3537_45260# a_5093_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X4086 VSS a_11189_46129# a_11608_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X4087 a_20835_44721# a_20640_44752# a_21145_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X4088 a_n327_42558# a_n97_42460# a_n473_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X4089 a_8147_43396# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X4090 VDD a_n3690_37440# a_n3420_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4091 a_19431_46494# a_18985_46122# a_19335_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4092 VDD a_12607_44458# a_n2661_43922# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4093 VDD a_17324_43396# a_17499_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4094 a_8685_42308# a_8515_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4095 a_1414_42308# a_1067_42314# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X4096 VDD a_4883_46098# a_10355_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4097 a_n2216_37690# a_n2810_45028# a_n2302_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X4098 VDD a_10193_42453# a_9885_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4099 VDD a_21356_42826# a_n357_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4100 a_16977_43638# a_16759_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4101 VSS a_n4334_40480# a_n4064_40160# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4102 VSS a_n237_47217# a_8270_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4103 a_10555_43940# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4104 a_1049_43396# a_458_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4105 EN_VIN_BSTR_P VDD a_n217_35174# VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.9
X4106 VSS a_22775_42308# a_22485_38105# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4107 VDD a_n443_42852# a_742_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4108 a_8145_46902# a_7927_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4109 a_21613_42308# a_21335_42336# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X4110 VDD a_n23_45546# a_7_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4111 VSS a_16019_45002# a_15903_45785# VSS sky130_fd_pr__nfet_01v8 ad=0.160875 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X4112 VCM a_5342_30871# C8_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4113 VDD a_2698_46116# a_2804_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X4114 a_20935_43940# a_18479_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4115 a_2713_42308# a_n755_45592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4116 VDD a_n699_43396# a_4743_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4117 DATA[1] a_1431_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4118 a_17591_47464# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X4119 a_9223_42460# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X4120 a_12741_44636# a_14537_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4121 a_2684_37794# a_1666_39587# a_1666_39043# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4122 VDD a_20202_43084# a_21335_42336# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X4123 a_564_42282# a_743_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4124 a_15367_44484# a_13556_45296# a_15004_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4125 VSS a_n2302_40160# a_n4315_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4126 VSS a_n452_47436# a_n815_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4127 VDD a_2063_45854# a_9863_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X4128 a_2981_46116# a_2804_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X4129 VSS a_6511_45714# a_6472_45840# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4130 VSS a_13159_45002# a_13105_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4131 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4132 a_9223_42460# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4133 VSS a_19987_42826# a_n2017_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.08775 ps=0.92 w=0.65 l=0.15
X4134 a_20692_30879# a_22959_46124# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4135 a_21188_45572# a_20273_45572# a_20841_45814# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4136 a_9028_43914# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X4137 VDD a_17715_44484# a_17737_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4138 VSS a_n2840_44458# a_n4318_40392# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4139 VSS a_15004_44636# a_14815_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4140 a_16759_43396# a_16243_43396# a_16664_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4141 a_4574_45260# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X4142 a_17829_46910# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4143 VSS a_n443_46116# a_4880_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X4144 a_n4064_38528# a_n4334_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4145 VDD a_1799_45572# a_1983_46706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X4146 VDD a_21363_45546# a_21350_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4147 a_n4064_40160# a_n4334_40480# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X4148 VDD a_22775_42308# a_22485_38105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4149 a_13259_45724# a_17583_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4150 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4151 C1_P_btm a_n4064_37440# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4152 VIN_P EN_VIN_BSTR_P C4_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X4153 a_6575_47204# a_6545_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4154 VSS a_765_45546# a_380_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X4155 VSS a_327_44734# a_501_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4156 a_104_43370# a_n699_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4157 VDD a_22959_42860# a_14097_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4158 a_n2293_42282# a_3357_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4159 VSS a_6171_42473# a_5379_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4160 a_3935_42891# a_2382_45260# a_3935_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4161 VSS a_9067_47204# DATA[4] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4162 VDD a_8145_46902# a_8035_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X4163 VDD a_n863_45724# a_327_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X4164 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4165 a_17141_43172# a_n1059_45260# a_16795_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4166 VDD a_9127_43156# a_5891_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4167 a_15433_44458# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4168 VSS a_10193_42453# a_11897_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X4169 VSS a_4791_45118# a_5066_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4170 VDD a_5691_45260# a_n2109_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X4171 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X4172 VDD a_1983_46706# a_n2661_46098# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4173 a_15227_46910# a_15368_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4174 a_18753_44484# a_18374_44850# a_18681_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X4175 a_15486_42560# a_15803_42450# a_15761_42308# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X4176 a_n1641_43230# a_n1991_42858# a_n1736_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4177 a_6682_46987# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X4178 a_n1079_45724# a_n755_45592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X4179 a_12429_44172# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.118125 ps=1.04 w=0.42 l=0.15
X4180 a_1568_43370# a_1847_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4181 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X4182 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4183 VDD a_7227_42308# a_6123_31319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4184 VSS a_1123_46634# a_584_46384# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4185 a_3457_43396# a_3232_43370# a_3626_43646# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4186 a_7174_31319# a_20107_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4187 a_8952_43230# a_8037_42858# a_8605_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4188 VSS a_167_45260# a_n37_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4189 a_13490_45067# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X4190 a_4181_44734# a_3090_45724# a_n2497_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4191 VSS a_6171_45002# a_11909_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4192 VSS a_n2302_39866# a_n4209_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4193 a_33_46660# a_n133_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4194 a_16388_46812# a_17957_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.112125 ps=0.995 w=0.65 l=0.15
X4195 VDD a_3218_45724# a_3175_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4196 a_8283_46482# a_n1151_42308# a_7920_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4197 a_8953_45002# CLK VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4198 VSS a_n809_44244# a_n755_45592# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4199 VDD a_15279_43071# a_14579_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4200 VDD a_16763_47508# a_5807_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4201 VDD a_310_45028# a_509_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X4202 a_n23_47502# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4203 a_n1099_45572# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X4204 VDD a_10903_43370# a_10907_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X4205 a_3935_43218# a_3681_42891# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X4206 a_14949_46494# a_13759_46122# a_14840_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4207 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4208 a_6851_47204# a_6491_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4209 a_13556_45296# a_6755_46942# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4210 VDD a_n4315_30879# a_n4334_40480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X4211 VSS a_15227_44166# a_14539_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X4212 a_19987_42826# a_18494_42460# a_20356_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
X4213 a_n2833_47464# a_n2497_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X4214 a_3524_46660# a_2609_46660# a_3177_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4215 VSS a_n1696_35090# a_n217_35174# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X4216 a_n4209_39304# a_n2302_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X4217 VSS a_22223_47212# a_21588_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4218 VSS a_6151_47436# a_6229_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X4219 a_18533_43940# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X4220 a_14205_43396# a_13667_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X4221 VREF a_n3565_39590# C8_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4222 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4223 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4224 a_n4064_37440# a_n4334_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4225 a_16377_45572# a_16333_45814# a_16211_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X4226 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X4227 a_10044_46482# a_n743_46660# a_9823_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4228 a_19113_45348# a_18911_45144# a_3090_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4229 VSS a_13720_44458# a_12607_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X4230 a_n2860_37984# a_n2956_38216# a_n2946_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X4231 a_2266_47570# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4232 a_5837_43396# a_5111_44636# a_5147_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4233 a_5934_30871# a_8791_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4234 a_10861_46660# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X4235 VSS a_7920_46348# a_7715_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4236 a_14383_46116# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X4237 a_2809_45348# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4238 a_2905_42968# a_742_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4239 a_6540_46812# a_6755_46942# a_6682_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X4240 a_6709_45028# a_6431_45366# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X4241 a_8953_45002# CLK VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4242 VSS a_18494_42460# a_20193_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4243 a_n2442_46660# a_n2472_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4244 C7_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X4245 a_13249_42308# a_13070_42354# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X4246 a_n1991_42858# a_n2157_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4247 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X4248 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4249 a_13348_45260# a_12891_46348# a_13490_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X4250 w_11334_34010# a_11530_34132# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.54375 pd=4.04 as=0 ps=0 w=3.75 l=15
X4251 VREF_GND a_n4064_39616# C9_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4252 a_17061_44484# a_11691_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4253 comp_n a_1169_39043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4254 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X4255 VDD a_18443_44721# a_18374_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X4256 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4257 a_1512_43396# a_n443_46116# a_1209_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X4258 VDD a_n3565_39304# a_n3690_39392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X4259 VDD a_22591_44484# a_17730_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4260 VDD a_22581_37893# a_22537_39537# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4261 VSS a_15803_42450# a_15764_42576# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4262 a_11901_46660# a_11735_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4263 EN_VIN_BSTR_N a_18194_35068# w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X4264 a_21076_30879# a_22959_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4265 a_3877_44458# a_3699_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X4266 VDD a_n4064_39072# a_n2216_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X4267 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4268 a_11691_44458# a_5807_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4269 a_15368_46634# a_15143_45578# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X4270 VSS a_9028_43914# a_8975_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X4271 a_2813_43396# a_n443_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X4272 C8_N_btm a_17538_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4273 a_5093_45028# a_4558_45348# a_5009_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4274 VSS a_10193_42453# a_13921_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X4275 a_15597_42852# a_15567_42826# a_15095_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X4276 a_2553_47502# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4277 VDD a_13059_46348# a_12839_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4278 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4279 a_3823_42558# a_3065_45002# a_3905_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X4280 VDD a_526_44458# a_5193_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4281 VSS a_1667_45002# a_n863_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X4282 a_1307_43914# a_2779_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4283 VDD a_n3690_38528# a_n3420_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X4284 VDD a_21177_47436# a_20990_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X4285 a_16855_45546# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4286 a_5495_43940# a_5244_44056# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X4287 VDD a_5815_47464# a_n1613_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X4288 VSS a_19787_47423# a_19594_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4289 VDD a_22365_46825# a_20202_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4290 a_5063_47570# a_4915_47217# a_4700_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4291 a_n1736_46482# a_n1853_46287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4292 VDD a_11459_47204# DATA[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X4293 a_11322_45546# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4294 a_19787_47423# START VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4295 a_3754_39466# a_7754_39632# VSS sky130_fd_pr__res_high_po_0p35 l=18
X4296 a_n4251_39616# a_n4318_39768# a_n4334_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X4297 VDD a_9127_43156# a_9114_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4298 a_10384_47026# a_9863_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4299 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X4300 VSS a_11525_45546# a_11189_46129# VSS sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X4301 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4302 a_10729_43914# a_11750_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4303 a_4921_42308# a_n913_45002# a_4933_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4304 VSS a_n23_47502# a_n89_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4305 a_20528_46660# a_20411_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4306 VSS a_8568_45546# a_8162_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X4307 a_13657_42558# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X4308 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X4309 VSS a_4223_44672# a_5205_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4310 a_18005_44484# a_17970_44736# a_17767_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X4311 a_13837_43396# a_13259_45724# a_13749_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X4312 a_19177_43646# a_17339_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X4313 a_196_42282# a_375_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4314 a_791_42968# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4315 VSS a_327_47204# DATA[0] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4316 a_11309_47204# a_11031_47542# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X4317 VSS a_4646_46812# a_7871_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4318 VSS a_5815_47464# a_n1613_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X4319 a_n23_45546# a_n356_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X4320 a_18691_45572# a_18175_45572# a_18596_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4321 a_9885_42558# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X4322 VSS a_4700_47436# a_3785_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4323 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X4324 a_4361_42308# a_3823_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X4325 VDD a_n2840_46634# a_n2956_39768# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4326 a_4817_46660# a_4651_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4327 VDD a_13635_43156# a_13622_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4328 VDD a_n2438_43548# a_n2157_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4329 a_8415_44056# a_5343_44458# a_8333_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4330 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4331 VSS a_1307_43914# a_4156_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X4332 a_n1699_44726# a_n1917_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4333 a_1525_44260# a_1467_44172# a_1115_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X4334 VDD a_n2946_39866# a_n3565_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4335 a_14976_45028# a_14797_45144# a_15060_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X4336 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X4337 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4338 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X4339 a_n3565_39304# a_n2946_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X4340 VSS a_15959_42545# a_15890_42674# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X4341 a_n2312_39304# a_n1920_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X4342 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4343 VIN_N EN_VIN_BSTR_N C7_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X4344 VDD a_1666_39587# a_1666_39043# VDD sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X4345 VDD a_n3690_37440# a_n3420_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X4346 VSS a_21363_45546# a_21297_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4347 VDD a_n452_44636# a_n2129_44697# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X4348 a_19443_46116# a_18819_46122# a_19335_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4349 VDD a_7112_43396# a_7287_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4350 VSS a_21753_35634# SMPL_ON_N VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4351 a_310_45028# a_n37_45144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X4352 VDD a_5111_44636# a_5518_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X4353 VDD EN_VIN_BSTR_N w_11334_34010# w_11334_34010# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4354 a_17719_45144# a_17613_45144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X4355 a_17499_43370# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4356 VDD a_12563_42308# a_5534_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4357 VSS a_13747_46662# a_19466_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4358 a_14112_44734# a_768_44030# a_13857_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X4359 VSS a_n2946_38778# a_n3565_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4360 a_n357_42282# a_21356_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4361 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X4362 VDD a_3483_46348# a_15037_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4363 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4364 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X4365 VDD a_13635_43156# a_9290_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X4366 VDD a_13487_47204# a_768_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4367 a_14097_32519# a_22959_42860# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4368 a_3094_47570# a_2905_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4369 a_8270_45546# a_n237_47217# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4370 a_8781_46436# a_8199_44636# a_8034_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4371 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4372 VSS a_3232_43370# a_11541_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X4373 DATA[4] a_9067_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X4374 a_20841_46902# a_20623_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4375 a_13527_45546# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4376 a_10533_42308# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4377 a_17896_45144# a_16922_45042# a_17801_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
X4378 DATA[1] a_1431_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X4379 a_18817_42826# a_18599_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4380 a_104_43370# a_n699_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X4381 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4382 a_16211_45572# a_15765_45572# a_16115_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4383 VDD a_4223_44672# a_4181_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4384 VSS a_20835_44721# a_20766_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X4385 a_19741_43940# a_19478_44306# a_19328_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4386 VDD a_13747_46662# a_14495_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4387 a_2487_47570# a_2063_45854# a_2124_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4388 VSS a_10809_44734# a_22959_46124# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4389 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4390 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4391 VSS a_7754_38470# a_6886_37412# VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4392 VSS a_20567_45036# a_12549_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4393 a_21359_45002# a_21513_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4394 a_18451_43940# a_18579_44172# a_18533_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X4395 a_13904_45546# a_13249_42308# a_14033_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X4396 VSS a_13661_43548# a_18587_45118# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4397 a_6547_43396# a_6031_43396# a_6452_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
C0 a_13467_32519# VDD 0.353373f
C1 a_20273_46660# VDD 0.247553f
C2 a_19321_45002# a_11967_42832# 0.266816f
C3 a_5937_45572# a_7229_43940# 0.126047f
C4 a_13259_45724# a_15861_45028# 0.16873f
C5 a_11599_46634# a_15507_47210# 0.267808f
C6 a_12861_44030# a_16327_47482# 0.120085f
C7 a_n971_45724# a_n1613_43370# 0.6298f
C8 a_3090_45724# a_19328_44172# 0.153704f
C9 a_15227_44166# a_14955_43940# 0.134177f
C10 a_20273_45572# a_21188_45572# 0.125324f
C11 C6_P_btm C0_P_btm 0.139059f
C12 C5_P_btm C1_P_btm 0.127408f
C13 C4_P_btm C2_P_btm 7.72909f
C14 a_12549_44172# a_6755_46942# 0.553062f
C15 a_n971_45724# a_n2293_46098# 0.110318f
C16 a_4883_46098# a_15227_44166# 0.176028f
C17 a_n1550_35608# VDD 0.366274f
C18 EN_VIN_BSTR_N C6_N_btm 0.118916f
C19 C7_P_btm C0_dummy_P_btm 0.119061f
C20 a_22315_44484# VDD 0.213791f
C21 a_7499_43078# a_8685_43396# 0.153217f
C22 a_10057_43914# a_5891_43370# 0.197199f
C23 a_n2109_47186# VDD 2.71791f
C24 a_n755_45592# a_3318_42354# 0.152654f
C25 a_310_45028# a_n356_45724# 0.12349f
C26 a_584_46384# a_2553_47502# 0.100103f
C27 a_n3565_39590# a_n3690_39616# 0.246863f
C28 a_22537_40625# a_22527_39145# 0.245895f
C29 a_n1613_43370# a_601_46902# 0.178721f
C30 a_5807_45002# a_19321_45002# 0.376188f
C31 a_3357_43084# SINGLE_ENDED 0.131897f
C32 a_22959_45572# VDD 0.304443f
C33 a_13348_45260# a_9482_43914# 0.352976f
C34 a_13017_45260# a_13777_45326# 0.195607f
C35 a_526_44458# a_n2661_42282# 0.191497f
C36 a_11901_46660# a_12251_46660# 0.219633f
C37 a_11735_46660# a_12816_46660# 0.102325f
C38 a_10835_43094# a_10991_42826# 0.105839f
C39 a_11691_44458# a_15004_44636# 0.221929f
C40 a_n971_45724# a_3429_45260# 0.171338f
C41 a_n2109_47186# a_5691_45260# 0.113268f
C42 a_19319_43548# VDD 0.561461f
C43 a_4185_45028# a_17303_42282# 0.235259f
C44 a_n1925_46634# VDD 0.783093f
C45 a_6109_44484# a_6453_43914# 0.165572f
C46 a_16327_47482# a_18287_44626# 0.552724f
C47 a_12549_44172# a_20193_45348# 0.587618f
C48 a_11415_45002# a_8696_44636# 0.10924f
C49 a_16795_42852# VDD 0.179044f
C50 a_n2956_38216# a_n3420_37984# 0.208204f
C51 a_10355_46116# VDD 0.222751f
C52 a_n2810_45572# a_n2302_37984# 0.130495f
C53 a_20692_30879# a_20447_31679# 9.02991f
C54 a_584_46384# a_1799_45572# 0.179456f
C55 a_4958_30871# VCM 0.642743f
C56 a_21335_42336# VDD 0.199586f
C57 a_7174_31319# RST_Z 0.216004f
C58 a_11599_46634# a_13747_46662# 0.25325f
C59 a_7411_46660# a_7715_46873# 0.162909f
C60 a_5807_45002# a_13059_46348# 0.1145f
C61 a_n971_45724# a_6945_45028# 0.247957f
C62 a_n1423_42826# a_n1641_43230# 0.209641f
C63 a_1307_43914# a_14539_43914# 0.131617f
C64 a_22365_46825# a_20202_43084# 0.115624f
C65 a_10949_43914# VDD 0.797824f
C66 a_20894_47436# VDD 0.188358f
C67 a_13661_43548# a_9482_43914# 0.127225f
C68 a_n2293_46098# a_2711_45572# 0.530463f
C69 a_17583_46090# a_13259_45724# 0.191869f
C70 a_13059_46348# a_15143_45578# 0.262261f
C71 a_n2293_42834# a_n2472_42826# 0.199703f
C72 a_20411_46873# VDD 0.348821f
C73 a_13259_45724# a_8696_44636# 0.259609f
C74 a_n4064_38528# a_n2302_38778# 0.239588f
C75 a_20107_45572# a_21188_45572# 0.102355f
C76 a_20841_45814# a_20623_45572# 0.209641f
C77 C6_P_btm C1_P_btm 0.127656f
C78 C7_P_btm C0_P_btm 0.140846f
C79 C4_P_btm C3_P_btm 9.61674f
C80 C5_P_btm C2_P_btm 0.13795f
C81 a_11453_44696# a_3090_45724# 0.232756f
C82 C8_P_btm C0_dummy_P_btm 0.234177f
C83 a_n2002_35608# VDD 0.522933f
C84 EN_VIN_BSTR_N C5_N_btm 0.115337f
C85 a_8696_44636# a_n2661_43922# 0.257466f
C86 a_10193_42453# a_3422_30871# 0.404849f
C87 a_4791_45118# a_2711_45572# 0.160646f
C88 a_3422_30871# VDD 1.12305f
C89 a_743_42282# a_564_42282# 0.169821f
C90 a_n2288_47178# VDD 0.29372f
C91 a_18479_45785# a_19319_43548# 0.102555f
C92 a_10903_43370# a_10809_44734# 0.353301f
C93 a_768_44030# a_2437_43646# 0.137571f
C94 a_17715_44484# a_15861_45028# 0.184272f
C95 a_584_46384# a_2063_45854# 0.406382f
C96 a_n4209_39590# a_n3420_39616# 0.234699f
C97 a_2324_44458# a_949_44458# 0.323116f
C98 a_8696_44636# a_17478_45572# 0.185985f
C99 a_22589_40599# a_22527_39145# 1.41544f
C100 a_n1613_43370# a_33_46660# 0.599895f
C101 a_n97_42460# a_n1853_43023# 0.151542f
C102 a_15095_43370# a_14955_43396# 0.130374f
C103 a_19963_31679# VDD 0.605523f
C104 a_3090_45724# a_9145_43396# 0.189557f
C105 a_3232_43370# a_1423_45028# 0.396815f
C106 a_11901_46660# a_12469_46902# 0.175891f
C107 a_10835_43094# a_10796_42968# 0.671797f
C108 a_7640_43914# VDD 0.196713f
C109 a_n2293_45010# a_895_43940# 0.283316f
C110 a_n971_45724# a_3065_45002# 0.220337f
C111 a_13259_45724# a_22400_42852# 0.34531f
C112 a_4185_45028# a_4958_30871# 0.121495f
C113 a_n2312_38680# VDD 0.540248f
C114 a_n913_45002# a_12281_43396# 0.28203f
C115 a_16414_43172# VDD 0.201389f
C116 a_9823_46155# VDD 0.102474f
C117 a_15493_43396# a_15493_43940# 0.188034f
C118 a_20205_31679# a_20447_31679# 9.01329f
C119 a_7174_31319# VDD 0.670432f
C120 a_4883_46098# a_n881_46662# 0.193691f
C121 a_12549_44172# a_4190_30871# 0.270972f
C122 VREF_GND VCM 2.79113f
C123 a_16137_43396# a_16414_43172# 0.179708f
C124 a_n1991_42858# a_n1641_43230# 0.229804f
C125 a_n2840_42826# a_n3674_39304# 0.16082f
C126 a_n2157_42858# a_n1076_43230# 0.102325f
C127 a_5111_44636# a_5891_43370# 0.702087f
C128 en_comp a_n2293_43922# 0.412872f
C129 a_1423_45028# a_8975_43940# 0.331942f
C130 a_13059_46348# a_3483_46348# 0.319214f
C131 a_765_45546# a_1176_45822# 0.241847f
C132 a_10729_43914# VDD 0.681371f
C133 a_19787_47423# VDD 0.256911f
C134 a_21487_43396# VDD 0.222231f
C135 a_n784_42308# a_7174_31319# 1.93626f
C136 a_20107_46660# VDD 0.442554f
C137 a_1138_42852# a_1307_43914# 0.123153f
C138 a_5937_45572# a_5205_44484# 0.481405f
C139 a_n2293_46634# a_14673_44172# 0.100552f
C140 a_4646_46812# a_7640_43914# 0.183308f
C141 a_3483_46348# a_13556_45296# 0.375978f
C142 a_5932_42308# VDD 0.534768f
C143 a_5934_30871# C5_N_btm 0.139996f
C144 a_n2129_43609# a_n2012_43396# 0.183186f
C145 a_n1177_43370# a_n1352_43396# 0.233657f
C146 a_20273_45572# a_20623_45572# 0.219856f
C147 a_16327_47482# a_15743_43084# 1.21037f
C148 a_n357_42282# a_18184_42460# 0.106442f
C149 C6_P_btm C2_P_btm 0.137206f
C150 C7_P_btm C1_P_btm 0.128479f
C151 C5_P_btm C3_P_btm 0.135528f
C152 a_12861_44030# a_16388_46812# 0.11634f
C153 C8_P_btm C0_P_btm 0.146541f
C154 a_13507_46334# a_15227_44166# 0.235687f
C155 C9_P_btm C0_dummy_P_btm 0.111645f
C156 EN_VIN_BSTR_N C4_N_btm 0.116925f
C157 a_1423_45028# VDD 4.06861f
C158 a_11967_42832# a_4958_30871# 0.239255f
C159 a_19692_46634# a_20411_46873# 0.215749f
C160 a_3080_42308# a_7174_31319# 0.22305f
C161 a_n2497_47436# VDD 1.33346f
C162 a_17583_46090# a_17715_44484# 0.22771f
C163 a_n1613_43370# a_n2661_45010# 0.223356f
C164 a_n784_42308# a_5932_42308# 0.151611f
C165 a_n755_45592# a_2713_42308# 0.243663f
C166 a_n1899_43946# a_n984_44318# 0.118759f
C167 a_n2661_45546# a_n443_42852# 0.141363f
C168 a_19692_46634# a_3422_30871# 0.208985f
C169 a_8696_44636# a_15861_45028# 0.26484f
C170 a_n1613_43370# a_171_46873# 0.11335f
C171 a_8128_46384# a_n1925_46634# 0.21095f
C172 a_5807_45002# a_13747_46662# 0.103485f
C173 a_14205_43396# a_14955_43396# 0.157423f
C174 a_22591_45572# VDD 0.314172f
C175 a_13159_45002# a_13348_45260# 0.105274f
C176 a_11735_46660# a_12251_46660# 0.105995f
C177 a_10518_42984# a_10796_42968# 0.118759f
C178 a_6109_44484# VDD 0.243629f
C179 a_3080_42308# a_5932_42308# 14.0282f
C180 a_n1177_44458# a_n1352_44484# 0.233657f
C181 a_n1151_42308# a_n913_45002# 0.395136f
C182 a_n971_45724# a_2680_45002# 0.108251f
C183 a_3232_43370# a_3457_43396# 0.131408f
C184 a_n2104_46634# VDD 0.286113f
C185 a_n2438_43548# a_n2661_43370# 0.147387f
C186 a_16327_47482# a_17970_44736# 0.219775f
C187 a_12891_46348# a_11691_44458# 0.141379f
C188 a_4646_46812# a_1423_45028# 0.415897f
C189 a_15567_42826# VDD 0.163583f
C190 a_n2956_38216# a_n3565_38216# 0.307285f
C191 a_9569_46155# VDD 0.19288f
C192 a_10193_42453# a_20712_42282# 0.157661f
C193 a_20365_43914# a_20623_43914# 0.22264f
C194 a_13259_45724# en_comp 0.19355f
C195 a_3754_39134# a_3754_38802# 0.296258f
C196 a_n4064_39616# C9_P_btm 0.215899f
C197 a_12861_44030# a_19321_45002# 0.10527f
C198 a_20712_42282# VDD 0.282526f
C199 a_11599_46634# a_5807_45002# 0.303048f
C200 a_7754_39964# a_7754_38470# 0.241119f
C201 a_n356_44636# a_1606_42308# 0.282657f
C202 a_3357_43084# a_3232_43370# 0.118744f
C203 a_12549_44172# a_765_45546# 0.118284f
C204 VREF VCM 44.262398f
C205 a_n1991_42858# a_n1423_42826# 0.186387f
C206 en_comp a_n2661_43922# 0.237031f
C207 a_7499_43078# a_11750_44172# 0.195997f
C208 a_15227_44166# a_17701_42308# 0.172697f
C209 a_765_45546# a_1208_46090# 0.134766f
C210 a_22959_42860# a_14097_32519# 0.166017f
C211 a_10405_44172# VDD 0.408512f
C212 a_19386_47436# VDD 0.121241f
C213 a_13059_46348# a_13249_42308# 0.306398f
C214 a_12861_44030# a_18184_42460# 0.266953f
C215 a_768_44030# a_1307_43914# 1.13357f
C216 a_20556_43646# VDD 0.34939f
C217 a_19551_46910# VDD 0.226848f
C218 a_5937_45572# a_6431_45366# 0.129839f
C219 a_13661_43548# a_11967_42832# 0.165876f
C220 a_3483_46348# a_9482_43914# 0.130172f
C221 a_6171_42473# VDD 0.184622f
C222 a_4791_45118# a_4883_46098# 0.135093f
C223 a_12861_44030# a_15811_47375# 0.144648f
C224 a_11967_42832# a_10835_43094# 0.263495f
C225 a_20107_45572# a_20623_45572# 0.103168f
C226 a_20273_45572# a_20841_45814# 0.175891f
C227 a_526_44458# a_n356_44636# 0.142971f
C228 C6_P_btm C3_P_btm 0.133742f
C229 C7_P_btm C2_P_btm 0.138288f
C230 C5_P_btm C4_P_btm 18.6196f
C231 a_12861_44030# a_13059_46348# 0.504219f
C232 C8_P_btm C1_P_btm 0.129306f
C233 C10_P_btm C0_dummy_P_btm 0.749362f
C234 EN_VIN_BSTR_N C3_N_btm 0.100325f
C235 C9_P_btm C0_P_btm 0.146135f
C236 a_18429_43548# a_16823_43084# 0.130506f
C237 a_19692_46634# a_20107_46660# 0.126737f
C238 a_20980_44850# VDD 0.132317f
C239 a_n2833_47464# VDD 0.461379f
C240 a_6969_46634# VDD 0.154507f
C241 a_n1331_43914# a_n1549_44318# 0.209641f
C242 a_n452_45724# a_n356_45724# 0.318161f
C243 a_n4064_40160# a_n4064_39616# 5.80519f
C244 a_n4209_39590# a_n3565_39590# 6.15218f
C245 a_2124_47436# a_584_46384# 0.220021f
C246 a_n1741_47186# a_4915_47217# 0.128899f
C247 a_n2302_37984# VDD 0.350854f
C248 a_n1613_43370# a_n133_46660# 0.347805f
C249 a_3726_37500# CAL_P 0.102027f
C250 a_3357_43084# VDD 1.66202f
C251 a_n4318_39304# a_n3674_39304# 2.9537f
C252 a_2437_43646# SINGLE_ENDED 0.117817f
C253 a_7499_43078# a_5891_43370# 1.00892f
C254 a_n2438_43548# a_n2157_46122# 0.270054f
C255 a_11813_46116# a_11901_46660# 0.211542f
C256 a_13507_46334# a_10809_44734# 0.603934f
C257 a_10518_42984# a_10835_43094# 0.102355f
C258 a_13747_46662# a_14495_45572# 0.288916f
C259 a_n1151_42308# a_n1059_45260# 0.16984f
C260 a_3483_46348# a_4419_46090# 0.218073f
C261 a_11599_46634# a_20107_45572# 0.246047f
C262 a_375_42282# a_n1557_42282# 0.450989f
C263 a_526_44458# a_3823_42558# 0.183187f
C264 a_n2293_46634# VDD 1.52629f
C265 a_10193_42453# a_5342_30871# 0.151919f
C266 a_16327_47482# a_17767_44458# 0.269619f
C267 a_9290_44172# a_7499_43078# 0.597117f
C268 a_5342_30871# VDD 0.496295f
C269 a_9625_46129# VDD 0.996485f
C270 a_20205_31679# a_19963_31679# 9.023429f
C271 VDAC_Pi a_3754_38470# 0.389564f
C272 a_10227_46804# a_12549_44172# 0.360691f
C273 a_20107_42308# VDD 0.284252f
C274 a_5937_45572# a_6453_43914# 0.144397f
C275 a_n1741_47186# a_10809_44734# 0.332771f
C276 VIN_N VCM 1.7189f
C277 a_11453_44696# a_12741_44636# 1.02327f
C278 VREF VREF_GND 44.051197f
C279 a_16237_45028# VDD 0.248452f
C280 a_n2157_42858# a_n1641_43230# 0.110532f
C281 a_16922_45042# a_18494_42460# 0.242236f
C282 a_18315_45260# a_18587_45118# 0.13675f
C283 a_7499_43078# a_10807_43548# 0.119721f
C284 a_9672_43914# VDD 0.150499f
C285 a_10193_42453# a_743_42282# 1.1645f
C286 a_18597_46090# VDD 0.930122f
C287 a_18479_47436# START 0.313639f
C288 a_3357_43084# a_3080_42308# 0.233522f
C289 a_12861_44030# a_19778_44110# 0.113118f
C290 a_12549_44172# a_1307_43914# 1.82879f
C291 a_743_42282# VDD 0.597869f
C292 a_19123_46287# VDD 0.336379f
C293 a_5937_45572# a_6171_45002# 0.206948f
C294 a_12549_44172# a_18579_44172# 0.154956f
C295 a_n1741_47186# a_n881_46662# 0.179671f
C296 a_5755_42308# VDD 0.229304f
C297 a_n3420_38528# a_n4064_38528# 8.203589f
C298 a_2277_45546# VDD 0.209584f
C299 C6_P_btm C4_P_btm 0.143514f
C300 C7_P_btm C3_P_btm 0.134911f
C301 a_n2293_46634# a_4646_46812# 0.135642f
C302 C8_P_btm C2_P_btm 0.138777f
C303 EN_VIN_BSTR_N C2_N_btm 0.118072f
C304 C9_P_btm C1_P_btm 0.132506f
C305 C10_P_btm C0_P_btm 0.365593f
C306 a_5807_45002# a_5257_43370# 0.683815f
C307 a_626_44172# VDD 0.621601f
C308 a_16137_43396# a_743_42282# 0.183525f
C309 a_19692_46634# a_20556_43646# 0.118928f
C310 a_413_45260# a_n2661_44458# 0.69469f
C311 a_n2312_38680# a_n2956_38680# 6.25577f
C312 a_11453_44696# a_16375_45002# 0.104273f
C313 a_11691_44458# a_14673_44172# 0.371587f
C314 a_6755_46942# VDD 1.05713f
C315 a_n1899_43946# a_n1549_44318# 0.218775f
C316 a_n2065_43946# a_n984_44318# 0.102325f
C317 a_n755_45592# a_997_45618# 0.133124f
C318 a_n237_47217# a_n1151_42308# 0.63407f
C319 a_n4209_39590# a_n4334_39616# 0.25243f
C320 a_8049_45260# VDD 1.89366f
C321 a_n2293_46634# a_14021_43940# 0.202404f
C322 a_n4064_37984# VDD 1.70621f
C323 a_22589_40599# a_22537_40625# 1.96968f
C324 a_n881_46662# a_n743_46660# 0.527182f
C325 a_n1613_43370# a_n2438_43548# 1.04064f
C326 a_2437_43646# START 0.12936f
C327 a_19479_31679# VDD 0.579933f
C328 a_13017_45260# a_13159_45002# 0.160415f
C329 a_n2438_43548# a_n2293_46098# 0.409291f
C330 a_11735_46660# a_11901_46660# 0.579036f
C331 a_13661_43548# a_3483_46348# 0.381471f
C332 a_3539_42460# a_3318_42354# 0.161793f
C333 a_n2293_45010# a_453_43940# 0.181603f
C334 a_413_45260# a_19237_31679# 0.119197f
C335 a_13259_45724# a_13667_43396# 0.160676f
C336 a_13747_46662# a_13249_42308# 0.134714f
C337 a_3483_46348# a_4185_45028# 0.430982f
C338 a_15037_43940# VDD 0.190221f
C339 a_8975_43940# a_9028_43914# 0.184602f
C340 a_10057_43914# a_9672_43914# 0.143523f
C341 a_11823_42460# a_12089_42308# 0.335983f
C342 a_n2442_46660# VDD 0.693209f
C343 a_n2293_43922# a_n2472_43914# 0.189122f
C344 a_526_44458# a_3316_45546# 0.128261f
C345 a_768_44030# a_11827_44484# 0.831344f
C346 a_5937_45572# a_8746_45002# 0.121678f
C347 a_19321_45002# a_16922_45042# 0.493823f
C348 a_15279_43071# VDD 0.189193f
C349 a_17124_42282# a_17303_42282# 0.172579f
C350 a_n3674_37592# a_n3420_37984# 0.172946f
C351 a_n2956_38216# a_n4209_38216# 0.232905f
C352 a_8953_45546# VDD 1.32809f
C353 a_20269_44172# a_20365_43914# 0.419086f
C354 a_3090_45724# a_9313_44734# 2.43867f
C355 a_9290_44172# a_n2661_43370# 0.185465f
C356 a_11525_45546# a_11682_45822# 0.18824f
C357 a_n443_46116# a_n743_46660# 0.532861f
C358 a_7754_39300# a_7754_38968# 0.296258f
C359 a_12861_44030# a_13747_46662# 0.139424f
C360 a_13258_32519# VDD 3.19378f
C361 a_7754_40130# a_7754_38470# 0.112286f
C362 a_5937_45572# a_5663_43940# 0.177912f
C363 a_10193_42453# a_20193_45348# 0.305022f
C364 a_n863_45724# a_n356_44636# 0.301674f
C365 VIN_N VREF_GND 16.4969f
C366 VIN_P VCM 1.7189f
C367 a_3877_44458# a_6969_46634# 0.101189f
C368 a_4646_46812# a_6755_46942# 0.362783f
C369 a_20193_45348# VDD 0.793111f
C370 a_n1853_43023# a_n1991_42858# 0.237526f
C371 a_7499_43078# a_10949_43914# 0.152939f
C372 a_22223_42860# a_22400_42852# 0.154104f
C373 a_9028_43914# VDD 0.17194f
C374 a_18989_43940# a_19006_44850# 0.168452f
C375 a_18780_47178# VDD 0.245515f
C376 a_12861_44030# a_18911_45144# 0.169f
C377 a_9803_42558# a_9885_42558# 0.171361f
C378 a_n784_42308# a_13258_32519# 0.140549f
C379 a_20301_43646# VDD 0.296691f
C380 a_18184_42460# a_15743_43084# 0.182123f
C381 a_18285_46348# VDD 0.259614f
C382 a_5937_45572# a_3232_43370# 0.662525f
C383 a_8199_44636# a_6171_45002# 0.163434f
C384 a_12861_44030# a_11599_46634# 0.169929f
C385 a_6123_31319# C4_N_btm 0.132906f
C386 a_n3420_38528# a_n2946_38778# 0.236674f
C387 a_1609_45822# VDD 0.270106f
C388 a_n2129_43609# a_n447_43370# 0.119518f
C389 a_n2267_43396# a_n1352_43396# 0.124988f
C390 a_20107_45572# a_20273_45572# 0.667378f
C391 a_3483_46348# a_11967_42832# 0.264293f
C392 C6_P_btm C5_P_btm 22.305399f
C393 C7_P_btm C4_P_btm 0.145303f
C394 C8_P_btm C3_P_btm 0.134581f
C395 EN_VIN_BSTR_N C1_N_btm 0.110046f
C396 a_1983_46706# a_n2661_46098# 0.147223f
C397 C9_P_btm C2_P_btm 0.141891f
C398 C10_P_btm C1_P_btm 0.31753f
C399 a_19692_46634# a_743_42282# 0.150479f
C400 a_3232_43370# a_11691_44458# 0.251483f
C401 a_n2312_38680# a_n2956_39304# 5.96956f
C402 a_n2312_38680# a_n3565_39304# 0.418567f
C403 a_5883_43914# a_5891_43370# 0.216958f
C404 a_9290_44172# a_10809_44734# 0.239594f
C405 SMPL_ON_N a_413_45260# 0.199669f
C406 a_3090_45724# a_2711_45572# 0.555348f
C407 a_10249_46116# VDD 1.03004f
C408 a_n1899_43946# a_n1331_43914# 0.171939f
C409 a_n746_45260# a_n1151_42308# 0.116939f
C410 a_n2109_47186# a_4915_47217# 0.352259f
C411 a_22959_43948# a_17538_32519# 0.168682f
C412 a_16855_45546# a_8696_44636# 0.112262f
C413 a_n2946_37984# VDD 0.38275f
C414 a_n881_46662# a_n1021_46688# 0.15991f
C415 a_n1613_43370# a_n743_46660# 0.521102f
C416 a_14358_43442# a_14205_43396# 0.163543f
C417 a_9803_43646# a_10341_43396# 0.11445f
C418 a_14579_43548# a_15095_43370# 0.109081f
C419 a_22223_45572# VDD 0.287831f
C420 a_n357_42282# a_11967_42832# 0.153035f
C421 a_6171_45002# a_16751_45260# 0.104212f
C422 a_n2017_45002# a_n2293_42834# 0.28698f
C423 a_13507_46334# a_6945_45028# 0.187229f
C424 a_n743_46660# a_n2293_46098# 0.213418f
C425 a_11735_46660# a_11813_46116# 0.162547f
C426 a_10083_42826# a_10518_42984# 0.234322f
C427 a_n2267_44484# a_n1352_44484# 0.118759f
C428 a_413_45260# a_22959_44484# 0.202222f
C429 a_n2312_39304# a_n3565_39590# 0.491833f
C430 a_n746_45260# a_327_44734# 0.256943f
C431 a_13661_43548# a_13249_42308# 0.486588f
C432 a_13565_43940# VDD 0.175245f
C433 a_10193_42453# a_5534_30871# 0.136243f
C434 a_n2472_46634# VDD 0.287589f
C435 a_20193_45348# a_14021_43940# 0.118757f
C436 a_12549_44172# a_11827_44484# 1.40268f
C437 a_8199_44636# a_8746_45002# 0.680077f
C438 a_5534_30871# VDD 0.513761f
C439 a_17124_42282# a_4958_30871# 0.20224f
C440 en_comp a_22400_42852# 0.721871f
C441 a_5937_45572# VDD 2.20055f
C442 a_n2810_45572# a_n3565_38216# 0.104999f
C443 VDAC_Pi VDAC_Ni 3.18068f
C444 a_12861_44030# a_13661_43548# 0.8566f
C445 a_n3565_39590# C8_P_btm 0.384801f
C446 a_19647_42308# VDD 0.227331f
C447 a_3357_43084# a_5111_44636# 0.318002f
C448 a_n745_45366# a_n467_45028# 0.110406f
C449 a_n1741_47186# a_6945_45028# 2.51584f
C450 VIN_N VREF 0.775904f
C451 a_3877_44458# a_6755_46942# 0.388535f
C452 VIN_P VREF_GND 16.4969f
C453 a_11691_44458# VDD 3.25709f
C454 a_n2157_42858# a_n1991_42858# 0.905962f
C455 a_10227_46804# a_15890_42674# 0.159412f
C456 a_3537_45260# a_5891_43370# 0.359819f
C457 a_14537_43396# a_14539_43914# 0.135541f
C458 a_7499_43078# a_10729_43914# 0.23002f
C459 a_8333_44056# VDD 0.124235f
C460 a_5534_30871# a_n784_42308# 9.92256f
C461 a_18479_47436# VDD 1.47669f
C462 a_n913_45002# a_n97_42460# 0.109647f
C463 a_10193_42453# a_4190_30871# 0.305842f
C464 a_n971_45724# a_n699_43396# 0.139047f
C465 a_n2293_46634# a_5111_44636# 0.130609f
C466 a_4190_30871# VDD 1.36846f
C467 a_n356_44636# a_2982_43646# 0.434193f
C468 a_1307_43914# a_3935_42891# 0.318189f
C469 a_17829_46910# VDD 0.37446f
C470 a_8199_44636# a_3232_43370# 0.32342f
C471 a_3483_46348# a_13017_45260# 0.51131f
C472 a_n3565_38502# a_n4064_38528# 0.228245f
C473 a_n443_42852# VDD 3.69394f
C474 a_n1699_43638# a_n1917_43396# 0.209641f
C475 a_16327_47482# a_17324_43396# 0.216094f
C476 a_4791_45118# a_4361_42308# 0.111224f
C477 C7_P_btm C5_P_btm 0.151416f
C478 VDAC_P VCM 11.743501f
C479 C8_P_btm C4_P_btm 0.145646f
C480 EN_VIN_BSTR_N C0_N_btm 0.12803f
C481 C9_P_btm C3_P_btm 0.137552f
C482 C10_P_btm C2_P_btm 0.327137f
C483 a_13507_46334# a_15559_46634# 0.216791f
C484 a_16137_43396# a_4190_30871# 0.113768f
C485 a_375_42282# VDD 0.591443f
C486 a_n913_45002# a_742_44458# 0.302053f
C487 a_19692_46634# a_20301_43646# 0.110092f
C488 a_4646_46812# a_5937_45572# 0.105447f
C489 a_2063_45854# a_6472_45840# 0.545607f
C490 a_n4318_39304# a_n3420_39616# 0.256393f
C491 a_22165_42308# a_22223_42860# 0.171681f
C492 a_2324_44458# a_15682_46116# 0.343876f
C493 a_6655_43762# VDD 0.132357f
C494 a_10554_47026# VDD 0.205847f
C495 a_n2065_43946# a_n1549_44318# 0.110816f
C496 a_12861_44030# a_11967_42832# 0.209245f
C497 a_n357_42282# a_n755_45592# 0.664842f
C498 a_14635_42282# VDD 0.369964f
C499 a_n971_45724# a_n1151_42308# 0.682801f
C500 a_1209_47178# a_584_46384# 0.104123f
C501 a_n913_45002# a_10533_42308# 0.246621f
C502 a_n2661_42834# a_n2840_42826# 0.174935f
C503 a_16855_45546# a_16680_45572# 0.233657f
C504 a_15903_45785# a_16020_45572# 0.157972f
C505 a_n3420_37984# VDD 0.930532f
C506 a_n881_46662# a_n1925_46634# 0.467945f
C507 a_6151_47436# a_6755_46942# 0.361724f
C508 a_9803_43646# a_9885_43646# 0.171361f
C509 a_3422_30871# COMP_P 0.208163f
C510 a_2437_43646# VDD 1.17411f
C511 a_n1699_44726# a_n1917_44484# 0.209641f
C512 a_3357_43084# a_3905_42865# 0.125186f
C513 a_5807_45002# a_13249_42308# 0.725941f
C514 a_n1925_46634# a_8162_45546# 0.104508f
C515 a_n2661_46634# a_10193_42453# 0.351509f
C516 a_18479_45785# a_4190_30871# 0.123942f
C517 a_n2661_43922# a_n2840_43914# 0.171265f
C518 a_n2661_46634# VDD 2.23057f
C519 a_8199_44636# a_10193_42453# 0.236934f
C520 a_8049_45260# a_20205_31679# 0.301209f
C521 a_14543_43071# VDD 0.18866f
C522 a_8199_44636# VDD 1.43837f
C523 a_10193_42453# a_19511_42282# 0.133376f
C524 a_13259_45724# a_n913_45002# 0.142601f
C525 a_19511_42282# VDD 0.244902f
C526 a_12861_44030# a_5807_45002# 0.214011f
C527 a_7754_40130# a_3754_38470# 0.191861f
C528 a_7754_39964# VDAC_Ni 0.207118f
C529 a_5343_44458# a_7963_42308# 0.108654f
C530 a_13661_43548# a_19268_43646# 0.136251f
C531 VIN_P VREF 0.775904f
C532 a_11453_44696# a_11415_45002# 0.123733f
C533 a_n2157_42858# a_n1853_43023# 0.290902f
C534 a_10227_46804# a_15959_42545# 0.152289f
C535 a_1423_45028# a_9838_44484# 0.254741f
C536 a_3537_45260# a_8375_44464# 0.10437f
C537 a_7499_43078# a_10405_44172# 0.132405f
C538 a_10227_46804# a_8746_45002# 0.117547f
C539 a_1823_45246# a_3823_42558# 0.137565f
C540 a_18287_44626# a_11967_42832# 0.789765f
C541 a_18143_47464# VDD 0.388551f
C542 a_n1059_45260# a_n97_42460# 0.869353f
C543 a_1823_45246# a_3503_45724# 0.295715f
C544 a_21259_43561# VDD 0.192954f
C545 a_765_45546# VDD 2.19953f
C546 a_1307_43914# a_3681_42891# 0.236785f
C547 a_6667_45809# a_6598_45938# 0.209641f
C548 a_6511_45714# a_7227_45028# 0.213161f
C549 a_8953_45546# a_5111_44636# 0.181796f
C550 a_1606_42308# VCM 0.152876f
C551 a_1273_38525# a_2113_38308# 0.325472f
C552 a_4921_42308# VDD 0.214995f
C553 a_n4209_38502# a_n2302_38778# 0.406492f
C554 a_n3565_38502# a_n2946_38778# 0.406164f
C555 a_n3690_38528# a_n3420_38528# 0.431104f
C556 a_n4334_38528# a_n4064_38528# 0.449049f
C557 a_n2433_43396# a_n1352_43396# 0.102325f
C558 a_509_45822# VDD 0.190119f
C559 a_n2267_43396# a_n1917_43396# 0.227165f
C560 a_16327_47482# a_17499_43370# 0.34052f
C561 C7_P_btm C6_P_btm 26.0771f
C562 CAL_P RST_Z 0.551895f
C563 VDAC_P VREF_GND 0.203715f
C564 C8_P_btm C5_P_btm 0.145019f
C565 a_22629_38406# VDD 0.315181f
C566 C9_P_btm C4_P_btm 0.154834f
C567 C10_P_btm C3_P_btm 0.321945f
C568 a_16751_45260# VDD 0.121848f
C569 a_413_45260# a_19721_31679# 0.116395f
C570 a_19333_46634# a_19123_46287# 0.113955f
C571 a_11453_44696# a_13259_45724# 0.251534f
C572 a_n2661_44458# a_n2661_43922# 6.64988f
C573 a_18287_44626# a_18989_43940# 0.193279f
C574 a_18443_44721# a_18374_44850# 0.209641f
C575 a_1307_43914# a_5663_43940# 0.11718f
C576 a_4185_45028# a_n1925_42282# 0.638728f
C577 a_5534_30871# a_n3420_39072# 0.339008f
C578 a_10623_46897# VDD 0.189083f
C579 a_n1761_44111# a_n1899_43946# 0.737653f
C580 a_20202_43084# a_n913_45002# 0.322116f
C581 a_13291_42460# VDD 0.546706f
C582 a_1239_47204# a_1431_47204# 0.219138f
C583 a_n2109_47186# a_4791_45118# 0.34446f
C584 a_375_42282# a_196_42282# 0.165785f
C585 a_1138_42852# a_n356_44636# 0.29814f
C586 a_8199_44636# a_10057_43914# 0.113262f
C587 a_n3690_38304# VDD 0.363068f
C588 a_n1613_43370# a_n1925_46634# 0.33524f
C589 a_14579_43548# a_14358_43442# 0.142377f
C590 a_21513_45002# VDD 0.416919f
C591 a_3232_43370# a_1307_43914# 0.14252f
C592 a_3090_45724# a_8685_43396# 2.11639f
C593 a_11453_44696# a_18189_46348# 0.534507f
C594 a_n2267_44484# a_n1917_44484# 0.212549f
C595 a_13259_45724# a_9145_43396# 0.155949f
C596 a_n2433_44484# a_n1352_44484# 0.102355f
C597 a_n971_45724# a_413_45260# 0.937818f
C598 a_n2293_46634# a_7499_43078# 0.14773f
C599 a_3147_46376# a_3483_46348# 0.207919f
C600 a_5342_30871# a_14113_42308# 0.203397f
C601 a_4190_30871# a_n3420_39072# 0.10848f
C602 a_n2956_39768# VDD 0.697168f
C603 a_3483_46348# a_13249_42308# 0.338396f
C604 a_8199_44636# a_10180_45724# 0.216999f
C605 a_19692_46634# a_2437_43646# 0.293918f
C606 a_13460_43230# VDD 0.276534f
C607 a_8349_46414# VDD 0.209819f
C608 a_n2810_45572# a_n4209_38216# 0.195791f
C609 a_13259_45724# a_n1059_45260# 0.390886f
C610 a_2063_45854# a_2107_46812# 0.214026f
C611 a_n3420_37984# a_n4064_37440# 7.43287f
C612 a_n1059_45260# a_n467_45028# 0.229142f
C613 a_12465_44636# a_12741_44636# 0.914049f
C614 a_22959_45036# VDD 0.30999f
C615 a_2711_45572# a_15493_43940# 0.128282f
C616 a_n2017_45002# a_n2293_43922# 0.654835f
C617 a_10227_46804# a_15803_42450# 0.296174f
C618 a_18248_44752# a_11967_42832# 0.500539f
C619 a_10227_46804# VDD 2.77567f
C620 a_n2017_45002# a_n97_42460# 0.169401f
C621 a_13059_46348# a_11823_42460# 0.256727f
C622 a_4190_30871# C10_N_btm 0.446355f
C623 a_17339_46660# VDD 0.555596f
C624 a_6472_45840# a_7227_45028# 0.208286f
C625 a_13259_45724# a_15599_45572# 0.205417f
C626 a_5742_30871# EN_VIN_BSTR_N 0.643089f
C627 a_1666_39043# a_2684_37794# 0.193789f
C628 a_n3565_38502# a_n3420_38528# 0.278952f
C629 a_n4209_38502# a_n4064_38528# 0.265711f
C630 a_12861_44030# a_13487_47204# 0.127147f
C631 a_n2267_43396# a_n1699_43638# 0.179796f
C632 a_16327_47482# a_16759_43396# 0.152273f
C633 CAL_P VDD 22.4816f
C634 VDAC_N VCM 11.7445f
C635 C8_P_btm C6_P_btm 0.163943f
C636 C10_P_btm C4_P_btm 0.703336f
C637 C9_P_btm C5_P_btm 0.150576f
C638 a_18597_46090# a_15227_44166# 0.150202f
C639 a_1307_43914# VDD 3.92807f
C640 a_10193_42453# a_18579_44172# 0.12582f
C641 a_14180_46812# a_14513_46634# 0.253235f
C642 a_18579_44172# VDD 0.38178f
C643 a_5111_44636# a_8333_44056# 0.280148f
C644 a_18248_44752# a_18989_43940# 0.207562f
C645 a_11827_44484# a_14673_44172# 0.150125f
C646 a_8103_44636# a_8375_44464# 0.13675f
C647 a_4185_45028# a_526_44458# 0.162857f
C648 a_12465_44636# a_413_45260# 0.28925f
C649 a_9396_43370# VDD 0.288403f
C650 a_10467_46802# VDD 0.401016f
C651 a_n755_45592# a_1755_42282# 1.52791f
C652 a_n2065_43946# a_n1899_43946# 0.614122f
C653 a_n746_45260# a_175_44278# 0.159759f
C654 a_n1099_45572# a_n755_45592# 0.193775f
C655 a_310_45028# a_n357_42282# 0.113929f
C656 a_13003_42852# VDD 0.132655f
C657 a_n971_45724# a_2905_45572# 0.118495f
C658 a_11967_42832# a_15743_43084# 0.180938f
C659 a_8034_45724# VDD 0.812726f
C660 a_15903_45785# a_15861_45028# 0.232345f
C661 a_n443_42852# a_5111_44636# 0.584506f
C662 a_n3565_38216# VDD 0.901085f
C663 a_11787_45002# a_11963_45334# 0.185422f
C664 a_6755_46942# a_15227_44166# 0.288173f
C665 a_n2267_44484# a_n1699_44726# 0.172319f
C666 a_20202_43084# a_19987_42826# 0.177726f
C667 a_3357_43084# a_2998_44172# 0.119142f
C668 a_16327_47482# a_19256_45572# 0.235006f
C669 a_n1151_42308# a_n2661_45010# 0.155007f
C670 a_n2840_46634# VDD 0.306342f
C671 a_3483_46348# a_13904_45546# 0.125708f
C672 a_n2293_46634# a_n2661_43370# 2.59564f
C673 a_8016_46348# a_10193_42453# 0.125497f
C674 a_5937_45572# a_9049_44484# 0.311862f
C675 a_8953_45546# a_7499_43078# 0.108436f
C676 a_13635_43156# VDD 0.463701f
C677 a_3483_46348# CLK 0.408122f
C678 a_8016_46348# VDD 1.42798f
C679 a_10490_45724# a_10907_45822# 0.229517f
C680 a_n971_45724# a_104_43370# 0.156156f
C681 a_n4209_39590# C9_P_btm 0.786375f
C682 a_16327_47482# a_12549_44172# 0.123271f
C683 a_6151_47436# a_n2661_46634# 0.140541f
C684 a_n237_47217# a_1799_45572# 0.417887f
C685 a_11682_45822# VDD 0.316586f
C686 a_22223_45036# VDD 0.300162f
C687 a_17591_47464# VDD 0.421992f
C688 a_167_45260# a_1848_45724# 0.359783f
C689 a_5934_30871# a_5742_30871# 16.7261f
C690 a_6453_43914# a_n2661_42282# 0.122766f
C691 a_6472_45840# a_6598_45938# 0.178024f
C692 a_6511_45714# a_6667_45809# 0.113977f
C693 a_n2497_47436# a_n1613_43370# 0.402561f
C694 a_3905_42558# VDD 0.176395f
C695 a_n1151_42308# a_4883_46098# 0.407909f
C696 a_n3565_38502# a_n3690_38528# 0.246863f
C697 a_n2433_43396# a_n1917_43396# 0.108815f
C698 a_16327_47482# a_16977_43638# 0.15941f
C699 VDAC_N VREF_GND 0.203821f
C700 a_10227_46804# a_19692_46634# 0.239326f
C701 a_6151_47436# a_765_45546# 0.191559f
C702 a_12861_44030# a_14180_46812# 0.238709f
C703 C9_P_btm C6_P_btm 0.165353f
C704 C10_P_btm C5_P_btm 0.51798f
C705 C8_P_btm C7_P_btm 31.072699f
C706 a_n2661_42282# a_n3674_37592# 0.12829f
C707 a_16019_45002# VDD 0.174085f
C708 a_10341_43396# a_22591_43396# 0.172197f
C709 a_4791_45118# a_5932_42308# 0.212275f
C710 a_2982_43646# a_17303_42282# 0.139588f
C711 a_8103_44636# a_7640_43914# 0.101633f
C712 a_18287_44626# a_18443_44721# 0.10279f
C713 a_18248_44752# a_18374_44850# 0.170059f
C714 a_1307_43914# a_5013_44260# 0.358053f
C715 a_3483_46348# a_n1925_42282# 0.536704f
C716 a_4791_45118# a_1423_45028# 0.721318f
C717 a_8791_43396# VDD 0.191045f
C718 a_10428_46928# VDD 0.278873f
C719 a_n755_45592# a_1606_42308# 0.104938f
C720 a_n2065_43946# a_n1761_44111# 0.617556f
C721 a_1209_47178# a_1239_47204# 0.264529f
C722 a_n237_47217# a_2063_45854# 0.947844f
C723 a_22223_43948# a_14401_32519# 0.157135f
C724 a_15765_45572# a_16680_45572# 0.118759f
C725 a_n4334_38304# VDD 0.385989f
C726 a_4915_47217# a_6755_46942# 0.260675f
C727 a_9145_43396# a_15095_43370# 0.213415f
C728 a_8696_44636# a_n2661_44458# 1.37553f
C729 a_8128_46384# a_8349_46414# 0.101217f
C730 a_9127_43156# a_8952_43230# 0.234322f
C731 a_n2433_44484# a_n1917_44484# 0.113784f
C732 a_16327_47482# a_19431_45546# 0.344862f
C733 a_13747_46662# a_11823_42460# 0.521845f
C734 a_1823_45246# a_4704_46090# 0.164557f
C735 a_11453_44696# a_8696_44636# 2.67247f
C736 a_n1059_45260# a_15095_43370# 0.108103f
C737 a_9290_44172# a_13070_42354# 0.140007f
C738 a_22612_30879# VDD 3.23778f
C739 a_8953_45546# a_8568_45546# 0.136365f
C740 a_12549_44172# a_20567_45036# 0.176249f
C741 a_8016_46348# a_10180_45724# 0.259851f
C742 a_12895_43230# VDD 0.212352f
C743 a_9313_44734# a_10341_43396# 0.175125f
C744 a_7920_46348# VDD 0.100184f
C745 a_14955_43940# a_15493_43940# 0.110232f
C746 a_13904_45546# a_13249_42308# 0.13587f
C747 a_n971_45724# a_n97_42460# 0.581616f
C748 a_15811_47375# a_15928_47570# 0.161235f
C749 a_n3420_37984# a_n3420_37440# 0.132162f
C750 a_10193_42453# a_11827_44484# 0.121679f
C751 a_n2810_45028# a_n2956_37592# 6.13705f
C752 a_n913_45002# a_n967_45348# 1.00127f
C753 a_n1151_42308# a_11387_46155# 0.195225f
C754 a_11827_44484# VDD 0.615802f
C755 a_2711_45572# a_11341_43940# 1.54309f
C756 a_16922_45042# a_17719_45144# 0.22253f
C757 a_10227_46804# a_15486_42560# 0.227612f
C758 a_16588_47582# VDD 0.282243f
C759 a_n443_42852# a_685_42968# 0.104532f
C760 a_n2293_46634# a_3537_45260# 0.155982f
C761 a_1307_43914# a_1847_42826# 0.428505f
C762 a_9313_44734# a_n97_42460# 1.76217f
C763 a_6472_45840# a_6667_45809# 0.215953f
C764 a_n443_42852# a_7499_43078# 0.375366f
C765 a_15227_44166# a_11691_44458# 0.443265f
C766 a_1666_39587# a_2113_38308# 0.100592f
C767 a_n1435_47204# a_13487_47204# 0.135076f
C768 a_13717_47436# a_12861_44030# 0.319645f
C769 a_n4209_38502# a_n3420_38528# 0.230544f
C770 a_n2129_43609# a_n2267_43396# 0.230013f
C771 VDAC_P VIN_P 0.255243f
C772 a_12861_44030# a_14035_46660# 0.153051f
C773 C9_P_btm C7_P_btm 0.22201f
C774 C10_P_btm C6_P_btm 0.895671f
C775 a_18479_47436# a_15227_44166# 0.199537f
C776 a_15595_45028# VDD 0.156299f
C777 a_18834_46812# a_18285_46348# 0.144972f
C778 a_13885_46660# a_14513_46634# 0.101344f
C779 a_21195_42852# a_21671_42860# 0.177876f
C780 a_2982_43646# a_4958_30871# 0.136637f
C781 a_n443_42852# a_15781_43660# 0.22553f
C782 a_5343_44458# a_5891_43370# 1.06553f
C783 a_18248_44752# a_18443_44721# 0.206455f
C784 a_n1613_43370# a_3357_43084# 0.228593f
C785 a_3483_46348# a_526_44458# 0.134907f
C786 a_15015_46420# a_14840_46494# 0.233657f
C787 a_1606_42308# a_2351_42308# 0.191324f
C788 a_8147_43396# VDD 0.393534f
C789 a_10150_46912# VDD 0.284144f
C790 a_n1099_45572# a_310_45028# 0.333219f
C791 a_n2293_46098# a_3357_43084# 0.16657f
C792 a_n237_47217# a_584_46384# 0.645142f
C793 a_n971_45724# a_2553_47502# 0.23907f
C794 a_n443_46116# a_2813_43396# 0.124521f
C795 a_8953_45546# a_5883_43914# 0.262126f
C796 a_16333_45814# a_16115_45572# 0.209641f
C797 a_n4209_38216# VDD 0.834113f
C798 a_n1613_43370# a_n2293_46634# 0.103089f
C799 VDAC_P a_11206_38545# 0.101449f
C800 a_9145_43396# a_14205_43396# 0.13322f
C801 a_5111_44636# a_1307_43914# 0.114933f
C802 a_n2129_44697# a_n2267_44484# 0.698671f
C803 a_2711_45572# a_n97_42460# 0.137121f
C804 a_16327_47482# a_18691_45572# 0.162157f
C805 a_13661_43548# a_11823_42460# 0.116839f
C806 a_1823_45246# a_4419_46090# 0.340207f
C807 a_4791_45118# a_3357_43084# 0.144996f
C808 a_17517_44484# a_20640_44752# 0.54753f
C809 a_5111_44636# a_9396_43370# 0.203348f
C810 a_21588_30879# VDD 1.7842f
C811 a_8199_44636# a_7499_43078# 0.859274f
C812 a_15227_44166# a_2437_43646# 0.167451f
C813 a_12549_44172# a_18494_42460# 0.331306f
C814 a_526_44458# a_n357_42282# 0.220537f
C815 a_13113_42826# VDD 0.217254f
C816 a_15493_43396# a_19478_44306# 0.154347f
C817 a_3090_45724# a_5891_43370# 0.166094f
C818 a_5937_45572# a_n2661_43370# 0.202031f
C819 a_n971_45724# a_n447_43370# 0.113797f
C820 a_18214_42558# VDD 0.295211f
C821 a_584_46384# a_1123_46634# 0.370049f
C822 a_3754_39466# a_3754_39134# 0.296258f
C823 a_14401_32519# a_10341_43396# 0.133035f
C824 a_10907_45822# VDD 0.352181f
C825 a_16147_45260# a_1307_43914# 0.150161f
C826 a_12465_44636# a_11415_45002# 0.375509f
C827 a_n1151_42308# a_11133_46155# 0.162011f
C828 a_21359_45002# VDD 0.319372f
C829 a_13556_45296# a_15004_44636# 0.127354f
C830 a_1423_45028# a_6298_44484# 0.103777f
C831 a_16922_45042# a_17613_45144# 0.10967f
C832 a_10227_46804# a_15051_42282# 0.361922f
C833 a_3090_45724# a_9290_44172# 0.196232f
C834 a_12861_44030# a_13527_45546# 0.274077f
C835 a_n2661_42282# VDD 0.406474f
C836 a_16763_47508# VDD 0.392885f
C837 a_768_44030# a_13556_45296# 0.267809f
C838 a_167_45260# a_n755_45592# 1.02724f
C839 a_12861_44030# a_16922_45042# 0.120012f
C840 a_11415_45002# a_2711_45572# 0.337384f
C841 a_6123_31319# a_5742_30871# 0.106954f
C842 a_16823_43084# VDD 0.159922f
C843 a_3483_46348# a_8953_45002# 0.121322f
C844 a_6472_45840# a_6511_45714# 0.781352f
C845 a_19321_45002# a_17517_44484# 0.264473f
C846 a_5742_30871# EN_VIN_BSTR_P 0.645741f
C847 a_5932_42308# C3_N_btm 0.121156f
C848 a_13381_47204# a_13487_47204# 0.152045f
C849 a_n2433_43396# a_n2267_43396# 0.756435f
C850 C9_P_btm C8_P_btm 39.4538f
C851 a_22537_39537# VDD 0.313136f
C852 C10_P_btm C7_P_btm 1.39624f
C853 VDAC_N VIN_N 0.256435f
C854 a_15415_45028# VDD 0.191729f
C855 a_6293_42852# a_5755_42852# 0.114235f
C856 a_11823_42460# a_11967_42832# 0.573139f
C857 a_4185_45028# a_2982_43646# 0.243496f
C858 a_13885_46660# a_14180_46812# 0.150851f
C859 a_17609_46634# a_18285_46348# 0.115413f
C860 a_14209_32519# a_14097_32519# 10.7606f
C861 a_19279_43940# VDD 0.302681f
C862 a_18248_44752# a_18287_44626# 0.633819f
C863 a_1307_43914# a_3905_42865# 0.224019f
C864 a_3147_46376# a_526_44458# 0.352f
C865 a_7112_43396# VDD 0.273193f
C866 a_9863_46634# VDD 0.411318f
C867 a_13661_43548# a_14539_43914# 0.193767f
C868 a_12465_44636# a_n2661_43922# 0.17969f
C869 a_n863_45724# a_n755_45592# 1.76733f
C870 a_13259_45724# a_2711_45572# 1.26722f
C871 a_n4315_30879# a_n4209_39590# 4.31257f
C872 a_11136_42852# VDD 0.132515f
C873 a_n1741_47186# a_n1151_42308# 2.98024f
C874 a_n2109_47186# a_3785_47178# 0.190973f
C875 a_n746_45260# a_584_46384# 0.491308f
C876 a_n971_45724# a_2063_45854# 0.164981f
C877 a_20512_43084# a_10341_43396# 0.758407f
C878 a_n2661_42282# a_3080_42308# 0.161683f
C879 a_15765_45572# a_16115_45572# 0.20669f
C880 a_15599_45572# a_16680_45572# 0.102355f
C881 a_10809_44734# a_11691_44458# 0.354084f
C882 a_5937_45572# a_5883_43914# 0.454323f
C883 a_2324_44458# a_n2661_44458# 0.134417f
C884 a_12549_44172# a_19321_45002# 0.238866f
C885 a_8912_37509# a_11206_38545# 1.26605f
C886 a_19862_44208# a_20922_43172# 0.164553f
C887 a_n881_46662# a_5937_45572# 0.195456f
C888 a_8128_46384# a_7920_46348# 0.197919f
C889 a_n97_42460# a_5934_30871# 0.221607f
C890 a_n2312_40392# a_n2302_40160# 0.151095f
C891 a_n2433_44484# a_n2267_44484# 0.730194f
C892 a_16327_47482# a_18909_45814# 0.16767f
C893 a_4915_47217# a_2437_43646# 0.114772f
C894 a_2698_46116# a_2804_46116# 0.313533f
C895 a_5342_30871# a_14456_42282# 0.160195f
C896 a_9801_43940# VDD 0.19512f
C897 a_5883_43914# a_8333_44056# 0.152643f
C898 a_n913_45002# a_14579_43548# 0.239851f
C899 a_20916_46384# VDD 0.302226f
C900 a_22612_30879# C10_N_btm 1.5848f
C901 a_8199_44636# a_8568_45546# 0.141772f
C902 a_n971_45724# a_n2661_42834# 0.165951f
C903 a_n2438_43548# a_n2293_42834# 0.138621f
C904 a_12545_42858# VDD 0.285703f
C905 a_19328_44172# a_19478_44306# 0.188181f
C906 a_6165_46155# VDD 0.204296f
C907 a_11823_42460# a_15143_45578# 0.120787f
C908 a_8199_44636# a_n2661_43370# 0.126664f
C909 a_19332_42282# VDD 0.227361f
C910 a_n1151_42308# a_n743_46660# 0.195953f
C911 a_10210_45822# VDD 0.323342f
C912 a_16147_45260# a_16019_45002# 0.186254f
C913 a_3357_43084# a_3065_45002# 0.316449f
C914 a_12549_44172# a_13059_46348# 0.808395f
C915 a_13507_46334# a_12741_44636# 0.137731f
C916 a_n1151_42308# a_11189_46129# 0.12414f
C917 a_21101_45002# VDD 0.2903f
C918 a_13556_45296# a_13720_44458# 0.212774f
C919 a_9482_43914# a_15004_44636# 0.34299f
C920 a_9290_44172# a_12281_43396# 0.36475f
C921 a_10227_46804# a_14113_42308# 0.627404f
C922 a_22612_30879# a_20205_31679# 0.111294f
C923 a_16023_47582# VDD 0.201413f
C924 a_14539_43914# a_11967_42832# 0.512158f
C925 a_n1435_47204# CLK 1.41989f
C926 a_768_44030# a_9482_43914# 0.77718f
C927 a_167_45260# a_n357_42282# 0.148401f
C928 a_n2293_46634# a_3065_45002# 0.102991f
C929 a_8685_42308# a_9223_42460# 0.166964f
C930 a_6194_45824# a_6511_45714# 0.102325f
C931 a_10809_44734# a_2437_43646# 0.13907f
C932 a_5379_42460# VDD 0.213136f
C933 a_n1435_47204# a_13717_47436# 0.196889f
C934 a_n4209_38502# a_n3565_38502# 6.84323f
C935 a_n2433_43396# a_n2129_43609# 0.283605f
C936 a_n23_45546# VDD 0.150941f
C937 a_7499_43078# a_1307_43914# 0.109806f
C938 a_16327_47482# a_16243_43396# 0.295263f
C939 EN_VIN_BSTR_P C0_P_btm 0.12803f
C940 C10_P_btm C8_P_btm 2.07867f
C941 a_4915_47217# a_765_45546# 0.169406f
C942 a_171_46873# a_n2661_46098# 0.168482f
C943 a_22889_38993# VDD 0.495671f
C944 a_14797_45144# VDD 0.124624f
C945 a_n2661_45010# a_742_44458# 0.694478f
C946 a_13885_46660# a_14035_46660# 0.25868f
C947 a_17609_46634# a_17829_46910# 0.111805f
C948 a_2063_45854# a_2711_45572# 0.185507f
C949 a_15227_44166# a_17339_46660# 0.524034f
C950 a_n443_46116# a_n443_42852# 0.145452f
C951 a_20766_44850# VDD 0.197657f
C952 a_1307_43914# a_3600_43914# 0.153686f
C953 a_17970_44736# a_18287_44626# 0.102355f
C954 a_5343_44458# a_7640_43914# 0.152634f
C955 a_7287_43370# VDD 0.457521f
C956 a_1606_42308# a_1755_42282# 0.278431f
C957 a_8492_46660# VDD 0.273866f
C958 a_n1079_45724# a_n755_45592# 0.109544f
C959 a_n863_45724# a_n357_42282# 0.172013f
C960 a_380_45546# a_n1099_45572# 0.148825f
C961 a_n4064_40160# a_n2302_40160# 0.249627f
C962 a_n971_45724# a_584_46384# 0.152617f
C963 a_n2293_43922# a_5649_42852# 1.78418f
C964 a_15765_45572# a_16333_45814# 0.17072f
C965 a_3483_46348# a_16979_44734# 0.173123f
C966 a_n443_42852# a_3537_45260# 0.567413f
C967 VDAC_N a_11206_38545# 0.15219f
C968 a_768_44030# a_13747_46662# 0.434325f
C969 a_8912_37509# VDAC_P 3.15325f
C970 a_8685_43396# a_10341_43396# 2.41562f
C971 a_17715_44484# a_17737_43940# 0.289085f
C972 a_10775_45002# a_10951_45334# 0.185422f
C973 a_n1613_43370# a_5937_45572# 0.117604f
C974 a_8037_42858# a_8952_43230# 0.118759f
C975 a_4905_42826# a_5267_42460# 0.146764f
C976 a_n23_44458# VDD 0.169093f
C977 a_n1059_45260# a_n1761_44111# 0.535535f
C978 a_n2312_40392# a_n4064_40160# 0.103899f
C979 a_n755_45592# a_2982_43646# 0.221452f
C980 a_n2433_44484# a_n2129_44697# 0.130072f
C981 a_n443_46116# a_2437_43646# 0.410719f
C982 a_765_45546# a_10809_44734# 2.52248f
C983 a_9290_44172# a_11551_42558# 0.123803f
C984 a_n1059_45260# a_14579_43548# 0.250544f
C985 a_1307_43914# a_1756_43548# 0.267667f
C986 a_8199_44636# a_8162_45546# 0.119979f
C987 a_3483_46348# a_11823_42460# 0.377948f
C988 a_12549_44172# a_19778_44110# 0.294084f
C989 a_n4318_37592# a_n3420_37984# 0.404896f
C990 a_n3674_38216# a_n4064_37984# 0.65176f
C991 a_12089_42308# VDD 0.807892f
C992 a_7542_44172# a_7499_43940# 0.157633f
C993 a_5497_46414# VDD 0.200657f
C994 a_8162_45546# a_8192_45572# 0.134163f
C995 a_18907_42674# VDD 0.148872f
C996 a_n1151_42308# a_n1021_46688# 0.105326f
C997 a_n443_46116# a_n2661_46634# 0.121882f
C998 a_7754_39632# a_7754_39300# 0.296258f
C999 a_n2661_45010# a_n467_45028# 0.227953f
C1000 a_12891_46348# a_13059_46348# 0.372745f
C1001 a_4791_45118# a_5937_45572# 0.151145f
C1002 a_n1151_42308# a_9290_44172# 0.10853f
C1003 a_20916_46384# a_19692_46634# 0.117693f
C1004 a_n881_46662# a_765_45546# 0.333008f
C1005 a_21005_45260# VDD 0.184261f
C1006 a_n2661_45010# a_n2661_43922# 0.111071f
C1007 a_9482_43914# a_13720_44458# 0.188323f
C1008 a_1423_45028# a_5343_44458# 0.128331f
C1009 a_12861_44030# a_12791_45546# 0.248928f
C1010 a_22000_46634# a_20202_43084# 0.154237f
C1011 a_16327_47482# a_10193_42453# 0.163668f
C1012 a_16327_47482# VDD 2.81451f
C1013 a_10903_43370# a_13259_45724# 0.600111f
C1014 a_12891_46348# a_13556_45296# 0.29495f
C1015 a_1823_45246# a_n755_45592# 0.390511f
C1016 a_526_44458# a_n1925_42282# 0.213917f
C1017 a_8685_42308# a_8791_42308# 0.147376f
C1018 a_22400_42852# a_22485_38105# 0.198011f
C1019 a_6194_45824# a_6472_45840# 0.118423f
C1020 a_8199_44636# a_3537_45260# 0.199536f
C1021 a_5267_42460# VDD 0.170631f
C1022 a_n4209_38502# a_n4334_38528# 0.25243f
C1023 a_9313_44734# a_22959_42860# 0.174475f
C1024 a_n356_45724# VDD 0.719282f
C1025 a_n2956_37592# a_n4315_30879# 0.107228f
C1026 a_3090_45724# a_10729_43914# 0.135702f
C1027 a_20202_43084# a_20512_43084# 0.130366f
C1028 a_11823_42460# a_11963_45334# 0.110904f
C1029 a_22613_38993# VDD 0.533489f
C1030 EN_VIN_BSTR_P C1_P_btm 0.110046f
C1031 a_n443_46116# a_765_45546# 0.297346f
C1032 a_n2438_43548# a_2443_46660# 0.237765f
C1033 C10_P_btm C9_P_btm 53.3168f
C1034 a_8953_45002# CLK 0.310391f
C1035 a_14537_43396# VDD 0.779752f
C1036 a_n2956_37592# a_n4318_40392# 2.71462f
C1037 a_17609_46634# a_765_45546# 0.256159f
C1038 a_20835_44721# VDD 0.198384f
C1039 a_13887_32519# a_14097_32519# 10.5943f
C1040 a_20922_43172# a_21195_42852# 0.119168f
C1041 a_13259_45724# a_5649_42852# 1.92021f
C1042 a_1307_43914# a_2998_44172# 0.233292f
C1043 a_17970_44736# a_18248_44752# 0.117156f
C1044 a_5343_44458# a_6109_44484# 0.285594f
C1045 a_5937_45572# a_6945_45028# 0.22046f
C1046 a_2804_46116# a_2981_46116# 0.134298f
C1047 a_13925_46122# a_14840_46494# 0.118759f
C1048 a_6547_43396# VDD 0.219105f
C1049 a_8667_46634# VDD 0.39254f
C1050 a_3090_45724# a_1423_45028# 0.450367f
C1051 a_n2438_43548# a_949_44458# 1.62911f
C1052 a_n2109_47186# a_n1151_42308# 0.235661f
C1053 a_n237_47217# a_1239_47204# 0.203126f
C1054 a_n971_45724# a_2124_47436# 0.352461f
C1055 a_n785_47204# a_327_47204# 0.237391f
C1056 a_2479_44172# a_2813_43396# 0.115852f
C1057 a_15599_45572# a_16115_45572# 0.105995f
C1058 a_8199_44636# a_8701_44490# 0.25266f
C1059 a_3483_46348# a_14539_43914# 1.24006f
C1060 a_768_44030# a_13661_43548# 0.175469f
C1061 a_2684_37794# VDD 0.286899f
C1062 a_n1613_43370# a_n2661_46634# 0.279652f
C1063 a_n2497_47436# a_3090_45724# 0.16041f
C1064 VDAC_N VDAC_P 4.74149f
C1065 a_20731_45938# VDD 0.142103f
C1066 a_20202_43084# a_21381_43940# 0.108097f
C1067 a_10193_42453# a_n356_44636# 2.49128f
C1068 a_10227_46804# a_10809_44734# 0.17883f
C1069 a_18479_47436# a_6945_45028# 0.348097f
C1070 a_8605_42826# a_8387_43230# 0.209641f
C1071 a_3626_43646# a_1755_42282# 0.119352f
C1072 a_n356_44636# VDD 1.17667f
C1073 a_n97_42460# a_6123_31319# 0.182488f
C1074 a_n2293_42834# a_5891_43370# 0.669411f
C1075 a_n971_45724# a_n967_45348# 0.581053f
C1076 a_16327_47482# a_18479_45785# 0.841261f
C1077 a_2521_46116# a_2698_46116# 0.159555f
C1078 a_2982_43646# CAL_N 0.181412f
C1079 a_9165_43940# VDD 0.192035f
C1080 a_9290_44172# a_5742_30871# 0.118117f
C1081 a_19321_45002# START 0.10793f
C1082 a_1307_43914# a_1568_43370# 0.182552f
C1083 a_20843_47204# VDD 0.188032f
C1084 a_21588_30879# C9_N_btm 0.786375f
C1085 a_12379_42858# VDD 0.484153f
C1086 a_5204_45822# VDD 0.359177f
C1087 a_13163_45724# a_13527_45546# 0.124682f
C1088 a_10053_45546# a_10210_45822# 0.18824f
C1089 a_11823_42460# a_13249_42308# 0.360411f
C1090 a_13507_46334# a_11341_43940# 0.162723f
C1091 a_10227_46804# a_n881_46662# 0.146883f
C1092 a_18727_42674# VDD 0.181095f
C1093 a_n1151_42308# a_n1925_46634# 0.105874f
C1094 a_2113_38308# VDAC_Ni 0.318652f
C1095 a_n4064_40160# C10_P_btm 0.460005f
C1096 a_8697_45822# VDD 0.189893f
C1097 a_20447_31679# a_413_45260# 0.226658f
C1098 a_7499_43078# a_11827_44484# 0.104754f
C1099 a_n2109_45247# en_comp 0.108653f
C1100 a_3357_43084# a_2382_45260# 0.219664f
C1101 a_4883_46098# a_20202_43084# 0.135688f
C1102 a_2063_45854# a_10903_43370# 0.277624f
C1103 a_4791_45118# a_8199_44636# 0.14611f
C1104 a_n1613_43370# a_765_45546# 0.205521f
C1105 a_20567_45036# VDD 0.237324f
C1106 a_9482_43914# a_13076_44458# 0.103066f
C1107 a_1307_43914# a_5883_43914# 0.289388f
C1108 a_526_44458# a_3539_42460# 0.213772f
C1109 a_12861_44030# a_11823_42460# 1.2465f
C1110 a_20273_46660# a_12741_44636# 0.540506f
C1111 a_16241_47178# VDD 0.208959f
C1112 a_1176_45822# a_997_45618# 0.140567f
C1113 a_12891_46348# a_9482_43914# 0.314487f
C1114 a_8325_42308# a_8791_42308# 0.173196f
C1115 a_16721_46634# VDD 0.186443f
C1116 a_6945_45028# a_2437_43646# 2.26888f
C1117 a_n2438_43548# a_n2293_43922# 0.575621f
C1118 a_12549_44172# a_19615_44636# 0.157395f
C1119 a_3823_42558# VDD 0.170296f
C1120 a_2063_45854# a_4883_46098# 0.116597f
C1121 en_comp a_22485_38105# 0.535686f
C1122 a_3503_45724# VDD 0.129733f
C1123 a_3090_45724# a_10405_44172# 0.126512f
C1124 a_10903_43370# a_n2661_42834# 0.269313f
C1125 a_11823_42460# a_11787_45002# 0.217891f
C1126 a_22581_37893# VDD 0.902719f
C1127 EN_VIN_BSTR_P C2_P_btm 0.118072f
C1128 a_2107_46812# a_1983_46706# 0.212212f
C1129 a_n2438_43548# a_n2661_46098# 0.391488f
C1130 a_18783_43370# a_15743_43084# 0.303966f
C1131 a_14180_45002# VDD 0.151315f
C1132 a_4791_45118# a_4921_42308# 0.172224f
C1133 a_20679_44626# VDD 0.439119f
C1134 a_3232_43370# a_3499_42826# 0.339727f
C1135 a_7499_43078# a_8147_43396# 0.227361f
C1136 a_n443_46116# a_1307_43914# 0.442637f
C1137 a_13759_46122# a_14840_46494# 0.102325f
C1138 a_14493_46090# a_14275_46494# 0.209641f
C1139 a_6765_43638# VDD 0.218204f
C1140 a_14635_42282# a_14456_42282# 0.172313f
C1141 a_7927_46660# VDD 0.187888f
C1142 a_n863_45724# a_n1099_45572# 0.172847f
C1143 a_8034_45724# a_8162_45546# 0.14162f
C1144 a_13661_43548# a_13720_44458# 0.122691f
C1145 a_n2438_43548# a_742_44458# 0.171623f
C1146 a_n4315_30879# a_n2302_40160# 0.407166f
C1147 a_n4334_40480# a_n4064_40160# 0.43652f
C1148 a_n23_47502# a_327_47204# 0.140943f
C1149 a_n237_47217# a_1209_47178# 0.206644f
C1150 a_5111_44636# a_5379_42460# 0.118194f
C1151 a_15493_43940# a_19319_43548# 0.36082f
C1152 a_15903_45785# a_15765_45572# 0.205788f
C1153 a_13059_46348# a_14673_44172# 0.108306f
C1154 a_8199_44636# a_8103_44636# 0.256009f
C1155 a_12549_44172# a_13661_43548# 0.149087f
C1156 a_1107_38525# VDD 0.374783f
C1157 VDAC_N a_8912_37509# 3.43288f
C1158 a_6151_47436# a_8492_46660# 0.302615f
C1159 a_8685_43396# a_14955_43396# 0.111211f
C1160 a_3537_45260# a_1307_43914# 0.290878f
C1161 a_8037_42858# a_8387_43230# 0.225358f
C1162 a_7871_42858# a_8952_43230# 0.102355f
C1163 a_n2293_45010# a_n1899_43946# 0.18948f
C1164 a_13556_45296# a_14673_44172# 0.137701f
C1165 a_n2312_40392# a_n4315_30879# 0.389397f
C1166 a_16327_47482# a_18175_45572# 0.346603f
C1167 a_765_45546# a_6945_45028# 4.99804f
C1168 a_17517_44484# a_11967_42832# 0.342031f
C1169 a_5111_44636# a_7287_43370# 0.104641f
C1170 a_19594_46812# VDD 0.349555f
C1171 a_3090_45724# a_3357_43084# 0.546562f
C1172 a_10341_42308# VDD 0.931019f
C1173 a_5164_46348# VDD 0.717083f
C1174 a_11453_44696# a_22959_47212# 0.182671f
C1175 a_18057_42282# VDD 0.130308f
C1176 a_11599_46634# a_12891_46348# 0.150715f
C1177 a_13507_46334# a_11415_45002# 0.160889f
C1178 a_n2293_46634# a_3090_45724# 1.2853f
C1179 a_18494_42460# VDD 0.73193f
C1180 a_10807_43548# a_11323_42473# 0.109765f
C1181 a_768_44030# a_n755_45592# 0.202175f
C1182 a_3499_42826# VDD 0.333472f
C1183 a_n357_42282# a_7227_42852# 0.185359f
C1184 a_15673_47210# VDD 0.569224f
C1185 a_1138_42852# a_n357_42282# 0.325445f
C1186 a_n2497_47436# a_n699_43396# 0.355158f
C1187 a_8325_42308# a_8685_42308# 0.141819f
C1188 a_18494_42460# a_16137_43396# 0.115144f
C1189 a_16388_46812# VDD 0.797417f
C1190 a_n2293_46098# a_1307_43914# 0.107603f
C1191 a_5907_45546# a_6194_45824# 0.233657f
C1192 a_12549_44172# a_11967_42832# 0.193926f
C1193 a_3318_42354# VDD 0.203036f
C1194 a_5934_30871# C5_P_btm 0.139996f
C1195 a_3316_45546# VDD 0.428912f
C1196 a_n743_46660# a_n2661_46098# 0.414618f
C1197 a_n2438_43548# a_1799_45572# 0.137623f
C1198 EN_VIN_BSTR_P C3_P_btm 0.100325f
C1199 a_16327_47482# a_19466_46812# 0.203994f
C1200 a_13777_45326# VDD 0.145151f
C1201 a_4955_46873# a_4704_46090# 0.109136f
C1202 a_20640_44752# VDD 0.246486f
C1203 a_1307_43914# a_2675_43914# 0.453622f
C1204 a_17767_44458# a_17970_44736# 0.233657f
C1205 a_626_44172# a_453_43940# 0.163589f
C1206 a_13925_46122# a_14275_46494# 0.20669f
C1207 a_6197_43396# VDD 0.408793f
C1208 a_1184_42692# a_2123_42473# 0.107417f
C1209 a_n863_45724# a_1606_42308# 0.20593f
C1210 a_8145_46902# VDD 0.199702f
C1211 a_15227_44166# a_15415_45028# 0.222342f
C1212 a_n2293_45546# a_310_45028# 0.113595f
C1213 a_n1079_45724# a_n1099_45572# 0.15766f
C1214 a_n2497_47436# a_n1151_42308# 0.156942f
C1215 a_n2109_47186# a_2905_45572# 0.124881f
C1216 a_n4315_30879# a_n4064_40160# 0.363059f
C1217 a_5066_45546# VDD 1.34058f
C1218 a_n913_45002# a_8325_42308# 0.233489f
C1219 a_15599_45572# a_15765_45572# 0.576512f
C1220 a_12549_44172# a_5807_45002# 0.675558f
C1221 a_6886_37412# a_8912_37509# 0.339465f
C1222 a_6151_47436# a_8667_46634# 0.357581f
C1223 a_n97_42460# a_4361_42308# 0.15989f
C1224 a_21188_45572# VDD 0.288663f
C1225 a_10227_46804# a_6945_45028# 0.220094f
C1226 a_768_44030# a_3483_46348# 0.281593f
C1227 a_8037_42858# a_8605_42826# 0.178024f
C1228 a_n2293_45010# a_n1761_44111# 0.148418f
C1229 a_9482_43914# a_14673_44172# 0.42967f
C1230 a_3090_45724# a_8049_45260# 1.23904f
C1231 a_167_45260# a_2521_46116# 0.328009f
C1232 a_19321_45002# VDD 1.01574f
C1233 a_2324_44458# a_2711_45572# 0.804101f
C1234 a_526_44458# a_n863_45724# 0.801581f
C1235 a_11453_44696# a_n2661_44458# 0.174607f
C1236 a_5742_30871# a_7174_31319# 0.34728f
C1237 a_10922_42852# VDD 0.216186f
C1238 a_n2293_46634# a_1414_42308# 0.260739f
C1239 a_13487_47204# a_768_44030# 0.371206f
C1240 a_n3565_38216# a_n4209_37414# 5.88577f
C1241 a_n4315_30879# C10_P_btm 1.5848f
C1242 a_17531_42308# VDD 0.262303f
C1243 a_10193_42453# a_18184_42460# 0.216199f
C1244 a_n1059_45260# a_n913_45002# 1.19505f
C1245 a_n2472_45002# en_comp 0.117861f
C1246 a_4646_46812# a_6197_43396# 0.601282f
C1247 a_20916_46384# a_15227_44166# 0.681561f
C1248 a_13507_46334# a_20202_43084# 0.205796f
C1249 a_19594_46812# a_19692_46634# 0.134424f
C1250 a_18184_42460# VDD 2.05053f
C1251 a_9482_43914# a_12607_44458# 0.151452f
C1252 a_9290_44172# a_10341_43396# 0.157042f
C1253 a_12861_44030# a_11962_45724# 0.184706f
C1254 a_20107_46660# a_12741_44636# 0.527863f
C1255 a_768_44030# a_n357_42282# 0.175577f
C1256 a_n357_42282# a_5755_42852# 0.179701f
C1257 a_15811_47375# VDD 0.979053f
C1258 a_13259_45724# a_17701_42308# 0.137488f
C1259 a_11459_47204# DATA[5] 0.370451f
C1260 a_n746_45260# a_n2129_44697# 0.17701f
C1261 a_5932_42308# a_5742_30871# 1.14154f
C1262 a_5891_43370# a_n97_42460# 0.957548f
C1263 a_13059_46348# VDD 0.955445f
C1264 a_2903_42308# VDD 0.22017f
C1265 a_6123_31319# C4_P_btm 0.132906f
C1266 a_n2840_43370# a_n4318_39304# 0.158695f
C1267 a_3218_45724# VDD 0.133843f
C1268 a_9290_44172# a_n2293_43922# 0.369185f
C1269 a_22527_39145# VDD 0.626886f
C1270 EN_VIN_BSTR_P C4_P_btm 0.116925f
C1271 a_13556_45296# VDD 0.569056f
C1272 a_18525_43370# a_18783_43370# 0.22264f
C1273 a_9290_44172# a_n97_42460# 0.351467f
C1274 a_21588_30879# a_10809_44734# 0.110956f
C1275 a_20362_44736# VDD 0.275577f
C1276 a_1307_43914# a_895_43940# 0.754684f
C1277 a_11691_44458# a_15433_44458# 0.110923f
C1278 a_19321_45002# a_18479_45785# 0.114441f
C1279 a_13759_46122# a_14275_46494# 0.105995f
C1280 a_13925_46122# a_14493_46090# 0.17072f
C1281 a_6293_42852# VDD 0.401011f
C1282 a_7577_46660# VDD 0.249866f
C1283 a_n2661_45546# a_n755_45592# 0.14317f
C1284 a_n4315_30879# a_n4334_40480# 0.253307f
C1285 a_15599_45572# a_15903_45785# 0.161702f
C1286 a_1609_45822# a_2274_45254# 0.11737f
C1287 a_5088_37509# VDAC_P 1.15441f
C1288 a_5700_37509# a_8912_37509# 15.051701f
C1289 a_6151_47436# a_7927_46660# 0.182356f
C1290 a_21363_45546# VDD 0.36538f
C1291 a_2324_44458# a_15682_43940# 0.321744f
C1292 a_413_45260# a_1423_45028# 0.194002f
C1293 a_3232_43370# a_9482_43914# 0.129525f
C1294 a_12549_44172# a_3483_46348# 0.185475f
C1295 a_7871_42858# a_8387_43230# 0.106107f
C1296 a_3080_42308# a_2903_42308# 0.154008f
C1297 a_n746_45260# a_n745_45366# 0.119822f
C1298 a_7499_43940# VDD 0.193884f
C1299 a_5534_30871# a_12563_42308# 0.179331f
C1300 a_5883_43914# a_n2661_42282# 0.107496f
C1301 a_19466_46812# a_20528_45572# 0.157758f
C1302 a_n3674_38216# a_n3565_38216# 0.128699f
C1303 a_10991_42826# VDD 0.201891f
C1304 a_18326_43940# a_18451_43940# 0.145292f
C1305 a_4704_46090# VDD 0.225404f
C1306 a_n971_45724# a_n2129_43609# 0.173854f
C1307 SMPL_ON_N a_11453_44696# 0.147722f
C1308 a_2063_45854# a_n743_46660# 1.58762f
C1309 a_12861_44030# a_768_44030# 0.260776f
C1310 a_17303_42282# VDD 0.37938f
C1311 a_3540_43646# a_3626_43646# 0.100706f
C1312 a_n2017_45002# a_n913_45002# 0.275686f
C1313 a_n2472_45002# a_n2956_37592# 0.152938f
C1314 a_n2661_45010# en_comp 0.10363f
C1315 a_19594_46812# a_19466_46812# 0.100902f
C1316 a_2063_45854# a_11189_46129# 0.294233f
C1317 a_22959_43396# a_17364_32525# 0.156288f
C1318 a_19778_44110# VDD 0.469922f
C1319 a_9482_43914# a_8975_43940# 0.186623f
C1320 a_20202_43084# a_4361_42308# 0.472299f
C1321 a_1423_45028# a_2779_44458# 0.246285f
C1322 SMPL_ON_N a_21753_35634# 0.39912f
C1323 a_13259_45724# a_17595_43084# 0.118887f
C1324 a_15507_47210# VDD 0.441662f
C1325 a_167_45260# a_n863_45724# 0.424358f
C1326 a_9290_44172# a_13259_45724# 0.272297f
C1327 a_12891_46348# a_13017_45260# 0.210934f
C1328 a_3483_46348# a_n2661_45546# 0.163728f
C1329 a_15227_46910# VDD 0.229766f
C1330 w_1575_34946# a_n1794_35242# 3.10971f
C1331 a_3090_45724# a_11691_44458# 0.245063f
C1332 a_13661_43548# a_14673_44172# 0.36897f
C1333 a_2713_42308# VDD 0.208275f
C1334 a_2957_45546# VDD 0.192471f
C1335 a_22589_40055# VDD 1.08898f
C1336 a_19998_35138# a_21753_35634# 0.150805f
C1337 EN_VIN_BSTR_P C5_P_btm 0.115337f
C1338 a_16327_47482# a_15227_44166# 0.239667f
C1339 a_9482_43914# VDD 1.75061f
C1340 a_n97_42460# a_16795_42852# 0.126591f
C1341 a_1823_45246# a_3539_42460# 0.678673f
C1342 a_20159_44458# VDD 0.345429f
C1343 a_1307_43914# a_2479_44172# 0.300587f
C1344 a_3537_45260# a_n2661_42282# 0.105917f
C1345 a_13747_46662# a_18341_45572# 0.554429f
C1346 a_19123_46287# a_19240_46482# 0.157972f
C1347 a_3090_45724# a_n443_42852# 0.269331f
C1348 a_1823_45246# a_526_44458# 1.93329f
C1349 a_6031_43396# VDD 0.47547f
C1350 a_13291_42460# a_13070_42354# 0.155164f
C1351 a_1184_42692# a_1606_42308# 0.125247f
C1352 a_1576_42282# a_1755_42282# 0.168925f
C1353 a_7715_46873# VDD 0.414019f
C1354 a_22959_44484# a_19237_31679# 0.155744f
C1355 a_15227_44166# a_14537_43396# 0.105881f
C1356 a_n746_45260# a_n785_47204# 0.198992f
C1357 a_11967_42832# a_16547_43609# 0.176385f
C1358 a_19862_44208# a_21381_43940# 0.113704f
C1359 a_5700_37509# VDAC_N 1.09421f
C1360 a_5088_37509# a_8912_37509# 16.1906f
C1361 a_n2302_38778# VDD 0.35162f
C1362 a_3726_37500# a_11206_38545# 0.11542f
C1363 a_6151_47436# a_8145_46902# 0.178565f
C1364 a_n1151_42308# a_6755_46942# 0.142929f
C1365 a_20623_45572# VDD 0.200978f
C1366 a_n4318_40392# a_n4315_30879# 0.151169f
C1367 a_327_44734# a_626_44172# 0.120093f
C1368 a_7765_42852# a_8037_42858# 0.309282f
C1369 a_n1809_44850# VDD 0.132538f
C1370 a_n2840_44458# a_n2661_44458# 0.179135f
C1371 a_n755_45592# a_n1557_42282# 0.199254f
C1372 a_11599_46634# a_18341_45572# 0.588263f
C1373 a_2202_46116# a_167_45260# 0.159883f
C1374 a_6671_43940# VDD 0.227011f
C1375 a_13747_46662# VDD 3.70214f
C1376 a_3483_46348# a_11322_45546# 0.554731f
C1377 a_10796_42968# VDD 0.270235f
C1378 a_5663_43940# a_5829_43940# 0.143754f
C1379 a_10729_43914# a_11341_43940# 0.243062f
C1380 a_10193_42453# a_4958_30871# 0.108497f
C1381 a_4419_46090# VDD 0.664887f
C1382 VDAC_Pi a_3754_39466# 0.308867f
C1383 a_4958_30871# VDD 1.06745f
C1384 a_584_46384# a_n743_46660# 0.42078f
C1385 a_12861_44030# a_12549_44172# 1.20253f
C1386 a_2982_43646# a_3626_43646# 6.553431f
C1387 a_n2017_45002# a_n1059_45260# 6.27837f
C1388 a_3357_43084# a_413_45260# 7.24598f
C1389 a_n2661_45010# a_n2956_37592# 0.163638f
C1390 a_n2293_46098# a_n2661_42282# 0.182071f
C1391 a_4646_46812# a_6031_43396# 0.849684f
C1392 a_n1151_42308# a_8953_45546# 0.120628f
C1393 a_2063_45854# a_9290_44172# 0.655982f
C1394 a_4791_45118# a_6419_46155# 0.371259f
C1395 a_18597_46090# a_12741_44636# 0.267775f
C1396 a_768_44030# a_14035_46660# 0.270355f
C1397 VDD VCM 1.50561f
C1398 a_19321_45002# a_19466_46812# 0.130025f
C1399 a_18911_45144# VDD 0.218047f
C1400 a_9482_43914# a_10057_43914# 0.401746f
C1401 a_20202_43084# a_13467_32519# 0.333168f
C1402 a_11599_46634# a_10193_42453# 0.100544f
C1403 a_11599_46634# VDD 5.64965f
C1404 a_n2497_47436# a_949_44458# 0.127971f
C1405 a_10903_43370# a_12839_46116# 0.115226f
C1406 a_5807_45002# a_6171_45002# 0.193427f
C1407 a_n2293_46634# a_413_45260# 0.497204f
C1408 a_n2017_45002# a_19987_42826# 0.142839f
C1409 a_3090_45724# a_19113_45348# 0.128103f
C1410 a_9313_45822# a_11459_47204# 0.210847f
C1411 a_n784_42308# VCM 0.195503f
C1412 a_1848_45724# VDD 0.100884f
C1413 a_n1613_43370# a_7112_43396# 0.245085f
C1414 EN_VIN_BSTR_P C6_P_btm 0.118916f
C1415 a_10227_46804# a_14976_45028# 0.536884f
C1416 a_1123_46634# a_948_46660# 0.234322f
C1417 a_18429_43548# a_18525_43370# 0.419086f
C1418 a_13507_46334# a_22400_42852# 0.235269f
C1419 a_n443_42852# a_1414_42308# 0.193113f
C1420 a_n2661_45010# a_n2267_44484# 0.260289f
C1421 a_n443_46116# a_n23_45546# 0.118272f
C1422 a_18597_46090# a_16375_45002# 0.105669f
C1423 a_768_44030# a_n1925_42282# 0.145535f
C1424 a_6755_46942# a_12741_44636# 0.131965f
C1425 a_19615_44636# VDD 0.203841f
C1426 a_1307_43914# a_2127_44172# 0.127867f
C1427 a_n2442_46660# a_n2302_39866# 0.161638f
C1428 a_13759_46122# a_13925_46122# 0.576786f
C1429 a_1576_42282# a_1606_42308# 0.176925f
C1430 a_3080_42308# VCM 0.148824f
C1431 a_7411_46660# VDD 0.41059f
C1432 a_n746_45260# a_n23_47502# 0.148631f
C1433 a_n971_45724# a_n785_47204# 0.385455f
C1434 a_11967_42832# a_16243_43396# 0.269605f
C1435 a_8049_45260# a_n2293_42834# 0.224469f
C1436 a_5700_37509# a_6886_37412# 0.13762f
C1437 a_5088_37509# VDAC_N 0.420254f
C1438 a_4338_37500# a_8912_37509# 0.331796f
C1439 a_n4064_38528# VDD 1.69517f
C1440 a_n237_47217# a_8270_45546# 0.552109f
C1441 a_6151_47436# a_7577_46660# 0.578207f
C1442 a_20841_45814# VDD 0.209907f
C1443 a_17538_32519# a_17364_32525# 9.64512f
C1444 a_n2293_43922# a_5932_42308# 0.178011f
C1445 a_2382_45260# a_1307_43914# 0.53878f
C1446 a_13259_45724# a_3422_30871# 0.587088f
C1447 a_6755_46942# a_13607_46688# 0.129798f
C1448 a_7871_42858# a_8037_42858# 0.772842f
C1449 a_n2840_44458# a_n4318_40392# 0.161548f
C1450 a_n357_42282# a_n1557_42282# 0.384406f
C1451 a_1823_45246# a_167_45260# 0.155648f
C1452 a_12891_46348# a_13249_42308# 0.166217f
C1453 a_19123_46287# a_18985_46122# 0.215692f
C1454 a_n971_45724# a_n913_45002# 0.101346f
C1455 a_n746_45260# a_n1059_45260# 0.138039f
C1456 a_13661_43548# a_10193_42453# 0.211481f
C1457 a_5829_43940# VDD 0.156797f
C1458 a_13661_43548# VDD 3.93017f
C1459 a_20193_45348# a_15493_43940# 0.10893f
C1460 a_7499_43078# a_10341_42308# 0.42152f
C1461 a_3537_45260# a_7287_43370# 0.400907f
C1462 a_20202_43084# a_21335_42336# 0.227943f
C1463 a_3483_46348# a_10490_45724# 0.207668f
C1464 a_4185_45028# a_10193_42453# 3.16135f
C1465 a_15764_42576# a_4958_30871# 0.413236f
C1466 a_10835_43094# VDD 0.43308f
C1467 a_18079_43940# a_18326_43940# 0.152347f
C1468 a_4185_45028# VDD 1.65665f
C1469 a_11962_45724# a_13163_45724# 0.113317f
C1470 a_12427_45724# a_12791_45546# 0.124682f
C1471 a_8049_45260# a_413_45260# 0.140877f
C1472 a_22731_47423# SMPL_ON_N 0.194951f
C1473 a_16327_47482# a_n881_46662# 0.195459f
C1474 a_5257_43370# a_4905_42826# 0.254437f
C1475 a_n443_42852# a_n699_43396# 0.333516f
C1476 a_n1151_42308# a_5937_45572# 0.11638f
C1477 a_4791_45118# a_6165_46155# 0.291653f
C1478 VDD VREF_GND 0.482759f
C1479 a_4646_46812# a_7411_46660# 0.266058f
C1480 a_375_42282# a_n699_43396# 0.127058f
C1481 a_14311_47204# RST_Z 0.184572f
C1482 a_18248_44752# a_17517_44484# 0.561898f
C1483 a_14955_47212# VDD 0.301751f
C1484 a_n2497_47436# a_742_44458# 0.153038f
C1485 a_1823_45246# a_n863_45724# 0.207189f
C1486 a_n2438_43548# en_comp 0.915368f
C1487 a_167_45260# a_n2293_45546# 0.681309f
C1488 a_8515_42308# a_8685_42308# 0.108744f
C1489 a_5934_30871# a_8791_42308# 0.223675f
C1490 a_3600_43914# a_3499_42826# 0.125876f
C1491 a_19466_46812# a_19778_44110# 0.116901f
C1492 a_3483_46348# a_6171_45002# 0.153232f
C1493 a_2063_45854# a_10949_43914# 0.129837f
C1494 a_997_45618# VDD 0.12359f
C1495 a_20202_43084# a_3422_30871# 0.527141f
C1496 a_n1613_43370# a_7287_43370# 0.337957f
C1497 a_22537_40625# VDD 0.534319f
C1498 EN_VIN_BSTR_P C7_P_btm 0.115875f
C1499 a_171_46873# a_288_46660# 0.159893f
C1500 a_10227_46804# a_3090_45724# 0.320681f
C1501 a_13159_45002# VDD 0.321035f
C1502 a_21381_43940# a_21195_42852# 0.238789f
C1503 a_16547_43609# a_16664_43396# 0.161376f
C1504 a_11967_42832# a_15803_42450# 0.258862f
C1505 a_4791_45118# a_5379_42460# 0.197725f
C1506 a_10193_42453# a_11967_42832# 0.752992f
C1507 a_n2661_45010# a_n2129_44697# 0.18531f
C1508 a_n443_46116# a_n356_45724# 0.113738f
C1509 a_768_44030# a_526_44458# 0.341438f
C1510 a_11967_42832# VDD 2.67441f
C1511 a_14539_43914# a_16979_44734# 0.132799f
C1512 a_626_44172# a_644_44056# 0.126386f
C1513 a_n2442_46660# a_n4064_39616# 0.224005f
C1514 a_n357_42282# a_n3674_37592# 0.327427f
C1515 a_n863_45724# a_1184_42692# 0.563857f
C1516 a_5257_43370# VDD 0.922495f
C1517 a_n2293_45546# a_n863_45724# 0.17075f
C1518 a_3090_45724# a_1307_43914# 2.66267f
C1519 a_n2109_47186# a_584_46384# 0.352889f
C1520 a_n971_45724# a_n23_47502# 0.225828f
C1521 a_n746_45260# a_n237_47217# 0.285294f
C1522 a_1337_46116# VDD 0.20087f
C1523 a_11967_42832# a_16137_43396# 0.300696f
C1524 a_13661_43548# a_14021_43940# 0.103152f
C1525 a_n2293_46634# a_11341_43940# 0.487839f
C1526 a_3090_45724# a_18579_44172# 0.16932f
C1527 a_5088_37509# a_6886_37412# 0.136505f
C1528 a_3726_37500# a_8912_37509# 0.267651f
C1529 a_6491_46660# a_5257_43370# 0.1719f
C1530 a_n2946_38778# VDD 0.383009f
C1531 a_20273_45572# VDD 0.571099f
C1532 a_13507_46334# a_22165_42308# 0.126777f
C1533 a_n2438_43548# a_n2157_42858# 0.266513f
C1534 a_18597_46090# a_18819_46122# 0.230891f
C1535 a_7871_42858# a_7765_42852# 0.379881f
C1536 a_18989_43940# VDD 0.342796f
C1537 a_11599_46634# a_18175_45572# 0.844188f
C1538 a_1138_42852# a_167_45260# 0.250282f
C1539 a_1823_45246# a_2202_46116# 0.25354f
C1540 a_19123_46287# a_18819_46122# 0.172712f
C1541 a_n971_45724# a_n1059_45260# 0.322275f
C1542 a_5745_43940# VDD 0.144352f
C1543 a_5807_45002# VDD 1.75047f
C1544 a_5111_44636# a_6031_43396# 0.207345f
C1545 a_4223_44672# a_8333_44056# 0.122173f
C1546 a_n1925_42282# a_n2661_45546# 0.181908f
C1547 a_12549_44172# a_16922_45042# 0.803336f
C1548 a_3483_46348# a_8746_45002# 0.605995f
C1549 a_10518_42984# VDD 0.273357f
C1550 a_n2810_45572# a_n3565_38502# 0.409424f
C1551 a_3699_46348# VDD 0.208984f
C1552 a_12741_44636# a_11691_44458# 0.81445f
C1553 a_n2497_47436# a_n447_43370# 0.192476f
C1554 a_11962_45724# a_12791_45546# 0.124167f
C1555 a_12427_45724# a_11823_42460# 0.17307f
C1556 a_7754_39964# a_7754_39632# 0.296522f
C1557 a_n1151_42308# a_n2661_46634# 0.832521f
C1558 a_15143_45578# VDD 0.12071f
C1559 a_n2109_45247# a_n2017_45002# 0.193269f
C1560 a_n2840_45002# a_n2810_45028# 0.161831f
C1561 a_n2293_46634# a_10341_43396# 2.04894f
C1562 a_13747_46662# a_19466_46812# 0.869986f
C1563 a_n1151_42308# a_8199_44636# 0.161616f
C1564 a_19321_45002# a_15227_44166# 0.145462f
C1565 VDD VREF 4.8299f
C1566 C10_N_btm VCM 10.5945f
C1567 a_18315_45260# VDD 0.12623f
C1568 a_n443_42852# a_15493_43940# 0.301211f
C1569 a_14311_47204# VDD 0.241476f
C1570 a_3357_43084# a_n97_42460# 0.113127f
C1571 a_18114_32519# a_19237_31679# 8.86269f
C1572 a_5807_45002# a_5691_45260# 0.19412f
C1573 a_2324_44458# a_10586_45546# 0.436403f
C1574 a_1138_42852# a_n863_45724# 0.135594f
C1575 a_17364_32525# EN_VIN_BSTR_N 1.00234f
C1576 a_8515_42308# a_8325_42308# 0.134955f
C1577 a_5934_30871# a_8685_42308# 0.186981f
C1578 a_16867_43762# VDD 0.132317f
C1579 a_3483_46348# a_3232_43370# 0.220803f
C1580 a_n3420_39072# a_n4064_38528# 7.47287f
C1581 a_1666_39043# a_2112_39137# 0.553829f
C1582 a_1273_38525# a_2684_37794# 0.224374f
C1583 a_5932_42308# C3_P_btm 0.121156f
C1584 a_n755_45592# VDD 2.41485f
C1585 a_n2438_43548# a_n2267_43396# 0.120634f
C1586 a_n2293_46634# a_n97_42460# 0.108602f
C1587 a_n443_42852# a_n2293_42834# 1.60683f
C1588 a_n1613_43370# a_6547_43396# 0.154311f
C1589 a_22589_40599# VDD 0.821011f
C1590 a_11599_46634# a_19466_46812# 0.453656f
C1591 a_n1151_42308# a_765_45546# 1.7705f
C1592 a_13017_45260# VDD 0.263701f
C1593 a_21381_43940# a_21356_42826# 0.196864f
C1594 a_4791_45118# a_5267_42460# 0.138738f
C1595 a_n2661_45010# a_n2433_44484# 0.217176f
C1596 a_3877_44458# a_4185_45028# 0.338483f
C1597 a_20916_46384# a_21137_46414# 0.118131f
C1598 a_7227_42852# a_7309_42852# 0.171361f
C1599 a_19339_43156# a_19164_43230# 0.233657f
C1600 a_526_44458# a_5111_42852# 0.265994f
C1601 a_1307_43914# a_1414_42308# 0.147738f
C1602 a_5807_45002# a_18479_45785# 0.174313f
C1603 a_1184_42692# a_961_42354# 0.100246f
C1604 a_n755_45592# a_n784_42308# 0.711298f
C1605 a_n2438_43548# a_n2267_44484# 0.120608f
C1606 a_n815_47178# a_n785_47204# 0.123817f
C1607 a_n971_45724# a_n237_47217# 0.134971f
C1608 a_n913_45002# a_5934_30871# 0.126791f
C1609 a_4338_37500# a_6886_37412# 1.95816f
C1610 a_6151_47436# a_7411_46660# 0.330209f
C1611 a_n3420_38528# VDD 0.522772f
C1612 a_5088_37509# a_5700_37509# 1.48771f
C1613 a_n971_45724# a_8270_45546# 0.251101f
C1614 a_20107_45572# VDD 0.458237f
C1615 a_14401_32519# a_17364_32525# 7.49646f
C1616 a_n97_42460# a_743_42282# 0.107736f
C1617 a_413_45260# a_375_42282# 0.112554f
C1618 a_n1741_47186# a_12839_46116# 0.113988f
C1619 a_16327_47482# a_6945_45028# 0.111399f
C1620 a_7227_42852# a_7765_42852# 0.118623f
C1621 a_18374_44850# VDD 0.203584f
C1622 a_n755_45592# a_3080_42308# 0.237742f
C1623 a_12549_44172# a_13163_45724# 0.172293f
C1624 a_16131_47204# VDD 0.142103f
C1625 a_20193_45348# a_11341_43940# 0.21261f
C1626 a_3483_46348# a_10193_42453# 0.359034f
C1627 a_10083_42826# VDD 0.461256f
C1628 a_n4318_38216# a_n4209_38216# 0.135236f
C1629 a_17973_43940# a_18079_43940# 0.419086f
C1630 a_17730_32519# a_17538_32519# 9.37324f
C1631 a_3483_46348# VDD 2.29096f
C1632 a_11962_45724# a_11823_42460# 0.177935f
C1633 a_n2438_43548# a_n2065_43946# 0.265458f
C1634 a_13381_47204# a_12549_44172# 0.135267f
C1635 a_4958_30871# C9_N_btm 0.209166f
C1636 a_14495_45572# VDD 0.238674f
C1637 a_2896_43646# a_2982_43646# 0.100706f
C1638 w_1575_34946# VDD 1.59781f
C1639 a_2437_43646# a_413_45260# 0.20387f
C1640 VDD VIN_N 1.44851f
C1641 C9_N_btm VCM 6.06251f
C1642 C10_N_btm VREF_GND 10.3207f
C1643 a_3877_44458# a_5257_43370# 0.142219f
C1644 a_17719_45144# VDD 0.1297f
C1645 a_22591_43396# a_14209_32519# 0.158752f
C1646 a_9482_43914# a_10157_44484# 0.321004f
C1647 a_13487_47204# VDD 0.273369f
C1648 a_12861_44030# RST_Z 0.290405f
C1649 a_9067_47204# DATA[4] 0.354356f
C1650 a_n443_42852# a_n13_43084# 0.13203f
C1651 a_1823_45246# a_n2293_45546# 0.234971f
C1652 a_5934_30871# a_8325_42308# 0.173576f
C1653 a_14513_46634# VDD 0.223375f
C1654 a_n357_42282# a_10193_42453# 0.634772f
C1655 a_2351_42308# VDD 0.188239f
C1656 a_1273_38525# a_1107_38525# 0.236832f
C1657 a_6151_47436# a_14955_47212# 0.192081f
C1658 a_n1151_42308# a_10227_46804# 0.458569f
C1659 SMPL_ON_P a_n2312_40392# 4.89949f
C1660 a_n357_42282# VDD 1.90108f
C1661 a_n1613_43370# a_6765_43638# 0.164755f
C1662 CAL_N VDD 26.0839f
C1663 a_11206_38545# RST_Z 0.382319f
C1664 EN_VIN_BSTR_N a_19998_35138# 0.573047f
C1665 a_18194_35068# a_19250_35138# 0.559484f
C1666 EN_VIN_BSTR_P C9_P_btm 0.226529f
C1667 a_33_46660# a_948_46660# 0.117156f
C1668 a_11963_45334# VDD 0.229584f
C1669 a_16409_43396# a_15743_43084# 0.586918f
C1670 a_n881_46662# a_5066_45546# 0.801045f
C1671 a_20916_46384# a_20708_46348# 0.189941f
C1672 a_18588_44850# VDD 0.132317f
C1673 a_n357_42282# a_16137_43396# 1.09442f
C1674 a_16112_44458# a_14539_43914# 0.13299f
C1675 a_526_44458# a_4520_42826# 0.247914f
C1676 a_1307_43914# a_1467_44172# 0.228571f
C1677 a_11415_45002# a_8049_45260# 0.426371f
C1678 a_4915_47217# a_13556_45296# 0.146395f
C1679 a_22165_42308# a_21887_42336# 0.110763f
C1680 a_22591_44484# a_17730_32519# 0.156987f
C1681 a_n863_45724# a_1067_42314# 0.289393f
C1682 a_11415_45002# a_19479_31679# 0.224531f
C1683 a_n971_45724# a_n746_45260# 0.393354f
C1684 a_20269_44172# a_19319_43548# 0.12985f
C1685 a_n443_42852# a_n37_45144# 0.137227f
C1686 a_3726_37500# a_6886_37412# 0.702909f
C1687 a_n3690_38528# VDD 0.363159f
C1688 a_4338_37500# a_5700_37509# 2.69237f
C1689 a_4883_46098# a_2107_46812# 2.95673f
C1690 a_7229_43940# a_7705_45326# 0.203098f
C1691 a_n443_46116# a_5066_45546# 0.130975f
C1692 a_18443_44721# VDD 0.193515f
C1693 a_18285_46348# a_17957_46116# 0.12677f
C1694 a_3537_45260# a_6197_43396# 0.337459f
C1695 a_19466_46812# a_20273_45572# 0.328586f
C1696 a_8049_45260# a_13259_45724# 0.895805f
C1697 a_5257_43370# a_5111_44636# 0.22597f
C1698 a_8952_43230# VDD 0.273404f
C1699 a_n1059_45260# a_16245_42852# 0.130348f
C1700 a_3147_46376# VDD 0.341038f
C1701 a_n4064_40160# EN_VIN_BSTR_P 0.149512f
C1702 a_13249_42308# VDD 0.653917f
C1703 a_20512_43084# a_19987_42826# 0.11919f
C1704 a_5807_45002# a_19466_46812# 0.178376f
C1705 a_n1151_42308# a_8016_46348# 0.580516f
C1706 a_4791_45118# a_5164_46348# 0.42219f
C1707 a_10227_46804# a_12741_44636# 0.188309f
C1708 C10_N_btm VREF 14.773f
C1709 C8_N_btm VCM 2.61094f
C1710 C9_N_btm VREF_GND 5.18245f
C1711 VDD VIN_P 1.46295f
C1712 a_n881_46662# a_13059_46348# 0.642888f
C1713 a_15095_43370# a_15567_42826# 0.167909f
C1714 a_n443_42852# a_11341_43940# 0.51832f
C1715 a_9482_43914# a_9838_44484# 0.175591f
C1716 a_20202_43084# a_743_42282# 0.135735f
C1717 a_526_44458# a_n1557_42282# 0.31675f
C1718 a_1307_43914# a_4223_44672# 0.747516f
C1719 a_n1441_43940# VDD 0.142719f
C1720 a_16979_44734# a_17517_44484# 0.109784f
C1721 a_12861_44030# VDD 3.56689f
C1722 a_13717_47436# RST_Z 4.51263f
C1723 a_6575_47204# DATA[4] 0.15718f
C1724 a_18114_32519# a_17730_32519# 9.15095f
C1725 a_5807_45002# a_5111_44636# 0.204193f
C1726 a_19700_43370# VDD 0.28578f
C1727 a_14180_46812# VDD 0.755623f
C1728 a_3357_43084# a_n2293_42282# 0.146926f
C1729 a_n2956_38680# a_n2946_38778# 0.14863f
C1730 a_18579_44172# a_15493_43940# 0.377126f
C1731 a_n4318_39768# a_n3674_39768# 3.06574f
C1732 a_2711_45572# a_4099_45572# 0.176427f
C1733 a_n3420_39072# a_n3420_38528# 0.127439f
C1734 a_n1920_47178# a_n2312_39304# 0.157528f
C1735 a_6151_47436# a_14311_47204# 0.136645f
C1736 a_2123_42473# VDD 0.1936f
C1737 a_n2293_43922# a_5534_30871# 0.271171f
C1738 a_310_45028# VDD 0.360949f
C1739 a_n2438_43548# a_n2433_43396# 0.415301f
C1740 a_11599_46634# a_15227_44166# 0.101252f
C1741 a_11206_38545# VDD 8.87267f
C1742 a_11530_34132# a_19998_35138# 0.201872f
C1743 EN_VIN_BSTR_N a_19250_35138# 0.651354f
C1744 EN_VIN_BSTR_P C10_P_btm 0.320569f
C1745 VDAC_P RST_Z 0.158793f
C1746 a_601_46902# a_383_46660# 0.209641f
C1747 a_n97_42460# a_5534_30871# 0.109695f
C1748 a_11787_45002# VDD 0.153399f
C1749 a_17499_43370# a_17324_43396# 0.234322f
C1750 a_16292_46812# a_16388_46812# 0.318472f
C1751 a_5755_42852# a_5837_42852# 0.171361f
C1752 a_n443_42852# a_10341_43396# 0.23026f
C1753 a_1307_43914# a_1115_44172# 0.115939f
C1754 a_n2293_46098# a_5066_45546# 0.140248f
C1755 a_4915_47217# a_9482_43914# 0.269756f
C1756 a_1067_42314# a_961_42354# 0.13675f
C1757 a_n784_42308# a_2123_42473# 0.216332f
C1758 a_n2438_43548# a_n2433_44484# 0.421822f
C1759 a_14976_45028# a_14797_45144# 0.137651f
C1760 a_n452_47436# a_n746_45260# 0.187792f
C1761 a_8495_42852# VDD 0.132018f
C1762 a_3065_45002# a_3823_42558# 0.198186f
C1763 a_n913_45002# a_6123_31319# 0.21316f
C1764 a_5257_43370# a_3905_42865# 0.106385f
C1765 a_3316_45546# a_3429_45260# 0.142842f
C1766 a_16375_45002# a_1307_43914# 0.101951f
C1767 a_584_46384# a_3457_43396# 0.120485f
C1768 a_n443_42852# a_n143_45144# 0.104427f
C1769 a_n3565_38502# VDD 0.762011f
C1770 a_4338_37500# a_5088_37509# 0.896828f
C1771 a_3726_37500# a_5700_37509# 0.574743f
C1772 a_2063_45854# a_6755_46942# 0.131005f
C1773 a_14401_32519# a_14209_32519# 10.7535f
C1774 a_n97_42460# a_4190_30871# 0.140814f
C1775 a_5891_43370# a_9223_42460# 0.13879f
C1776 a_8685_43396# a_9145_43396# 0.201058f
C1777 a_7229_43940# a_6709_45028# 0.136786f
C1778 a_4791_45118# a_5066_45546# 0.238282f
C1779 a_768_44030# a_1823_45246# 0.287407f
C1780 a_21588_30879# a_21076_30879# 8.21286f
C1781 a_18287_44626# VDD 0.389383f
C1782 en_comp a_3422_30871# 0.357746f
C1783 a_n443_42852# a_n97_42460# 0.822111f
C1784 a_18285_46348# a_18189_46348# 0.118603f
C1785 a_12549_44172# a_11823_42460# 0.624462f
C1786 a_n971_45724# a_n2293_45010# 0.549225f
C1787 a_20202_43084# a_13258_32519# 0.685083f
C1788 a_19466_46812# a_20107_45572# 0.283769f
C1789 a_5257_43370# a_5147_45002# 0.836149f
C1790 a_9127_43156# VDD 0.468721f
C1791 a_17737_43940# a_17973_43940# 0.22264f
C1792 a_2804_46116# VDD 0.159351f
C1793 a_20202_43084# a_20193_45348# 0.116706f
C1794 a_17124_42282# VDD 0.28176f
C1795 a_12465_44636# a_22223_47212# 0.175138f
C1796 a_4915_47217# a_13747_46662# 0.710704f
C1797 a_584_46384# a_n2293_46634# 0.374996f
C1798 a_13904_45546# VDD 0.135068f
C1799 a_n443_42852# a_742_44458# 0.168627f
C1800 C10_N_btm VIN_N 3.66034f
C1801 VDD CLK 0.49309f
C1802 a_13661_43548# a_15227_44166# 0.805606f
C1803 C9_N_btm VREF 7.369471f
C1804 C7_N_btm VCM 1.58335f
C1805 C8_N_btm VREF_GND 2.58605f
C1806 a_5907_46634# a_5732_46660# 0.233657f
C1807 a_15095_43370# a_5342_30871# 0.238762f
C1808 a_1307_43914# a_2779_44458# 0.332183f
C1809 a_9290_44172# a_13667_43396# 0.136018f
C1810 a_1847_42826# a_2351_42308# 0.120686f
C1811 a_16979_44734# a_17061_44734# 0.171361f
C1812 a_13717_47436# VDD 0.314317f
C1813 a_n1435_47204# RST_Z 0.179508f
C1814 a_2437_43646# a_n97_42460# 0.201806f
C1815 a_n443_42852# a_n901_43156# 0.367747f
C1816 a_19268_43646# VDD 0.237793f
C1817 a_14035_46660# VDD 0.363878f
C1818 a_n2017_45002# a_18249_42858# 0.545311f
C1819 a_n1059_45260# a_17333_42852# 0.270324f
C1820 a_n2956_38680# a_n3420_38528# 0.233147f
C1821 a_3483_46348# a_5111_44636# 0.340106f
C1822 a_n237_47217# a_4883_46098# 0.181672f
C1823 a_1606_42308# RST_Z 1.44945f
C1824 a_1755_42282# VDD 0.215277f
C1825 a_1666_39587# a_2684_37794# 0.565516f
C1826 en_comp a_7174_31319# 5.65156f
C1827 a_n1099_45572# VDD 0.89411f
C1828 a_13259_45724# a_11691_44458# 0.337184f
C1829 a_4883_46098# a_8270_45546# 0.278829f
C1830 a_10227_46804# a_12816_46660# 0.253017f
C1831 EN_VIN_BSTR_N a_18194_35068# 0.336225f
C1832 a_11530_34132# a_19250_35138# 0.481434f
C1833 VDAC_P VDD 5.18919f
C1834 a_n133_46660# a_948_46660# 0.102355f
C1835 a_33_46660# a_383_46660# 0.20669f
C1836 a_n2438_43548# a_2107_46812# 0.111283f
C1837 a_10951_45334# VDD 0.226705f
C1838 a_16243_43396# a_15743_43084# 0.600668f
C1839 a_n971_45724# a_2711_45572# 0.214535f
C1840 a_18249_42858# a_19164_43230# 0.118759f
C1841 a_n2442_46660# a_n3565_39590# 0.134948f
C1842 a_13259_45724# a_4190_30871# 0.271537f
C1843 a_n2956_39768# a_n2946_39866# 0.14868f
C1844 a_584_46384# a_626_44172# 0.450256f
C1845 a_1067_42314# a_1184_42692# 0.147283f
C1846 a_n357_42282# a_n473_42460# 0.179066f
C1847 a_22485_44484# a_22591_44484# 0.15878f
C1848 a_12549_44172# a_14539_43914# 0.110516f
C1849 a_n2438_43548# a_n2661_44458# 0.136664f
C1850 a_n2472_45546# a_n2293_45546# 0.171197f
C1851 a_n452_47436# a_n971_45724# 0.330438f
C1852 a_n2109_47186# a_1209_47178# 0.226908f
C1853 a_3065_45002# a_3318_42354# 0.146272f
C1854 a_n1925_42282# VDD 0.728256f
C1855 en_comp a_5932_42308# 0.23313f
C1856 a_9313_44734# a_13887_32519# 0.191376f
C1857 a_15227_44166# a_11967_42832# 0.132673f
C1858 a_3316_45546# a_3065_45002# 0.141454f
C1859 a_n4334_38528# VDD 0.385889f
C1860 a_3726_37500# a_5088_37509# 0.189392f
C1861 a_n881_46662# a_13747_46662# 0.550574f
C1862 a_7276_45260# a_6709_45028# 0.215102f
C1863 a_6755_46942# a_11901_46660# 0.587021f
C1864 a_n2661_46634# a_11415_45002# 0.494836f
C1865 a_16327_47482# a_19900_46494# 0.216811f
C1866 a_18248_44752# VDD 0.251171f
C1867 a_765_45546# a_17957_46116# 0.133328f
C1868 a_1176_45822# a_1138_42852# 0.41217f
C1869 a_12549_44172# a_12427_45724# 0.152925f
C1870 a_n746_45260# a_n2661_45010# 0.400342f
C1871 a_3737_43940# VDD 0.18423f
C1872 a_n1925_42282# a_n784_42308# 0.235613f
C1873 a_18479_45785# a_19268_43646# 0.12682f
C1874 a_3483_46348# a_9049_44484# 0.117501f
C1875 a_8387_43230# VDD 0.200672f
C1876 a_22485_44484# a_20974_43370# 0.101193f
C1877 a_2698_46116# VDD 0.195879f
C1878 a_2324_44458# a_1423_45028# 0.154419f
C1879 a_18479_47436# a_20935_43940# 0.207572f
C1880 a_526_44458# a_3232_43370# 0.461444f
C1881 a_12741_44636# a_11827_44484# 0.305294f
C1882 a_11322_45546# a_11823_42460# 0.133185f
C1883 a_11599_46634# a_n881_46662# 0.100714f
C1884 a_n746_45260# a_171_46873# 0.120194f
C1885 a_11459_47204# a_11309_47204# 0.183357f
C1886 a_3422_30871# a_21671_42860# 0.199876f
C1887 a_13527_45546# VDD 0.1902f
C1888 a_n2472_45002# a_n2293_45010# 0.177252f
C1889 C9_N_btm VIN_N 1.82823f
C1890 a_n443_46116# a_4419_46090# 0.20069f
C1891 VDD EN_OFFSET_CAL 0.489629f
C1892 a_13661_43548# a_18834_46812# 0.1407f
C1893 C8_N_btm VREF 3.6701f
C1894 C7_N_btm VREF_GND 1.61142f
C1895 a_n2497_47436# a_2324_44458# 0.796031f
C1896 C6_N_btm VCM 0.877241f
C1897 a_18114_32519# EN_VIN_BSTR_N 0.149512f
C1898 a_n97_42460# a_13291_42460# 0.419357f
C1899 a_16922_45042# VDD 1.54713f
C1900 a_15095_43370# a_15279_43071# 0.105784f
C1901 SMPL_ON_P a_n4315_30879# 3.7092f
C1902 a_n1925_42282# a_3080_42308# 0.897997f
C1903 a_526_44458# a_4905_42826# 0.202895f
C1904 a_1307_43914# a_11341_43940# 2.31482f
C1905 a_n1435_47204# VDD 0.267875f
C1906 a_22612_30879# a_413_45260# 0.11791f
C1907 a_1823_45246# a_n2661_45546# 0.181403f
C1908 a_15743_43084# VDD 0.572249f
C1909 a_13885_46660# VDD 0.499249f
C1910 a_n2017_45002# a_17333_42852# 0.314084f
C1911 a_n755_45592# a_7499_43078# 0.157526f
C1912 a_15227_44166# a_18315_45260# 0.272047f
C1913 a_3483_46348# a_5147_45002# 0.363215f
C1914 a_1169_39043# comp_n 0.3874f
C1915 a_1606_42308# VDD 0.629724f
C1916 a_6151_47436# a_12861_44030# 0.39397f
C1917 a_14401_32519# a_20974_43370# 0.118041f
C1918 a_380_45546# VDD 0.154763f
C1919 a_10807_43548# a_10695_43548# 0.159782f
C1920 a_n913_45002# a_21613_42308# 0.259761f
C1921 a_2324_44458# a_6109_44484# 0.101116f
C1922 a_8746_45002# a_8953_45002# 0.257529f
C1923 a_10227_46804# a_10341_43396# 0.188948f
C1924 a_n1613_43370# a_6031_43396# 0.308901f
C1925 a_16327_47482# a_3090_45724# 1.00134f
C1926 a_10227_46804# a_12991_46634# 0.349162f
C1927 a_11530_34132# a_18194_35068# 0.419364f
C1928 VDAC_N RST_Z 0.154233f
C1929 a_8912_37509# VDD 18.3523f
C1930 a_33_46660# a_601_46902# 0.17072f
C1931 a_n743_46660# a_2107_46812# 0.72755f
C1932 a_10775_45002# VDD 0.148349f
C1933 a_n2661_42282# a_n2840_42282# 0.173771f
C1934 a_15559_46634# a_13059_46348# 0.167936f
C1935 a_5111_42852# a_5193_42852# 0.171361f
C1936 a_18817_42826# a_18599_43230# 0.209641f
C1937 a_n2956_39768# a_n3420_39616# 0.233256f
C1938 a_10903_43370# a_13351_46090# 0.181897f
C1939 a_n784_42308# a_1606_42308# 15.027599f
C1940 a_3539_42460# VDD 0.363092f
C1941 a_n913_45002# a_4361_42308# 0.250497f
C1942 a_n2472_45546# a_n2956_38216# 0.157892f
C1943 a_20202_43084# a_2437_43646# 0.129143f
C1944 a_3090_45724# a_14537_43396# 0.530123f
C1945 COMP_P a_22537_40625# 0.120662f
C1946 a_15493_43396# a_19319_43548# 0.120111f
C1947 a_526_44458# VDD 2.35177f
C1948 a_n913_45002# a_6761_42308# 0.350952f
C1949 a_10227_46804# a_n97_42460# 0.18445f
C1950 a_n4209_38502# VDD 0.811731f
C1951 a_3726_37500# a_4338_37500# 0.212154f
C1952 a_7276_45260# a_7229_43940# 0.322065f
C1953 a_1799_45572# a_765_45546# 0.225248f
C1954 a_16327_47482# a_20075_46420# 0.270434f
C1955 a_3080_42308# a_1606_42308# 4.87174f
C1956 a_17970_44736# VDD 0.27753f
C1957 a_2063_45854# a_2437_43646# 0.392331f
C1958 a_14401_32519# EN_VIN_BSTR_N 0.814814f
C1959 a_16922_45042# a_14021_43940# 0.11663f
C1960 a_7499_43078# a_10083_42826# 0.375624f
C1961 a_3232_43370# a_3626_43646# 0.204337f
C1962 a_1307_43914# a_n97_42460# 0.23336f
C1963 a_3483_46348# a_7499_43078# 0.207714f
C1964 a_8605_42826# VDD 0.204898f
C1965 a_2521_46116# VDD 0.163553f
C1966 a_n2497_47436# a_n2267_43396# 0.222725f
C1967 a_16104_42674# VDD 0.134357f
C1968 a_2063_45854# a_n2661_46634# 1.75382f
C1969 a_4915_47217# a_5807_45002# 0.766023f
C1970 a_7754_40130# a_7754_39964# 0.301877f
C1971 a_3422_30871# a_21195_42852# 0.289298f
C1972 a_13163_45724# VDD 0.322298f
C1973 a_n2661_45010# a_n2293_45010# 0.400159f
C1974 C8_N_btm VIN_N 0.907642f
C1975 VDD DATA[5] 0.504354f
C1976 C7_N_btm VREF 1.818f
C1977 a_10227_46804# a_11415_45002# 0.139042f
C1978 C6_N_btm VREF_GND 0.836236f
C1979 C5_N_btm VCM 0.719982f
C1980 a_4955_46873# a_5072_46660# 0.17431f
C1981 a_22223_43396# a_13887_32519# 0.154411f
C1982 a_12281_43396# a_12089_42308# 0.210903f
C1983 a_n913_45002# a_5891_43370# 0.255618f
C1984 a_1307_43914# a_742_44458# 0.355379f
C1985 a_15227_44166# a_3483_46348# 0.595533f
C1986 a_6755_46942# a_15682_46116# 0.116442f
C1987 a_7227_47204# DATA[3] 0.357377f
C1988 a_13381_47204# VDD 0.130765f
C1989 a_n2438_43548# a_n2017_45002# 0.29197f
C1990 a_5934_30871# a_8515_42308# 0.222946f
C1991 a_18783_43370# VDD 0.289099f
C1992 a_n2956_38680# a_n3565_38502# 0.302523f
C1993 a_4185_45028# a_3537_45260# 1.06643f
C1994 a_n357_42282# a_7499_43078# 0.259858f
C1995 a_2324_44458# a_3357_43084# 0.216574f
C1996 a_15227_44166# a_17719_45144# 0.187414f
C1997 a_9290_44172# a_n913_45002# 0.632534f
C1998 a_n2288_47178# a_n2312_40392# 0.153632f
C1999 a_6151_47436# a_13717_47436# 0.17202f
C2000 a_n452_45724# VDD 0.112977f
C2001 a_11823_42460# a_6171_45002# 0.123118f
C2002 a_11530_34132# EN_VIN_BSTR_N 1.06713f
C2003 a_n3420_37440# VIN_P 0.143165f
C2004 a_n881_46662# a_5257_43370# 0.447042f
C2005 VDAC_N VDD 4.61811f
C2006 a_n133_46660# a_383_46660# 0.105995f
C2007 a_2063_45854# a_765_45546# 1.71006f
C2008 a_10227_46804# a_12251_46660# 0.188053f
C2009 a_8953_45002# VDD 1.24336f
C2010 a_16409_43396# a_17324_43396# 0.118759f
C2011 a_584_46384# a_n443_42852# 1.36389f
C2012 a_10227_46804# a_13259_45724# 0.335001f
C2013 a_15368_46634# a_13059_46348# 0.101997f
C2014 a_7765_42852# a_8292_43218# 0.157652f
C2015 a_18083_42858# a_19164_43230# 0.101963f
C2016 a_18249_42858# a_18599_43230# 0.210876f
C2017 a_10193_42453# a_3626_43646# 0.13905f
C2018 a_526_44458# a_2075_43172# 0.227071f
C2019 a_584_46384# a_375_42282# 0.480677f
C2020 a_10903_43370# a_12594_46348# 0.169312f
C2021 a_3626_43646# VDD 0.340378f
C2022 a_5275_47026# VDD 0.135766f
C2023 a_768_44030# a_13720_44458# 0.178939f
C2024 a_n2661_45546# a_n2956_38216# 0.15505f
C2025 a_20202_43084# a_21513_45002# 0.13666f
C2026 COMP_P a_22589_40599# 0.204694f
C2027 a_n815_47178# a_n452_47436# 0.107449f
C2028 a_n2109_47186# a_n785_47204# 0.43597f
C2029 a_18451_43940# a_18533_43940# 0.171361f
C2030 a_2981_46116# VDD 0.111597f
C2031 a_12549_44172# a_768_44030# 0.490163f
C2032 a_2112_39137# VDD 0.28506f
C2033 a_n881_46662# a_5807_45002# 0.243322f
C2034 a_n4209_39304# VREF 0.195875f
C2035 a_20974_43370# a_5649_42852# 0.186094f
C2036 a_8696_44636# a_11691_44458# 0.141053f
C2037 a_6431_45366# a_6709_45028# 0.112564f
C2038 a_n881_46662# a_3699_46348# 0.203393f
C2039 a_6755_46942# a_11735_46660# 0.61229f
C2040 a_16327_47482# a_19335_46494# 0.155998f
C2041 a_17767_44458# VDD 0.348803f
C2042 a_17339_46660# a_18189_46348# 0.170772f
C2043 a_765_45546# a_17715_44484# 0.117636f
C2044 a_1208_46090# a_1176_45822# 0.141891f
C2045 a_584_46384# a_2437_43646# 0.302508f
C2046 a_12089_42308# a_11551_42558# 0.109508f
C2047 a_11827_44484# a_11341_43940# 0.231114f
C2048 a_n356_44636# a_1414_42308# 0.179164f
C2049 a_n1151_42308# a_n23_44458# 0.101137f
C2050 a_3483_46348# a_8568_45546# 0.137016f
C2051 a_10903_43370# a_2711_45572# 0.213719f
C2052 a_8037_42858# VDD 0.344922f
C2053 a_9313_44734# a_8685_43396# 0.124273f
C2054 a_167_45260# VDD 1.41955f
C2055 a_3483_46348# a_n2661_43370# 0.953959f
C2056 a_n2497_47436# a_n2129_43609# 0.216536f
C2057 a_18597_46090# a_19862_44208# 0.536021f
C2058 a_10490_45724# a_12427_45724# 0.108721f
C2059 a_11525_45546# a_11652_45724# 0.138143f
C2060 a_11322_45546# a_11962_45724# 0.270736f
C2061 a_3754_39964# VDAC_Pi 0.296508f
C2062 a_n237_47217# a_n743_46660# 0.192378f
C2063 a_11031_47542# a_11309_47204# 0.110775f
C2064 a_4699_43561# a_3539_42460# 0.109444f
C2065 a_12791_45546# VDD 0.205486f
C2066 a_4817_46660# a_5732_46660# 0.118759f
C2067 a_n743_46660# a_8270_45546# 0.274248f
C2068 C7_N_btm VIN_N 1.52449f
C2069 VDD DATA[4] 0.326957f
C2070 C6_N_btm VREF 1.41944f
C2071 a_11453_44696# a_20273_46660# 0.545219f
C2072 C5_N_btm VREF_GND 0.676559f
C2073 C4_N_btm VCM 0.716447f
C2074 a_n1059_45260# a_5891_43370# 0.186322f
C2075 a_n1925_42282# a_4235_43370# 0.199349f
C2076 a_9290_44172# a_9145_43396# 0.103991f
C2077 a_327_44734# a_n23_44458# 0.141544f
C2078 a_6755_46942# a_2324_44458# 0.155169f
C2079 a_6851_47204# DATA[3] 0.146601f
C2080 a_14539_43914# a_14673_44172# 0.205935f
C2081 a_n863_45724# a_2905_42968# 0.269475f
C2082 a_11459_47204# VDD 0.34771f
C2083 a_18525_43370# VDD 0.263553f
C2084 a_n2017_45002# a_17701_42308# 0.132871f
C2085 a_7542_44172# a_7845_44172# 0.137004f
C2086 a_2063_45854# a_10227_46804# 0.186188f
C2087 a_n2497_47436# a_n2312_40392# 0.194574f
C2088 a_6575_47204# a_9067_47204# 0.210614f
C2089 a_10807_43548# a_9145_43396# 0.290878f
C2090 a_n863_45724# VDD 1.89058f
C2091 a_10180_45724# a_8953_45002# 0.107499f
C2092 a_6886_37412# VDD 0.235486f
C2093 a_171_46873# a_33_46660# 0.207108f
C2094 a_n1925_46634# a_2107_46812# 1.12874f
C2095 a_12861_44030# a_15227_44166# 0.810382f
C2096 a_10227_46804# a_12469_46902# 0.181535f
C2097 a_8191_45002# VDD 0.39677f
C2098 a_16977_43638# a_16759_43396# 0.209641f
C2099 a_n443_46116# a_n755_45592# 0.651643f
C2100 a_14976_45028# a_13059_46348# 0.209989f
C2101 a_18249_42858# a_18817_42826# 0.16939f
C2102 a_7229_43940# a_7281_43914# 0.164835f
C2103 a_n443_42852# a_14205_43396# 0.118229f
C2104 a_n2956_39768# a_n3565_39590# 0.302561f
C2105 a_526_44458# a_1847_42826# 0.154735f
C2106 a_10903_43370# a_12005_46116# 0.277468f
C2107 a_3540_43646# VDD 0.209044f
C2108 a_n863_45724# a_n784_42308# 0.358682f
C2109 a_8199_44636# a_8696_44636# 0.265919f
C2110 a_768_44030# a_13076_44458# 0.132449f
C2111 a_n2810_45572# a_n2956_38216# 6.20057f
C2112 a_22775_42308# a_22485_38105# 0.330766f
C2113 a_7309_42852# VDD 0.177437f
C2114 a_20193_45348# a_22165_42308# 0.252856f
C2115 a_4791_45118# a_5257_43370# 0.36404f
C2116 a_12891_46348# a_768_44030# 0.193145f
C2117 a_n881_46662# a_3483_46348# 0.5947f
C2118 a_13507_46334# a_13351_46090# 0.214666f
C2119 a_16327_47482# a_19553_46090# 0.172776f
C2120 a_16979_44734# VDD 0.256327f
C2121 a_1307_43914# a_n2661_42834# 3.43601f
C2122 a_13556_45296# a_15433_44458# 0.1084f
C2123 a_n913_45002# a_3422_30871# 0.145467f
C2124 a_n881_46662# a_14495_45572# 0.170589f
C2125 a_2455_43940# VDD 0.144352f
C2126 a_3232_43370# a_2982_43646# 0.416054f
C2127 a_7765_42852# VDD 0.333322f
C2128 a_2202_46116# VDD 0.20904f
C2129 a_11415_45002# a_11827_44484# 0.169126f
C2130 a_526_44458# a_5111_44636# 0.338508f
C2131 a_10490_45724# a_11962_45724# 0.114064f
C2132 a_10193_42453# a_11823_42460# 0.235429f
C2133 a_11322_45546# a_11652_45724# 0.26844f
C2134 a_n2497_47436# a_n2433_43396# 0.173242f
C2135 a_13487_47204# a_n881_46662# 0.108977f
C2136 a_4791_45118# a_5807_45002# 0.129041f
C2137 a_11823_42460# VDD 4.44574f
C2138 a_8696_44636# a_16751_45260# 0.265287f
C2139 a_5385_46902# a_5167_46660# 0.209641f
C2140 a_n2661_46634# a_11813_46116# 0.162517f
C2141 a_19321_45002# a_3090_45724# 0.163821f
C2142 a_n1151_42308# a_5204_45822# 0.487224f
C2143 C6_N_btm VIN_N 0.391905f
C2144 a_5807_45002# a_16292_46812# 0.202526f
C2145 C5_N_btm VREF 0.987144f
C2146 C4_N_btm VREF_GND 0.671882f
C2147 C3_N_btm VCM 0.716273f
C2148 a_13747_46662# a_15368_46634# 0.110984f
C2149 VDD DATA[3] 0.309692f
C2150 a_14579_43548# a_15279_43071# 0.108607f
C2151 a_5649_42852# a_22223_43396# 0.165664f
C2152 a_13678_32519# a_13887_32519# 10.751599f
C2153 a_8270_45546# a_9290_44172# 0.433963f
C2154 a_4915_47217# a_13249_42308# 0.161597f
C2155 a_9313_45822# VDD 0.5747f
C2156 a_6151_47436# DATA[5] 0.19492f
C2157 a_n443_42852# a_n1853_43023# 0.141267f
C2158 a_18429_43548# VDD 0.163446f
C2159 a_n1059_45260# a_16795_42852# 0.182174f
C2160 a_n2956_38680# a_n4209_38502# 0.235751f
C2161 a_3483_46348# a_3537_45260# 0.605469f
C2162 a_1823_45246# a_3232_43370# 0.344002f
C2163 a_20512_43084# a_5649_42852# 0.141324f
C2164 a_n1079_45724# VDD 0.172275f
C2165 a_10227_46804# a_15095_43370# 0.264777f
C2166 a_12861_44030# a_15681_43442# 0.137136f
C2167 a_19431_45546# a_19256_45572# 0.233657f
C2168 a_5700_37509# VDD 1.0734f
C2169 a_11599_46634# a_15368_46634# 0.320705f
C2170 a_n133_46660# a_33_46660# 0.580914f
C2171 VDAC_N C10_N_btm 0.883474p
C2172 a_16243_43396# a_17324_43396# 0.102355f
C2173 a_16409_43396# a_16759_43396# 0.20669f
C2174 a_7705_45326# VDD 0.211554f
C2175 a_4646_46812# a_7765_42852# 0.122773f
C2176 a_1823_45246# a_4905_42826# 0.110836f
C2177 a_3090_45724# a_13059_46348# 0.167043f
C2178 a_n443_46116# a_n357_42282# 0.153614f
C2179 a_18083_42858# a_18599_43230# 0.113784f
C2180 a_11827_44484# a_n2661_43922# 0.32722f
C2181 a_10193_42453# a_2982_43646# 0.231527f
C2182 a_584_46384# a_1307_43914# 0.314947f
C2183 a_5937_45572# a_2324_44458# 0.407894f
C2184 a_3090_45724# a_3218_45724# 0.100752f
C2185 a_2982_43646# VDD 1.40372f
C2186 a_n2293_43922# a_n2661_42282# 0.133253f
C2187 a_13507_46334# a_9313_44734# 0.145766f
C2188 a_5837_42852# VDD 0.1774f
C2189 a_n1741_47186# a_n971_45724# 0.157081f
C2190 a_n2109_47186# a_n237_47217# 0.730469f
C2191 a_n913_45002# a_5932_42308# 0.220872f
C2192 a_n357_42282# a_3537_45260# 0.200175f
C2193 a_12891_46348# a_12549_44172# 0.309821f
C2194 a_n2312_39304# a_n2442_46660# 0.15211f
C2195 a_n356_44636# a_5742_30871# 0.120133f
C2196 a_n97_42460# a_16823_43084# 0.205258f
C2197 a_526_44458# a_3905_42865# 0.321601f
C2198 a_10193_42453# a_14539_43914# 0.278963f
C2199 a_12861_44030# a_10809_44734# 0.156561f
C2200 a_10249_46116# a_11186_47026# 0.172467f
C2201 a_14539_43914# VDD 0.873589f
C2202 a_9482_43914# a_15433_44458# 0.20244f
C2203 a_13556_45296# a_14815_43914# 0.378519f
C2204 a_472_46348# a_1176_45822# 0.146555f
C2205 a_2253_43940# VDD 0.156797f
C2206 a_8953_45546# a_9223_42460# 0.166987f
C2207 a_14113_42308# a_16522_42674# 0.183181f
C2208 a_7871_42858# VDD 0.395222f
C2209 a_1823_45246# VDD 1.7584f
C2210 a_3600_43914# a_3737_43940# 0.126609f
C2211 a_18479_47436# a_19862_44208# 0.138185f
C2212 a_12861_44030# a_n881_46662# 0.135351f
C2213 a_n971_45724# a_n743_46660# 0.122713f
C2214 a_9313_45822# a_9804_47204# 0.171044f
C2215 a_12427_45724# VDD 0.33808f
C2216 a_n2840_45002# a_n2661_45010# 0.189331f
C2217 a_4817_46660# a_5167_46660# 0.218775f
C2218 a_n1925_46634# a_8270_45546# 0.109762f
C2219 a_n1151_42308# a_5164_46348# 0.110485f
C2220 C5_N_btm VIN_N 0.502041f
C2221 C4_N_btm VREF 0.98728f
C2222 C3_N_btm VREF_GND 0.67174f
C2223 C2_N_btm VCM 0.716172f
C2224 a_n1741_47186# a_12594_46348# 0.150956f
C2225 VDD DATA[2] 0.3216f
C2226 a_4651_46660# a_5732_46660# 0.102355f
C2227 a_14309_45028# VDD 0.189806f
C2228 a_526_44458# a_4093_43548# 0.107158f
C2229 a_1423_45028# a_n2661_44458# 0.164701f
C2230 a_6755_46942# a_15015_46420# 0.133517f
C2231 a_n3674_39768# VDD 0.398971f
C2232 a_6545_47178# DATA[3] 0.178561f
C2233 a_n863_45724# a_1847_42826# 0.216819f
C2234 a_11031_47542# VDD 0.214104f
C2235 a_4915_47217# CLK 0.198293f
C2236 a_n2497_47436# a_n2661_44458# 0.138848f
C2237 a_17324_43396# VDD 0.274722f
C2238 a_6123_31319# a_5934_30871# 15.8951f
C2239 a_15227_44166# a_16922_45042# 0.533576f
C2240 a_1184_42692# VDD 0.813074f
C2241 a_n3565_39304# a_n4209_38502# 5.79402f
C2242 a_n2293_45546# VDD 2.06545f
C2243 a_10227_46804# a_14205_43396# 0.422372f
C2244 a_5088_37509# VDD 1.15925f
C2245 VDAC_N C9_N_btm 0.44188p
C2246 a_n2438_43548# a_33_46660# 0.588568f
C2247 a_n133_46660# a_171_46873# 0.163873f
C2248 a_12861_44030# a_17609_46634# 0.183853f
C2249 a_16409_43396# a_16977_43638# 0.17072f
C2250 a_6709_45028# VDD 0.390566f
C2251 a_4646_46812# a_7871_42858# 0.26422f
C2252 a_15227_44166# a_15743_43084# 0.513622f
C2253 a_17333_42852# a_18249_42858# 0.311255f
C2254 a_n2956_39768# a_n4209_39590# 0.334714f
C2255 a_8199_44636# a_2324_44458# 0.412215f
C2256 a_3090_45724# a_2957_45546# 0.167712f
C2257 a_2896_43646# VDD 0.208317f
C2258 a_564_42282# a_n1794_35242# 0.156633f
C2259 a_5732_46660# VDD 0.277366f
C2260 a_526_44458# a_7499_43078# 0.2203f
C2261 a_10586_45546# a_2711_45572# 0.295169f
C2262 a_12891_46348# a_13076_44458# 0.182315f
C2263 a_768_44030# a_12607_44458# 0.215512f
C2264 a_5193_42852# VDD 0.187605f
C2265 a_n2109_47186# a_n746_45260# 0.295988f
C2266 comp_n VDD 0.504807f
C2267 a_n2312_40392# a_n2442_46660# 5.91846f
C2268 a_18799_45938# VDD 0.132317f
C2269 a_n2293_43922# a_5379_42460# 0.4571f
C2270 a_20974_43370# a_4361_42308# 0.122936f
C2271 a_3232_43370# a_7229_43940# 0.180766f
C2272 a_n1613_43370# a_8952_43230# 0.213002f
C2273 a_n1151_42308# a_5066_45546# 0.5423f
C2274 a_16327_47482# a_18819_46122# 0.324239f
C2275 a_14579_43548# a_14635_42282# 0.124652f
C2276 a_16112_44458# VDD 0.182397f
C2277 a_n1557_42282# a_n1794_35242# 0.865968f
C2278 a_n743_46660# a_2711_45572# 0.525746f
C2279 a_1443_43940# VDD 0.144342f
C2280 a_n3674_38216# a_n3420_38528# 0.152701f
C2281 a_7227_42852# VDD 0.254613f
C2282 a_1138_42852# VDD 0.397518f
C2283 a_12741_44636# a_18494_42460# 0.114105f
C2284 a_21496_47436# a_4883_46098# 0.257837f
C2285 a_2113_38308# VDAC_Pi 0.170941f
C2286 a_11962_45724# VDD 0.210594f
C2287 VDD DATA[1] 0.321585f
C2288 C4_N_btm VIN_N 0.50261f
C2289 C3_N_btm VREF 0.984942f
C2290 C2_N_btm VREF_GND 0.671742f
C2291 C1_N_btm VCM 0.716121f
C2292 a_n1741_47186# a_12005_46116# 0.174477f
C2293 a_4817_46660# a_5385_46902# 0.170485f
C2294 a_13747_46662# a_3090_45724# 0.139869f
C2295 a_13507_46334# a_22000_46634# 0.183978f
C2296 a_13661_43548# a_14976_45028# 0.162789f
C2297 a_3877_44458# a_6540_46812# 0.244975f
C2298 a_13678_32519# a_5649_42852# 0.506367f
C2299 w_11334_34010# a_18194_35068# 0.799648f
C2300 a_21363_46634# a_21188_46660# 0.233657f
C2301 a_2063_45854# a_10907_45822# 0.22153f
C2302 a_n4318_39768# VDD 0.469044f
C2303 a_9863_47436# VDD 0.207794f
C2304 a_n863_45724# a_791_42968# 0.338631f
C2305 a_n2438_43548# a_n2661_45010# 0.220364f
C2306 a_15368_46634# a_15143_45578# 0.105334f
C2307 a_768_44030# a_3232_43370# 0.224083f
C2308 a_17499_43370# VDD 0.453381f
C2309 a_6123_31319# a_7963_42308# 0.192155f
C2310 a_n913_45002# a_5342_30871# 0.122483f
C2311 a_3090_45724# a_18911_45144# 0.190188f
C2312 a_13507_46334# a_20512_43084# 0.497215f
C2313 a_1576_42282# VDD 0.26017f
C2314 a_n2956_38216# VDD 0.484692f
C2315 a_n2293_43922# a_12089_42308# 0.183316f
C2316 a_16327_47482# a_10341_43396# 0.159266f
C2317 a_9290_44172# a_9313_44734# 0.140741f
C2318 EN_VIN_BSTR_P a_n217_35174# 0.651354f
C2319 a_4338_37500# VDD 0.525635f
C2320 a_3726_37500# RST_Z 1.60318f
C2321 a_4915_47217# a_13885_46660# 0.179458f
C2322 VDAC_N C8_N_btm 0.220913p
C2323 a_10227_46804# a_11735_46660# 0.54163f
C2324 a_11599_46634# a_3090_45724# 0.133107f
C2325 a_16243_43396# a_16759_43396# 0.106647f
C2326 a_7229_43940# VDD 0.821851f
C2327 a_3877_44458# a_1823_45246# 0.231164f
C2328 a_n443_46116# a_n1099_45572# 0.368941f
C2329 a_2107_46812# a_9625_46129# 0.184645f
C2330 a_18083_42858# a_18249_42858# 0.699797f
C2331 a_12883_44458# a_13076_44458# 0.142643f
C2332 a_12607_44458# a_13720_44458# 0.122704f
C2333 a_18597_46090# a_n913_45002# 0.126328f
C2334 COMP_P a_1606_42308# 2.67743f
C2335 a_5907_46634# VDD 0.341121f
C2336 a_n913_45002# a_743_42282# 0.25834f
C2337 a_768_44030# a_8975_43940# 0.124155f
C2338 a_n2840_45546# a_n2661_45546# 0.175179f
C2339 a_4649_42852# VDD 0.194775f
C2340 SMPL_ON_P a_n1605_47204# 0.194856f
C2341 a_n2109_47186# a_n971_45724# 1.21934f
C2342 a_16327_47482# a_n97_42460# 0.113034f
C2343 a_3316_45546# a_413_45260# 0.110075f
C2344 a_2063_45854# a_9863_46634# 0.10786f
C2345 a_8530_39574# CAL_N 0.644218f
C2346 a_1666_39043# VDD 2.8964f
C2347 a_n2312_39304# a_n2661_46634# 0.105298f
C2348 a_n2661_42282# a_n2293_42282# 1.04835f
C2349 a_10903_43370# a_12429_44172# 0.116356f
C2350 a_n1613_43370# a_9127_43156# 0.267842f
C2351 a_20916_46384# a_20202_43084# 0.181561f
C2352 a_12861_44030# a_6945_45028# 0.108969f
C2353 a_19321_45002# a_12741_44636# 0.113088f
C2354 a_n2497_47436# a_n2017_45002# 0.125552f
C2355 a_472_46348# a_805_46414# 0.360492f
C2356 a_1241_43940# VDD 0.162129f
C2357 a_768_44030# VDD 1.53454f
C2358 a_7499_43078# a_8037_42858# 0.160087f
C2359 a_8953_45546# a_8685_42308# 0.250058f
C2360 a_4646_46812# a_7229_43940# 0.104864f
C2361 a_5755_42852# VDD 0.179985f
C2362 a_11823_42460# a_15051_42282# 0.367924f
C2363 a_1176_45822# VDD 0.781481f
C2364 a_10193_42453# a_11652_45724# 0.197229f
C2365 a_2324_44458# a_1307_43914# 0.129761f
C2366 a_10490_45724# a_11322_45546# 0.246478f
C2367 a_13507_46334# a_4883_46098# 4.09671f
C2368 a_n971_45724# a_n1925_46634# 0.163523f
C2369 a_9863_47436# a_9804_47204# 0.109361f
C2370 a_11652_45724# VDD 0.155048f
C2371 a_13507_46334# a_5649_42852# 0.136078f
C2372 a_n2293_46634# a_9145_43396# 0.238561f
C2373 a_16327_47482# a_11415_45002# 0.94171f
C2374 a_13661_43548# a_3090_45724# 0.177565f
C2375 C3_N_btm VIN_N 0.455045f
C2376 C2_N_btm VREF 0.987884f
C2377 VDD DATA[0] 1.05526f
C2378 a_4651_46660# a_5167_46660# 0.102946f
C2379 C0_N_btm VCM 0.717064f
C2380 C1_N_btm VREF_GND 0.673422f
C2381 a_526_44458# a_1568_43370# 0.220609f
C2382 w_11334_34010# EN_VIN_BSTR_N 3.97937f
C2383 a_3090_45724# a_4185_45028# 0.770164f
C2384 a_9313_45822# a_9049_44484# 0.119007f
C2385 a_7845_44172# VDD 0.11772f
C2386 a_9067_47204# VDD 0.47483f
C2387 a_4915_47217# DATA[5] 0.121371f
C2388 a_10903_43370# a_10586_45546# 0.238199f
C2389 a_6755_46942# a_15903_45785# 0.192397f
C2390 a_16759_43396# VDD 0.191873f
C2391 a_n356_44636# a_n97_42460# 1.46232f
C2392 a_1067_42314# VDD 0.128996f
C2393 a_n2472_45546# VDD 0.290266f
C2394 a_10227_46804# a_14579_43548# 0.118896f
C2395 a_18479_45785# a_18596_45572# 0.183223f
C2396 a_18341_45572# a_19256_45572# 0.116691f
C2397 a_n2438_43548# a_n133_46660# 0.848709f
C2398 a_n1057_35174# a_n217_35174# 0.481434f
C2399 a_3726_37500# VDD 0.341303f
C2400 VDAC_N C7_N_btm 0.11042p
C2401 a_16547_43609# a_16409_43396# 0.206231f
C2402 a_4905_42826# a_5111_42852# 0.105155f
C2403 a_n913_45002# a_20193_45348# 0.224918f
C2404 a_19963_31679# a_19721_31679# 9.01086f
C2405 a_16327_47482# a_13259_45724# 0.584328f
C2406 a_17517_44484# VDD 2.99662f
C2407 a_18083_42858# a_17333_42852# 0.284837f
C2408 a_742_44458# a_n356_44636# 0.207503f
C2409 a_12607_44458# a_13076_44458# 0.200168f
C2410 a_11189_46129# a_10903_43370# 0.151119f
C2411 a_5167_46660# VDD 0.203378f
C2412 a_22315_44484# a_22485_44484# 0.109468f
C2413 a_n1059_45260# a_743_42282# 0.198704f
C2414 a_n2840_45546# a_n2810_45572# 0.162234f
C2415 a_2107_46812# a_9028_43914# 0.110155f
C2416 a_3090_45724# a_11967_42832# 0.12811f
C2417 a_1169_39043# VDD 0.505762f
C2418 a_n2312_39304# a_n2956_39768# 5.91067f
C2419 a_4883_46098# a_n743_46660# 5.6639f
C2420 a_19256_45572# VDD 0.27151f
C2421 a_21381_43940# a_4361_42308# 0.195418f
C2422 a_10903_43370# a_11750_44172# 0.135933f
C2423 a_n1613_43370# a_8387_43230# 0.163582f
C2424 a_3232_43370# a_5205_44484# 0.217288f
C2425 a_10227_46804# a_14840_46494# 0.275527f
C2426 a_n443_46116# a_526_44458# 0.366438f
C2427 a_13720_44458# VDD 0.202097f
C2428 a_19479_31679# a_19237_31679# 9.049419f
C2429 a_2711_45572# a_19319_43548# 0.225335f
C2430 a_12549_44172# a_10193_42453# 0.116594f
C2431 a_12549_44172# VDD 3.08339f
C2432 a_3537_45260# a_3539_42460# 0.264936f
C2433 a_n4318_38216# a_n3420_38528# 0.31769f
C2434 a_n3674_38680# a_n4064_38528# 0.557806f
C2435 a_5111_42852# VDD 0.178652f
C2436 a_11823_42460# a_14113_42308# 0.103699f
C2437 a_1208_46090# VDD 0.178097f
C2438 a_15227_44166# a_16979_44734# 0.181002f
C2439 a_526_44458# a_3537_45260# 0.938783f
C2440 a_13507_46334# a_21496_47436# 0.167302f
C2441 a_11525_45546# VDD 0.133093f
C2442 a_n755_45592# a_5343_44458# 0.349527f
C2443 a_1823_45246# a_3905_42865# 0.218008f
C2444 VDD CLK_DATA 0.422202f
C2445 a_16327_47482# a_20202_43084# 0.475502f
C2446 a_4955_46873# a_4817_46660# 0.318259f
C2447 C2_N_btm VIN_N 0.502408f
C2448 C1_N_btm VREF 0.98698f
C2449 a_11453_44696# a_18285_46348# 0.236771f
C2450 C0_dummy_N_btm VCM 0.311452f
C2451 C0_N_btm VREF_GND 0.350401f
C2452 a_21855_43396# a_13678_32519# 0.17881f
C2453 a_526_44458# a_1049_43396# 0.121121f
C2454 w_11334_34010# a_11530_34132# 37.749f
C2455 a_20411_46873# a_20528_46660# 0.170785f
C2456 a_16795_42852# a_16877_42852# 0.171361f
C2457 a_7542_44172# VDD 0.412456f
C2458 a_6575_47204# VDD 1.32036f
C2459 a_16977_43638# VDD 0.206333f
C2460 a_7227_42308# a_6123_31319# 0.189956f
C2461 a_4190_30871# C10_P_btm 0.446355f
C2462 a_n913_45002# a_5534_30871# 0.274894f
C2463 a_8953_45546# a_n1059_45260# 0.318691f
C2464 a_12741_44636# a_9482_43914# 0.101234f
C2465 a_n1151_42308# a_11599_46634# 0.116147f
C2466 a_n1794_35242# VDD 3.20904f
C2467 a_n2661_45546# VDD 0.733118f
C2468 a_18909_45814# a_18691_45572# 0.209641f
C2469 a_n743_46660# a_n133_46660# 0.205551f
C2470 VDAC_N C6_N_btm 55.2142f
C2471 a_n1696_35090# a_n217_35174# 0.559484f
C2472 a_n1057_35174# EN_VIN_BSTR_P 1.06713f
C2473 a_5205_44484# VDD 0.508148f
C2474 a_16243_43396# a_16409_43396# 0.575934f
C2475 a_4905_42826# a_4520_42826# 0.147708f
C2476 a_1823_45246# a_4093_43548# 0.17443f
C2477 a_n1613_43370# a_526_44458# 0.826565f
C2478 a_n237_47217# a_2277_45546# 0.104529f
C2479 a_n443_46116# a_n452_45724# 0.188857f
C2480 a_17061_44734# VDD 0.17647f
C2481 a_3422_30871# EN_VIN_BSTR_N 0.182769f
C2482 a_n2442_46660# a_n4315_30879# 0.361271f
C2483 a_n452_44636# a_n356_44636# 0.318214f
C2484 a_12607_44458# a_12883_44458# 0.11453f
C2485 a_n443_42852# a_9803_43646# 0.102893f
C2486 a_9290_44172# a_10903_43370# 0.340316f
C2487 a_11189_46129# a_11387_46155# 0.320331f
C2488 a_12549_44172# a_18479_45785# 0.105486f
C2489 a_1427_43646# VDD 0.19291f
C2490 a_5385_46902# VDD 0.203316f
C2491 a_n2017_45002# a_743_42282# 7.84646f
C2492 a_n2497_47436# a_n971_45724# 0.229429f
C2493 a_n2109_47186# a_n815_47178# 0.160027f
C2494 a_n1741_47186# SMPL_ON_P 0.178214f
C2495 a_n1533_46116# VDD 0.143145f
C2496 a_n443_42852# a_n913_45002# 0.796158f
C2497 a_12549_44172# a_14021_43940# 0.150377f
C2498 a_19431_45546# VDD 0.342308f
C2499 a_10903_43370# a_10807_43548# 0.193971f
C2500 a_n1613_43370# a_8605_42826# 0.159791f
C2501 a_n237_47217# a_8049_45260# 0.109887f
C2502 a_n881_46662# a_167_45260# 0.108232f
C2503 a_10227_46804# a_15015_46420# 0.287571f
C2504 a_13076_44458# VDD 0.180665f
C2505 a_n863_45724# a_1568_43370# 0.202455f
C2506 a_n2661_45546# a_3080_42308# 0.155045f
C2507 a_1138_42852# a_791_42968# 0.100783f
C2508 a_1423_45028# a_9313_44734# 0.241551f
C2509 a_n2497_47436# a_n2293_45010# 0.233882f
C2510 a_376_46348# a_472_46348# 0.318161f
C2511 a_16388_46812# a_17957_46116# 0.140894f
C2512 a_8270_45546# a_8049_45260# 0.321896f
C2513 a_12891_46348# VDD 1.01428f
C2514 a_7499_43078# a_7871_42858# 0.146369f
C2515 a_8199_44636# a_8685_42308# 0.114007f
C2516 a_n2956_38680# a_n2956_38216# 0.10753f
C2517 a_5937_45572# a_5907_45546# 0.104991f
C2518 a_15959_42545# a_15890_42674# 0.209641f
C2519 a_4520_42826# VDD 0.142755f
C2520 a_n913_45002# a_14635_42282# 0.332583f
C2521 a_5891_43370# a_8685_43396# 0.145735f
C2522 a_21076_30879# VREF 0.417978f
C2523 a_13249_42308# a_13070_42354# 0.141799f
C2524 a_805_46414# VDD 0.154663f
C2525 a_768_44030# a_5244_44056# 0.167173f
C2526 a_15227_44166# a_14539_43914# 0.520312f
C2527 a_8746_45002# a_10490_45724# 0.116339f
C2528 a_5742_30871# VCM 0.211981f
C2529 a_11322_45546# VDD 0.370908f
C2530 a_n2810_45028# a_n3565_38216# 0.349341f
C2531 a_13747_46662# a_13607_46688# 0.168294f
C2532 VDD SINGLE_ENDED 0.210835f
C2533 a_12549_44172# a_19692_46634# 0.491923f
C2534 a_2063_45854# a_5204_45822# 0.174206f
C2535 a_n443_46116# a_167_45260# 0.794635f
C2536 C1_N_btm VIN_N 0.39234f
C2537 a_11599_46634# a_12741_44636# 0.183316f
C2538 C0_N_btm VREF 0.443884f
C2539 a_4651_46660# a_4817_46660# 0.57393f
C2540 C0_dummy_P_btm VCM 0.311452f
C2541 a_9290_44172# a_8685_43396# 0.207262f
C2542 a_20273_46660# a_21188_46660# 0.118759f
C2543 a_8270_45546# a_8953_45546# 1.06716f
C2544 a_7281_43914# VDD 0.198809f
C2545 a_7903_47542# VDD 0.202868f
C2546 a_2107_46812# a_2437_43646# 0.185914f
C2547 a_768_44030# a_5111_44636# 0.154519f
C2548 a_16409_43396# VDD 0.250832f
C2549 a_6761_42308# a_6123_31319# 0.187371f
C2550 a_12359_47026# VDD 0.142103f
C2551 a_4915_47217# a_9313_45822# 0.366722f
C2552 a_6851_47204# a_7227_47204# 0.241208f
C2553 a_6545_47178# a_6575_47204# 0.11927f
C2554 a_1273_38525# a_2112_39137# 0.225378f
C2555 a_564_42282# VDD 0.293756f
C2556 a_n356_44636# a_n2293_42282# 1.10197f
C2557 a_n913_45002# a_19511_42282# 0.120073f
C2558 a_n2810_45572# VDD 0.557886f
C2559 a_18175_45572# a_19256_45572# 0.102355f
C2560 a_18341_45572# a_18691_45572# 0.206455f
C2561 a_8270_45546# a_9028_43914# 0.233359f
C2562 VDAC_N C5_N_btm 27.606901f
C2563 a_n1696_35090# EN_VIN_BSTR_P 0.336639f
C2564 a_n743_46660# a_n2438_43548# 0.426835f
C2565 a_16243_43396# a_16547_43609# 0.165289f
C2566 a_6431_45366# VDD 0.203167f
C2567 a_n237_47217# a_1609_45822# 0.141985f
C2568 a_2905_45572# a_2957_45546# 0.137248f
C2569 a_11599_46634# a_16375_45002# 0.407484f
C2570 a_16241_44734# VDD 0.189894f
C2571 a_3422_30871# a_11530_34132# 0.127528f
C2572 en_comp a_n2661_42282# 0.103098f
C2573 a_n443_42852# a_9145_43396# 2.32123f
C2574 a_11189_46129# a_11133_46155# 0.203074f
C2575 a_11453_44696# a_2437_43646# 0.189184f
C2576 a_n1557_42282# VDD 0.355513f
C2577 a_4817_46660# VDD 0.370615f
C2578 a_n1059_45260# a_4190_30871# 0.133926f
C2579 a_3422_30871# a_20512_43084# 0.125955f
C2580 a_10809_44734# a_11823_42460# 0.215753f
C2581 a_21613_42308# a_22775_42308# 0.225363f
C2582 a_22400_42852# a_22889_38993# 0.13715f
C2583 a_n913_45002# a_4921_42308# 0.169235f
C2584 a_n443_42852# a_n1059_45260# 0.130036f
C2585 a_13661_43548# a_15493_43940# 1.28948f
C2586 a_n971_45724# a_6969_46634# 0.235123f
C2587 a_8530_39574# a_8912_37509# 0.426772f
C2588 a_18691_45572# VDD 0.191893f
C2589 a_10903_43370# a_10949_43914# 0.451961f
C2590 a_3232_43370# a_6171_45002# 0.314056f
C2591 a_4883_46098# a_10355_46116# 0.23167f
C2592 a_11599_46634# a_18985_46122# 0.570252f
C2593 a_10227_46804# a_14275_46494# 0.18614f
C2594 a_13661_43548# a_12741_44636# 0.13948f
C2595 a_12883_44458# VDD 0.263743f
C2596 a_n971_45724# a_3357_43084# 0.565799f
C2597 a_n1925_42282# a_n2104_42282# 0.166917f
C2598 a_11309_47204# VDD 0.358104f
C2599 a_7499_43078# a_7227_42852# 0.126148f
C2600 a_3065_45002# a_3539_42460# 0.300764f
C2601 a_584_46384# a_n356_44636# 0.268036f
C2602 a_5934_30871# a_7174_31319# 0.473128f
C2603 a_472_46348# VDD 0.706547f
C2604 a_20202_43084# a_18494_42460# 0.166633f
C2605 a_526_44458# a_3065_45002# 0.138202f
C2606 a_1823_45246# a_n2661_43370# 0.112095f
C2607 a_9313_45822# a_n881_46662# 1.00227f
C2608 a_15890_42674# VDD 0.203548f
C2609 a_5742_30871# VREF_GND 0.191352f
C2610 a_21177_47436# a_13507_46334# 0.329096f
C2611 a_n1151_42308# a_5807_45002# 1.52318f
C2612 a_6151_47436# a_12549_44172# 0.214024f
C2613 a_6575_47204# a_8128_46384# 0.105633f
C2614 a_n2956_37592# a_n4209_38216# 0.104159f
C2615 a_10490_45724# VDD 0.162001f
C2616 a_n755_45592# a_n699_43396# 0.185444f
C2617 VDD START 0.114358f
C2618 C0_N_btm VIN_N 0.529671f
C2619 C0_P_btm VCM 0.717283f
C2620 a_4651_46660# a_4955_46873# 0.140348f
C2621 a_4646_46812# a_4817_46660# 0.588038f
C2622 a_4361_42308# a_21855_43396# 0.167446f
C2623 a_13467_32519# a_13678_32519# 10.9526f
C2624 a_6171_45002# a_8975_43940# 0.175346f
C2625 a_13059_46348# a_11415_45002# 0.225168f
C2626 a_20841_46902# a_20623_46660# 0.209641f
C2627 a_8270_45546# a_5937_45572# 0.29626f
C2628 a_6453_43914# VDD 0.194953f
C2629 a_7227_47204# VDD 0.430714f
C2630 a_n2661_43370# a_n3674_39768# 0.144159f
C2631 a_768_44030# a_5147_45002# 0.191082f
C2632 a_16547_43609# VDD 0.31275f
C2633 a_6761_42308# a_7227_42308# 0.173849f
C2634 a_5932_42308# a_5934_30871# 1.37963f
C2635 a_11967_42832# a_15493_43940# 0.299734f
C2636 a_5111_44636# a_5111_42852# 0.148196f
C2637 a_11415_45002# a_13556_45296# 0.16025f
C2638 a_3503_45724# a_3775_45552# 0.13675f
C2639 a_4185_45028# a_413_45260# 0.191095f
C2640 a_4915_47217# a_11031_47542# 0.125943f
C2641 a_n4064_39072# a_n2302_39072# 0.250408f
C2642 a_n3674_37592# VDD 0.357168f
C2643 a_3422_30871# a_5649_42852# 0.291966f
C2644 a_n2840_45546# VDD 0.302566f
C2645 a_n2293_45546# a_n2661_43370# 0.131199f
C2646 a_10193_42453# a_6171_45002# 0.411891f
C2647 a_8746_45002# a_3232_43370# 0.439467f
C2648 a_18341_45572# a_18909_45814# 0.170692f
C2649 VDAC_N C4_N_btm 13.8047f
C2650 a_n1696_35090# a_n1057_35174# 0.419261f
C2651 a_n1550_35608# EN_VIN_BSTR_P 0.573047f
C2652 a_12861_44030# a_3090_45724# 0.496275f
C2653 a_16137_43396# a_16547_43609# 0.151161f
C2654 a_6171_45002# VDD 0.441339f
C2655 a_19479_31679# a_19721_31679# 9.039419f
C2656 a_14673_44172# VDD 0.381917f
C2657 a_16795_42852# a_17333_42852# 0.108694f
C2658 a_13059_46348# a_13259_45724# 0.812126f
C2659 a_10227_46804# a_n913_45002# 0.344574f
C2660 a_12465_44636# a_3357_43084# 1.30897f
C2661 a_n784_42308# a_n3674_37592# 0.254719f
C2662 a_4955_46873# VDD 0.467566f
C2663 a_n1920_47178# a_n1741_47186# 0.173125f
C2664 a_n443_46116# a_2982_43646# 0.140614f
C2665 a_n971_45724# a_6755_46942# 0.185154f
C2666 a_7754_38470# a_8912_37509# 0.575911f
C2667 a_n4064_39616# VREF_GND 0.241027f
C2668 a_n2302_39072# VDD 0.355374f
C2669 a_18909_45814# VDD 0.205795f
C2670 a_5111_44636# a_5205_44484# 0.200189f
C2671 a_n913_45002# a_1307_43914# 0.298747f
C2672 a_11599_46634# a_18819_46122# 0.314824f
C2673 a_10227_46804# a_14493_46090# 0.202633f
C2674 a_n881_46662# a_1823_45246# 0.155149f
C2675 a_12607_44458# VDD 0.188171f
C2676 a_n2497_47436# a_n2661_45010# 0.281004f
C2677 a_16327_47482# a_16680_45572# 0.223571f
C2678 a_768_44030# a_7499_43078# 0.101779f
C2679 a_3065_45002# a_3626_43646# 0.480498f
C2680 a_15803_42450# a_15959_42545# 0.110532f
C2681 a_15764_42576# a_15890_42674# 0.181217f
C2682 a_3681_42891# VDD 0.223661f
C2683 a_2711_45572# a_20107_42308# 0.164316f
C2684 a_376_46348# VDD 0.116284f
C2685 a_20202_43084# a_18184_42460# 0.299795f
C2686 a_526_44458# a_2680_45002# 0.119733f
C2687 a_768_44030# a_3600_43914# 0.182408f
C2688 a_10193_42453# a_8746_45002# 0.11003f
C2689 a_11031_47542# a_n881_46662# 0.183988f
C2690 a_15959_42545# VDD 0.19373f
C2691 a_6151_47436# a_12891_46348# 0.169139f
C2692 a_7903_47542# a_8128_46384# 0.109077f
C2693 a_8746_45002# VDD 0.970181f
C2694 VDD RST_Z 4.72787f
C2695 a_3160_47472# a_3699_46348# 0.109505f
C2696 C0_dummy_N_btm VIN_N 0.544204f
C2697 C1_P_btm VCM 0.716121f
C2698 C0_P_btm VREF_GND 0.350485f
C2699 a_n443_46116# a_1823_45246# 0.217935f
C2700 a_7499_43078# a_7845_44172# 0.112307f
C2701 a_3232_43370# a_8975_43940# 0.620589f
C2702 a_20273_46660# a_20623_46660# 0.20669f
C2703 a_20107_46660# a_21188_46660# 0.102355f
C2704 a_8270_45546# a_8199_44636# 0.95539f
C2705 a_5649_42852# a_5932_42308# 0.126438f
C2706 a_17333_42852# a_18504_43218# 0.157683f
C2707 a_5663_43940# VDD 0.133666f
C2708 a_6851_47204# VDD 0.287724f
C2709 a_9290_44172# a_10586_45546# 0.264957f
C2710 a_16243_43396# VDD 0.39865f
C2711 a_13259_45724# a_17303_42282# 0.460497f
C2712 a_18579_44172# a_18451_43940# 0.147572f
C2713 a_5495_43940# a_5663_43940# 0.227135f
C2714 a_11415_45002# a_9482_43914# 0.309633f
C2715 a_1823_45246# a_3537_45260# 0.482502f
C2716 a_n327_42558# VDD 0.198414f
C2717 a_6491_46660# a_6851_47204# 0.132946f
C2718 a_3422_30871# a_13678_32519# 0.452533f
C2719 a_18175_45572# a_18691_45572# 0.105995f
C2720 a_n237_47217# a_765_45546# 0.1364f
C2721 a_n1021_46688# a_n743_46660# 0.11001f
C2722 a_n1925_46634# a_n2438_43548# 0.166008f
C2723 VDAC_N C3_N_btm 6.907279f
C2724 a_n1550_35608# a_n1057_35174# 0.201872f
C2725 a_16137_43396# a_16243_43396# 0.182209f
C2726 a_3232_43370# VDD 2.96597f
C2727 a_19479_31679# a_18114_32519# 0.182316f
C2728 a_15009_46634# a_14180_46812# 0.123843f
C2729 a_n746_45260# a_n443_42852# 0.136813f
C2730 a_3422_30871# EN_VIN_BSTR_P 0.182769f
C2731 a_17595_43084# a_17701_42308# 0.141211f
C2732 SMPL_ON_P a_n2002_35608# 0.399535f
C2733 a_n746_45260# a_375_42282# 0.41439f
C2734 a_9290_44172# a_11189_46129# 0.199578f
C2735 a_6755_46942# a_2711_45572# 0.612305f
C2736 a_4905_42826# VDD 0.439034f
C2737 a_196_42282# a_n3674_37592# 0.1528f
C2738 a_14537_43396# a_14358_43442# 0.1418f
C2739 a_4651_46660# VDD 0.457722f
C2740 a_8049_45260# a_2711_45572# 2.31131f
C2741 a_n3674_37592# a_n4064_37440# 0.651412f
C2742 a_n2109_47186# a_n1741_47186# 0.18579f
C2743 a_13259_45724# a_9482_43914# 0.321549f
C2744 a_15227_44166# a_17517_44484# 0.104904f
C2745 a_13661_43548# a_11341_43940# 0.15891f
C2746 a_19321_45002# a_20623_43914# 0.294126f
C2747 a_3754_38470# VDAC_P 0.323951f
C2748 a_7754_38470# VDAC_N 0.110605f
C2749 a_8530_39574# a_6886_37412# 0.616015f
C2750 a_n4064_39072# VDD 1.74897f
C2751 a_22959_47212# a_22612_30879# 0.156518f
C2752 a_18341_45572# VDD 0.2432f
C2753 a_n1613_43370# a_7871_42858# 0.659491f
C2754 a_5691_45260# a_3232_43370# 0.123939f
C2755 a_n881_46662# a_1138_42852# 0.148785f
C2756 a_10227_46804# a_13925_46122# 0.635045f
C2757 a_8975_43940# VDD 0.257588f
C2758 a_n863_45724# a_458_43396# 0.122956f
C2759 a_n2661_45546# a_4093_43548# 0.343267f
C2760 a_9290_44172# a_4361_42308# 0.1126f
C2761 a_3090_45724# a_n1925_42282# 0.157861f
C2762 a_16327_47482# a_16855_45546# 0.305145f
C2763 a_n2293_46098# a_1823_45246# 0.107882f
C2764 a_2382_45260# a_3539_42460# 0.110439f
C2765 a_n2956_38680# a_n2810_45572# 5.73878f
C2766 a_4646_46812# a_3232_43370# 0.305673f
C2767 a_n3674_38680# a_n3565_38502# 0.128677f
C2768 a_6123_31319# a_7174_31319# 13.9919f
C2769 a_15764_42576# a_15959_42545# 0.21686f
C2770 a_2905_42968# VDD 0.142081f
C2771 a_20193_45348# a_13887_32519# 0.277027f
C2772 a_20820_30879# VREF 0.195875f
C2773 a_10949_43914# a_12429_44172# 0.156922f
C2774 a_n1076_46494# VDD 0.294742f
C2775 a_16327_47482# a_19862_44208# 0.209324f
C2776 a_2324_44458# a_14537_43396# 0.341957f
C2777 a_768_44030# a_2998_44172# 0.571981f
C2778 a_10180_45724# a_8746_45002# 0.304016f
C2779 a_15803_42450# VDD 0.448709f
C2780 a_20990_47178# a_21177_47436# 0.159555f
C2781 a_4915_47217# a_768_44030# 0.187438f
C2782 a_9863_47436# a_n881_46662# 0.164043f
C2783 a_10193_42453# VDD 2.18892f
C2784 a_15903_45785# a_16019_45002# 0.139976f
C2785 a_3160_47472# a_3483_46348# 0.154179f
C2786 a_4646_46812# a_4651_46660# 0.844575f
C2787 a_12549_44172# a_15227_44166# 0.354423f
C2788 C2_P_btm VCM 0.716172f
C2789 C1_P_btm VREF_GND 0.673422f
C2790 C0_P_btm VREF 0.443926f
C2791 a_13467_32519# a_4361_42308# 0.121732f
C2792 a_20273_46660# a_20841_46902# 0.17072f
C2793 a_5495_43940# VDD 0.173477f
C2794 a_6491_46660# VDD 0.436756f
C2795 a_10193_42453# a_16137_43396# 0.329316f
C2796 a_n755_45592# a_n13_43084# 0.113444f
C2797 a_5932_42308# a_6123_31319# 1.49414f
C2798 a_16137_43396# VDD 0.483673f
C2799 a_3090_45724# a_16922_45042# 0.206138f
C2800 a_1666_39587# a_2112_39137# 0.269764f
C2801 a_n784_42308# VDD 0.59759f
C2802 a_6545_47178# a_6851_47204# 0.134581f
C2803 a_16375_45002# a_17719_45144# 0.201099f
C2804 a_n357_42282# a_n2293_42834# 4.06139f
C2805 a_18479_45785# a_18341_45572# 0.21997f
C2806 a_9290_44172# a_5891_43370# 0.302383f
C2807 a_n1925_46634# a_n743_46660# 0.193773f
C2808 VDAC_N C2_N_btm 3.46253f
C2809 a_n2302_37690# VDD 0.350131f
C2810 a_n1613_43370# a_5732_46660# 0.268372f
C2811 a_5691_45260# VDD 0.205518f
C2812 a_2905_45572# a_n755_45592# 0.168143f
C2813 a_14084_46812# a_14180_46812# 0.318161f
C2814 a_n971_45724# a_n443_42852# 0.329303f
C2815 a_11599_46634# a_13259_45724# 0.249721f
C2816 a_3080_42308# VDD 0.849776f
C2817 a_20193_45348# a_14401_32519# 0.175398f
C2818 a_4646_46812# VDD 2.53408f
C2819 a_21335_42336# a_21613_42308# 0.110671f
C2820 a_n2497_47436# SMPL_ON_P 0.131317f
C2821 a_2063_45854# a_7715_46873# 0.178294f
C2822 a_7754_38470# a_6886_37412# 0.181496f
C2823 a_3754_38470# a_8912_37509# 1.88278f
C2824 a_n3420_39616# VREF_GND 0.117023f
C2825 a_8530_39574# a_5700_37509# 0.947638f
C2826 a_n2946_39072# VDD 0.383374f
C2827 a_18479_45785# VDD 0.536075f
C2828 a_20974_43370# a_4190_30871# 0.214288f
C2829 a_9290_44172# a_10807_43548# 0.364112f
C2830 a_13661_43548# a_11415_45002# 0.107787f
C2831 a_13747_46662# a_20202_43084# 0.308003f
C2832 a_4883_46098# a_9625_46129# 0.164961f
C2833 a_11599_46634# a_18189_46348# 0.101491f
C2834 a_10227_46804# a_13759_46122# 0.920747f
C2835 a_3080_42308# a_n784_42308# 0.170007f
C2836 a_10057_43914# VDD 0.399284f
C2837 a_n901_46420# a_n1076_46494# 0.234322f
C2838 a_16327_47482# a_16115_45572# 0.163022f
C2839 a_n971_45724# a_2437_43646# 0.204278f
C2840 a_14021_43940# VDD 1.60583f
C2841 a_9804_47204# VDD 0.410522f
C2842 a_n1059_45260# a_8791_43396# 0.196029f
C2843 a_8953_45546# a_5934_30871# 0.113715f
C2844 a_n2438_43548# a_1423_45028# 0.242599f
C2845 a_12465_44636# a_11691_44458# 0.15589f
C2846 a_11453_44696# a_11827_44484# 0.170003f
C2847 a_15764_42576# a_15803_42450# 0.901878f
C2848 a_21076_30879# EN_OFFSET_CAL 0.2809f
C2849 a_11967_42832# a_n97_42460# 0.489711f
C2850 a_n901_46420# VDD 0.518805f
C2851 a_12861_44030# a_15493_43940# 0.370814f
C2852 a_10180_45724# a_10193_42453# 0.145672f
C2853 a_15764_42576# VDD 0.258303f
C2854 a_n443_46116# a_768_44030# 0.177051f
C2855 a_n971_45724# a_n2661_46634# 0.190714f
C2856 a_4915_47217# a_12549_44172# 0.316329f
C2857 a_n2497_47436# a_n2438_43548# 0.206216f
C2858 a_22485_38105# a_22629_38406# 0.206945f
C2859 a_3905_42865# a_3935_42891# 0.240349f
C2860 en_comp a_1107_38525# 0.206093f
C2861 a_10180_45724# VDD 0.336512f
C2862 a_n2293_46634# a_8685_43396# 0.335608f
C2863 a_5257_43370# a_n97_42460# 0.167676f
C2864 a_22959_45572# a_20447_31679# 0.154273f
C2865 a_12861_44030# a_12741_44636# 0.366155f
C2866 a_n971_45724# a_8199_44636# 0.247183f
C2867 a_3160_47472# a_3147_46376# 0.208295f
C2868 C0_dummy_P_btm VIN_P 0.544204f
C2869 C3_P_btm VCM 0.716273f
C2870 C2_P_btm VREF_GND 0.671742f
C2871 C1_P_btm VREF 0.98698f
C2872 a_13661_43548# a_13259_45724# 0.250875f
C2873 a_20107_46660# a_20623_46660# 0.105914f
C2874 a_5013_44260# VDD 0.198233f
C2875 a_20193_45348# a_20512_43084# 0.160912f
C2876 a_6545_47178# VDD 0.386368f
C2877 a_n357_42282# a_n13_43084# 0.194173f
C2878 a_10903_43370# a_8049_45260# 0.114138f
C2879 a_768_44030# a_3537_45260# 0.341201f
C2880 a_4185_45028# a_13259_45724# 0.194989f
C2881 a_19692_46634# VDD 2.53528f
C2882 a_19279_43940# a_19328_44172# 0.120319f
C2883 a_5013_44260# a_5495_43940# 0.251039f
C2884 a_11415_45002# a_13159_45002# 0.141106f
C2885 a_1823_45246# a_3065_45002# 0.607468f
C2886 a_1273_38525# a_1666_39043# 0.297741f
C2887 a_196_42282# VDD 0.291844f
C2888 a_n3420_39072# a_n4064_39072# 4.91095f
C2889 a_2063_45854# a_11599_46634# 0.19861f
C2890 a_4915_47217# a_6575_47204# 0.849579f
C2891 a_6545_47178# a_6491_46660# 0.181574f
C2892 a_18184_42460# a_22400_42852# 0.16156f
C2893 a_20692_30879# VDD 0.499669f
C2894 a_n2661_45546# a_n2661_43370# 0.145941f
C2895 a_18175_45572# a_18341_45572# 0.577068f
C2896 a_n971_45724# a_765_45546# 0.140618f
C2897 VDAC_N C1_N_btm 1.7375f
C2898 a_n4064_37440# VDD 1.65981f
C2899 a_n1613_43370# a_5907_46634# 0.338694f
C2900 a_4927_45028# VDD 0.159822f
C2901 a_14401_32519# a_5534_30871# 0.339008f
C2902 a_4883_46098# a_8049_45260# 0.469963f
C2903 a_12549_44172# a_10809_44734# 2.27272f
C2904 a_n743_46660# a_9823_46155# 0.196587f
C2905 a_12465_44636# a_2437_43646# 0.18195f
C2906 COMP_P a_n1794_35242# 2.45645f
C2907 a_n473_42460# a_n327_42558# 0.171361f
C2908 a_4699_43561# VDD 0.262218f
C2909 a_3877_44458# VDD 0.786903f
C2910 a_22400_42852# a_22527_39145# 0.228292f
C2911 a_14955_43940# a_15037_43940# 0.171361f
C2912 a_15227_44166# a_16241_44734# 0.105126f
C2913 a_n863_45724# a_2382_45260# 0.119625f
C2914 a_3754_38470# VDAC_N 0.169096f
C2915 a_8530_39574# a_5088_37509# 0.166912f
C2916 a_7754_38470# a_5700_37509# 0.971846f
C2917 a_n881_46662# a_12549_44172# 0.225257f
C2918 a_n4064_37440# a_n2302_37690# 0.239588f
C2919 SMPL_ON_N a_22612_30879# 5.16049f
C2920 a_n3420_39072# VDD 1.01442f
C2921 a_18175_45572# VDD 0.38478f
C2922 a_14401_32519# a_4190_30871# 0.10855f
C2923 a_9290_44172# a_10949_43914# 0.113864f
C2924 a_13259_45724# a_11967_42832# 0.141918f
C2925 a_5111_44636# a_3232_43370# 0.134191f
C2926 a_10440_44484# VDD 0.159539f
C2927 a_22959_45036# a_19721_31679# 0.156264f
C2928 a_n755_45592# a_n97_42460# 1.02989f
C2929 a_16327_47482# a_16333_45814# 0.168559f
C2930 a_10341_42308# a_9803_42558# 0.108853f
C2931 a_8128_46384# VDD 0.403575f
C2932 a_5111_44636# a_4905_42826# 0.128918f
C2933 a_5883_43914# a_7542_44172# 0.187537f
C2934 a_1847_42826# VDD 0.527555f
C2935 a_15486_42560# a_15803_42450# 0.102355f
C2936 a_10729_43914# a_11750_44172# 0.144893f
C2937 a_2711_45572# a_19511_42282# 0.234026f
C2938 a_n1641_46494# VDD 0.226065f
C2939 a_15486_42560# VDD 0.275297f
C2940 a_20894_47436# a_20990_47178# 0.313533f
C2941 a_4915_47217# a_12891_46348# 0.156543f
C2942 a_6575_47204# a_n881_46662# 0.708623f
C2943 a_3905_42865# a_3681_42891# 0.101054f
C2944 a_4699_43561# a_3080_42308# 0.223965f
C2945 a_10053_45546# VDD 0.150582f
C2946 a_19692_46634# a_14021_43940# 0.775991f
C2947 C0_P_btm VIN_P 0.529671f
C2948 C10_N_btm VDD 2.40001f
C2949 a_12549_44172# a_17609_46634# 0.487224f
C2950 C3_P_btm VREF_GND 0.67174f
C2951 C4_P_btm VCM 0.716447f
C2952 C2_P_btm VREF 0.987884f
C2953 a_20411_46873# a_20273_46660# 0.219954f
C2954 a_5244_44056# VDD 0.146618f
C2955 a_4007_47204# DATA[2] 0.337596f
C2956 a_6151_47436# VDD 4.39915f
C2957 w_11334_34010# a_3422_30871# 1.91172f
C2958 a_5244_44056# a_5495_43940# 0.107037f
C2959 a_19466_46812# VDD 0.664497f
C2960 a_n913_45002# a_12545_42858# 0.548984f
C2961 a_3537_45260# a_5111_42852# 0.123919f
C2962 a_11415_45002# a_13017_45260# 0.100288f
C2963 a_n473_42460# VDD 0.27195f
C2964 a_n3420_39072# a_n2946_39072# 0.238708f
C2965 a_6151_47436# a_6491_46660# 0.31912f
C2966 a_3422_30871# a_13467_32519# 0.421402f
C2967 a_20205_31679# VDD 0.737408f
C2968 a_9049_44484# a_3232_43370# 0.17048f
C2969 a_526_44458# a_n699_43396# 0.285f
C2970 a_13259_45724# a_18315_45260# 0.144632f
C2971 a_18175_45572# a_18479_45785# 0.280208f
C2972 a_n2293_46634# a_n2438_43548# 0.807205f
C2973 VDAC_N C0_N_btm 0.901121f
C2974 VDAC_P C0_dummy_P_btm 0.88451f
C2975 a_n2002_35608# a_n1550_35608# 0.150805f
C2976 a_n2946_37690# VDD 0.38221f
C2977 a_n1151_42308# a_13885_46660# 0.333314f
C2978 a_n1613_43370# a_5167_46660# 0.177362f
C2979 a_5111_44636# VDD 1.28013f
C2980 a_12891_46348# a_10809_44734# 0.102888f
C2981 a_n443_46116# a_n2661_45546# 0.136593f
C2982 a_14084_46812# a_13885_46660# 0.237373f
C2983 a_n743_46660# a_9569_46155# 0.104962f
C2984 a_10903_43370# a_5534_30871# 0.134296f
C2985 a_13717_47436# a_413_45260# 4.36729f
C2986 a_n4318_37592# a_n1794_35242# 0.847279f
C2987 a_n4318_38680# a_n4209_38502# 0.105064f
C2988 a_4235_43370# VDD 0.229422f
C2989 a_n1059_45260# a_16823_43084# 0.318918f
C2990 a_3422_30871# a_22315_44484# 0.19914f
C2991 a_10227_46804# a_9313_44734# 0.875947f
C2992 a_10809_44734# a_11322_45546# 0.22629f
C2993 a_22400_42852# a_22589_40055# 0.663766f
C2994 a_n2288_47178# a_n2109_47186# 0.177673f
C2995 a_n2956_38680# VDD 0.871805f
C2996 a_n913_45002# a_5379_42460# 0.179494f
C2997 a_3905_42865# a_4905_42826# 0.404829f
C2998 a_310_45028# a_n37_45144# 0.112458f
C2999 a_n2661_45546# a_3537_45260# 0.780422f
C3000 a_10193_42453# a_16147_45260# 0.193225f
C3001 a_15227_44166# a_14673_44172# 0.357896f
C3002 a_18189_46348# a_18315_45260# 0.101775f
C3003 a_n755_45592# a_n467_45028# 0.26002f
C3004 a_n863_45724# a_2274_45254# 0.17549f
C3005 a_6151_47436# a_4646_46812# 0.153739f
C3006 a_2063_45854# a_5257_43370# 0.426517f
C3007 a_7754_38470# a_5088_37509# 0.394117f
C3008 SMPL_ON_N a_21588_30879# 0.119129f
C3009 a_n3690_39392# VDD 0.363068f
C3010 en_comp a_22527_39145# 0.393507f
C3011 a_16147_45260# VDD 0.197706f
C3012 a_5111_44636# a_5691_45260# 0.130044f
C3013 a_5147_45002# a_3232_43370# 0.253159f
C3014 a_10334_44484# VDD 0.19332f
C3015 a_5649_42852# a_5534_30871# 0.234793f
C3016 a_1847_42826# a_2075_43172# 0.103349f
C3017 a_n1557_42282# COMP_P 0.123881f
C3018 a_n357_42282# a_n97_42460# 0.900712f
C3019 a_1423_45028# a_5891_43370# 0.301629f
C3020 a_2382_45260# a_2982_43646# 0.468592f
C3021 a_8199_44636# a_5934_30871# 0.159294f
C3022 a_10903_43370# a_n443_42852# 0.176275f
C3023 a_791_42968# VDD 0.128737f
C3024 a_15486_42560# a_15764_42576# 0.118759f
C3025 a_n1423_46090# VDD 0.227012f
C3026 a_10729_43914# a_10807_43548# 0.238591f
C3027 a_2127_44172# a_2253_43940# 0.143754f
C3028 a_12741_44636# EN_OFFSET_CAL 0.230064f
C3029 a_7499_43078# a_8746_45002# 0.153858f
C3030 a_12741_44636# a_16922_45042# 0.139755f
C3031 a_10053_45546# a_10180_45724# 0.144403f
C3032 a_7903_47542# a_n881_46662# 0.178742f
C3033 a_15051_42282# VDD 0.461307f
C3034 a_9049_44484# VDD 0.680993f
C3035 a_15493_43940# a_15743_43084# 0.206331f
C3036 a_2437_43646# a_n2661_45010# 0.15182f
C3037 C1_P_btm VIN_P 0.39234f
C3038 C9_N_btm VDD 0.345685f
C3039 C4_P_btm VREF_GND 0.671882f
C3040 C5_P_btm VCM 0.719982f
C3041 C3_P_btm VREF 0.984942f
C3042 a_4190_30871# a_5649_42852# 0.434284f
C3043 a_21487_43396# a_13467_32519# 0.152042f
C3044 a_20107_46660# a_20273_46660# 0.608339f
C3045 a_10227_46804# a_2711_45572# 0.130695f
C3046 a_3905_42865# VDD 0.788273f
C3047 a_5815_47464# VDD 0.399354f
C3048 a_n2293_46098# a_n2661_45546# 3.03243f
C3049 a_n881_46662# a_6431_45366# 0.177591f
C3050 a_768_44030# a_3065_45002# 0.288972f
C3051 a_n1613_43370# a_5205_44484# 0.551795f
C3052 a_3483_46348# a_13259_45724# 0.230226f
C3053 a_1606_42308# a_5742_30871# 3.46204f
C3054 a_19333_46634# VDD 0.199048f
C3055 a_1823_45246# a_2382_45260# 0.801932f
C3056 a_n961_42308# VDD 0.24416f
C3057 a_n3565_39304# a_n4064_39072# 0.344587f
C3058 a_6151_47436# a_6545_47178# 0.39775f
C3059 a_2711_45572# a_1307_43914# 0.187968f
C3060 a_7499_43078# a_3232_43370# 0.318423f
C3061 a_16375_45002# a_16922_45042# 0.170835f
C3062 a_11599_46634# a_11813_46116# 0.106062f
C3063 VDAC_N C0_dummy_N_btm 0.885361f
C3064 VDAC_P C0_P_btm 0.901219f
C3065 a_n3420_37440# VDD 2.26579f
C3066 a_n1613_43370# a_5385_46902# 0.182522f
C3067 a_5147_45002# VDD 0.574918f
C3068 a_413_45260# EN_OFFSET_CAL 0.114452f
C3069 a_6171_45002# a_n2661_43370# 2.37006f
C3070 a_n863_45724# a_1414_42308# 0.711805f
C3071 a_13059_46348# a_14579_43548# 0.171744f
C3072 a_n755_45592# a_n809_44244# 0.404418f
C3073 a_2711_45572# a_18579_44172# 0.170319f
C3074 a_13607_46688# a_13885_46660# 0.11044f
C3075 a_n743_46660# a_9625_46129# 0.206271f
C3076 a_n2661_46634# a_10903_43370# 0.663878f
C3077 a_n443_42852# a_8685_43396# 0.281116f
C3078 a_16327_47482# a_n913_45002# 0.137194f
C3079 a_4883_46098# a_2437_43646# 0.458866f
C3080 a_n961_42308# a_n784_42308# 0.154417f
C3081 a_4093_43548# VDD 0.216874f
C3082 a_5891_43370# a_10405_44172# 0.15894f
C3083 a_n3674_37592# a_n3565_37414# 0.129086f
C3084 a_n784_42308# a_n3420_37440# 0.140549f
C3085 a_n2497_47436# a_n2109_47186# 0.197671f
C3086 a_13483_43940# a_13565_43940# 0.171361f
C3087 a_n2956_39304# VDD 0.455981f
C3088 a_n863_45724# a_1667_45002# 0.20954f
C3089 a_526_44458# a_n2293_42834# 1.7774f
C3090 a_n4209_39590# VCM 0.179761f
C3091 a_3754_38470# a_5700_37509# 0.124176f
C3092 a_7754_38470# a_4338_37500# 0.208561f
C3093 a_8530_39574# a_3726_37500# 1.35509f
C3094 a_n3565_39304# VDD 0.888861f
C3095 a_n3565_39590# VREF 0.417978f
C3096 en_comp a_22589_40055# 0.260977f
C3097 a_n97_42460# a_19700_43370# 0.154491f
C3098 a_5111_44636# a_4927_45028# 0.134309f
C3099 a_7499_43078# a_8975_43940# 0.519621f
C3100 a_4883_46098# a_8199_44636# 0.242f
C3101 a_11599_46634# a_15682_46116# 1.8289f
C3102 a_10157_44484# VDD 0.174233f
C3103 a_22223_45036# a_18114_32519# 0.15655f
C3104 a_n1991_46122# a_n1076_46494# 0.124988f
C3105 a_19778_44110# a_19862_44208# 0.213467f
C3106 a_n755_45592# a_n2293_42282# 0.208531f
C3107 a_13507_46334# a_20193_45348# 0.253904f
C3108 a_14113_42308# a_15803_42450# 0.289859f
C3109 a_20820_30879# EN_OFFSET_CAL 0.107181f
C3110 a_n1991_46122# VDD 0.581018f
C3111 a_10729_43914# a_10949_43914# 0.418928f
C3112 a_10809_44734# a_6171_45002# 0.244599f
C3113 a_7499_43078# a_10193_42453# 0.298293f
C3114 a_526_44458# a_413_45260# 0.103799f
C3115 a_14113_42308# VDD 0.365578f
C3116 a_7499_43078# VDD 1.87959f
C3117 a_1049_43396# a_n1557_42282# 0.211757f
C3118 a_n863_45724# a_n699_43396# 0.23135f
C3119 C2_P_btm VIN_P 0.502408f
C3120 C8_N_btm VDD 0.19922f
C3121 a_2063_45854# a_3483_46348# 0.164542f
C3122 C5_P_btm VREF_GND 0.676559f
C3123 C6_P_btm VCM 0.877162f
C3124 C4_P_btm VREF 0.98728f
C3125 a_3422_30871# a_7174_31319# 2.22059f
C3126 a_743_42282# a_4361_42308# 7.66647f
C3127 a_n913_45002# a_n356_44636# 0.640597f
C3128 a_20107_46660# a_20411_46873# 0.316529f
C3129 a_n743_46660# a_8049_45260# 2.07544f
C3130 a_3600_43914# VDD 0.22716f
C3131 a_5649_42852# a_4921_42308# 0.133152f
C3132 a_3785_47178# DATA[2] 0.119025f
C3133 a_5129_47502# VDD 0.20906f
C3134 a_10903_43370# a_13291_42460# 0.135558f
C3135 a_4185_45028# a_22400_42852# 0.105559f
C3136 a_15227_44166# a_10193_42453# 0.205591f
C3137 a_15781_43660# VDD 0.196099f
C3138 a_n2956_39304# a_n2946_39072# 0.150476f
C3139 a_3905_42865# a_5013_44260# 0.182997f
C3140 a_15227_44166# VDD 2.69945f
C3141 a_167_45260# a_327_44734# 0.199136f
C3142 a_n2293_46634# a_5891_43370# 0.105307f
C3143 a_n755_45592# a_3775_45552# 0.100709f
C3144 a_13259_45724# a_13249_42308# 0.358931f
C3145 a_1823_45246# a_2274_45254# 0.255985f
C3146 a_1666_39587# a_1666_39043# 1.95282f
C3147 a_n4334_39392# a_n4064_39072# 0.410653f
C3148 a_n4209_39304# a_n2302_39072# 0.407162f
C3149 a_n3690_39392# a_n3420_39072# 0.414961f
C3150 a_n3565_39304# a_n2946_39072# 0.410957f
C3151 a_n1329_42308# VDD 0.237697f
C3152 a_4915_47217# a_6851_47204# 0.172567f
C3153 a_16147_45260# a_18175_45572# 0.108647f
C3154 a_11599_46634# a_11735_46660# 0.268769f
C3155 a_n2104_46634# a_n1925_46634# 0.167849f
C3156 VDAC_P C1_P_btm 1.74268f
C3157 a_n3690_37440# VDD 0.363068f
C3158 a_n1613_43370# a_4817_46660# 0.330391f
C3159 a_4558_45348# VDD 0.25277f
C3160 a_12861_44030# a_13259_45724# 0.435853f
C3161 a_n2293_46634# a_9290_44172# 0.102393f
C3162 a_3626_43646# a_5742_30871# 0.168508f
C3163 a_5147_45002# a_5013_44260# 0.189328f
C3164 a_10334_44484# a_10440_44484# 0.313533f
C3165 a_4646_46812# a_7499_43078# 0.158236f
C3166 a_16327_47482# a_n1059_45260# 0.235708f
C3167 a_n4318_37592# a_n3674_37592# 3.06402f
C3168 a_n3674_38216# a_n1794_35242# 0.333493f
C3169 a_1756_43548# VDD 0.138878f
C3170 a_14537_43396# a_9145_43396# 0.129182f
C3171 a_22400_42852# a_22537_40625# 0.93502f
C3172 a_22959_46124# VDD 0.309939f
C3173 a_13747_46662# a_19862_44208# 0.15289f
C3174 a_n863_45724# a_327_44734# 0.353745f
C3175 a_n971_45724# a_8147_43396# 0.116186f
C3176 VDAC_Ni a_6886_37412# 0.178275f
C3177 a_n4334_39392# VDD 0.385989f
C3178 a_n443_46116# a_4955_46873# 0.126551f
C3179 a_3754_38470# a_5088_37509# 0.632585f
C3180 a_7754_38470# a_3726_37500# 0.124796f
C3181 a_n3420_37440# a_n4064_37440# 8.19012f
C3182 a_22223_47212# a_21588_30879# 0.164932f
C3183 a_20193_45348# a_21613_42308# 0.137559f
C3184 a_5147_45002# a_4927_45028# 0.168157f
C3185 a_7499_43078# a_10057_43914# 0.262644f
C3186 a_n357_42282# a_n2661_42834# 0.239713f
C3187 a_2905_45572# a_526_44458# 0.142766f
C3188 a_11599_46634# a_2324_44458# 0.428445f
C3189 a_9838_44484# VDD 0.242131f
C3190 a_n1557_42282# a_n1736_42282# 0.170341f
C3191 a_9290_44172# a_743_42282# 0.117511f
C3192 a_1423_45028# a_7640_43914# 0.105665f
C3193 a_16327_47482# a_15599_45572# 0.331892f
C3194 a_n1423_46090# a_n1641_46494# 0.209641f
C3195 a_n2109_47186# a_3357_43084# 0.170493f
C3196 a_5883_43914# a_5663_43940# 0.153361f
C3197 a_n881_46662# RST_Z 0.351994f
C3198 a_12465_44636# a_11827_44484# 0.785011f
C3199 a_15051_42282# a_15486_42560# 0.234322f
C3200 a_14113_42308# a_15764_42576# 0.229529f
C3201 a_5932_42308# a_7174_31319# 13.0265f
C3202 a_n1853_46287# VDD 0.645231f
C3203 a_11823_42460# a_11551_42558# 0.138126f
C3204 a_10809_44734# a_3232_43370# 0.158726f
C3205 a_13657_42558# VDD 0.195727f
C3206 a_10227_46804# a_4883_46098# 0.200137f
C3207 a_22485_38105# a_22537_39537# 0.559814f
C3208 a_1209_43370# a_n1557_42282# 0.113851f
C3209 a_8568_45546# VDD 0.182812f
C3210 a_22591_45572# a_19963_31679# 0.161955f
C3211 a_13507_46334# a_4190_30871# 0.186424f
C3212 a_n1925_42282# a_n2293_43922# 2.06056f
C3213 C7_P_btm VCM 1.58335f
C3214 C6_P_btm VREF_GND 0.836236f
C3215 C3_P_btm VIN_P 0.455045f
C3216 C9_N_btm C10_N_btm 53.3168f
C3217 C7_N_btm VDD 0.121904f
C3218 a_10227_46804# a_21188_46660# 0.22222f
C3219 C5_P_btm VREF 0.987144f
C3220 a_n2661_43370# VDD 1.53673f
C3221 a_7229_43940# a_5343_44458# 0.196399f
C3222 a_3232_43370# a_5883_43914# 0.337937f
C3223 a_2998_44172# VDD 0.362233f
C3224 a_4915_47217# VDD 3.43172f
C3225 a_15681_43442# VDD 0.159054f
C3226 a_n2956_39304# a_n3420_39072# 0.208204f
C3227 a_18834_46812# VDD 0.116625f
C3228 a_167_45260# a_413_45260# 0.120357f
C3229 a_1823_45246# a_1667_45002# 0.24808f
C3230 a_n4209_39304# a_n4064_39072# 0.19711f
C3231 a_n3565_39304# a_n3420_39072# 0.241179f
C3232 COMP_P VDD 3.52703f
C3233 a_4915_47217# a_6491_46660# 0.19739f
C3234 a_5815_47464# a_6151_47436# 0.235454f
C3235 a_n1059_45260# a_18727_42674# 0.20226f
C3236 a_4883_46098# a_9396_43370# 0.172323f
C3237 a_10227_46804# a_8685_43396# 0.227547f
C3238 a_n863_45724# a_n2293_42834# 0.107229f
C3239 a_10809_44734# a_8975_43940# 0.169586f
C3240 a_8953_45546# a_5891_43370# 0.321625f
C3241 a_n2661_46634# a_n2438_43548# 0.493975f
C3242 a_n2104_46634# a_n2312_38680# 0.154937f
C3243 VDAC_P C2_P_btm 3.46245f
C3244 a_n3565_37414# VDD 0.783444f
C3245 a_1414_42308# a_1184_42692# 0.115223f
C3246 a_4574_45260# VDD 0.122256f
C3247 a_10341_43396# a_15743_43084# 0.464206f
C3248 a_13661_43548# a_2324_44458# 0.307974f
C3249 a_584_46384# a_n357_42282# 0.107436f
C3250 a_15227_44166# a_19692_46634# 0.116169f
C3251 a_19333_46634# a_19466_46812# 0.167526f
C3252 a_5147_45002# a_5244_44056# 0.122327f
C3253 a_5883_43914# a_8975_43940# 0.50976f
C3254 a_n2497_47436# a_1423_45028# 1.36987f
C3255 a_8953_45546# a_9290_44172# 0.373944f
C3256 a_16327_47482# a_n2017_45002# 0.209709f
C3257 a_13507_46334# a_2437_43646# 0.117533f
C3258 COMP_P a_n784_42308# 0.109134f
C3259 a_1568_43370# VDD 0.433732f
C3260 a_20411_46873# a_3357_43084# 0.157199f
C3261 a_22400_42852# a_22589_40599# 0.135364f
C3262 a_10809_44734# VDD 2.67671f
C3263 a_n863_45724# a_413_45260# 0.140312f
C3264 a_n4209_39590# VREF 0.860047f
C3265 a_n237_47217# a_8667_46634# 0.171086f
C3266 a_n4209_39304# VDD 0.984278f
C3267 a_3754_38470# a_4338_37500# 0.473597f
C3268 a_n3420_37440# a_n2946_37690# 0.236674f
C3269 a_n97_42460# a_15743_43084# 0.205305f
C3270 a_20193_45348# a_21887_42336# 0.169001f
C3271 a_5147_45002# a_5111_44636# 0.562127f
C3272 a_4558_45348# a_4927_45028# 0.123258f
C3273 a_3537_45260# a_3232_43370# 0.530258f
C3274 a_16327_47482# a_19164_43230# 0.292734f
C3275 a_9290_44172# a_9028_43914# 0.169653f
C3276 a_4883_46098# a_8016_46348# 0.289691f
C3277 a_5883_43914# VDD 0.859221f
C3278 a_3080_42308# COMP_P 4.43537f
C3279 a_n743_46660# a_n443_42852# 0.378464f
C3280 a_n1741_47186# a_2437_43646# 4.86702f
C3281 a_n2157_46122# a_n1076_46494# 0.102355f
C3282 a_n1991_46122# a_n1641_46494# 0.219633f
C3283 a_13467_32519# a_13258_32519# 11.0084f
C3284 a_5343_44458# a_7845_44172# 0.103601f
C3285 a_3537_45260# a_4905_42826# 0.339989f
C3286 a_n881_46662# VDD 2.6692f
C3287 a_22959_46124# a_20692_30879# 0.155635f
C3288 a_5204_45822# a_5263_45724# 0.109078f
C3289 a_11415_45002# EN_OFFSET_CAL 0.14622f
C3290 a_n2157_46122# VDD 0.42567f
C3291 a_8049_45260# a_22959_45572# 0.176374f
C3292 a_768_44030# a_453_43940# 0.110708f
C3293 a_n1741_47186# a_n2661_46634# 0.22396f
C3294 a_4093_43548# a_4235_43370# 0.515101f
C3295 a_8162_45546# VDD 0.266272f
C3296 a_n2293_46098# a_5663_43940# 0.142661f
C3297 C7_P_btm VREF_GND 1.61142f
C3298 C4_P_btm VIN_P 0.50261f
C3299 C8_N_btm C10_N_btm 2.07867f
C3300 C6_N_btm VDD 0.210613f
C3301 a_768_44030# a_3090_45724# 0.115303f
C3302 C8_P_btm VCM 2.61094f
C3303 a_n1925_46634# a_6755_46942# 0.12389f
C3304 a_10227_46804# a_21363_46634# 0.273017f
C3305 C6_P_btm VREF 1.41944f
C3306 a_526_44458# a_n97_42460# 0.277959f
C3307 a_5205_44484# a_5518_44484# 0.135771f
C3308 a_2889_44172# VDD 0.1447f
C3309 a_2063_45854# CLK 0.271193f
C3310 a_n443_46116# VDD 3.87014f
C3311 a_n2956_39304# a_n2956_38680# 0.163045f
C3312 a_6171_42473# a_5932_42308# 0.224949f
C3313 a_17609_46634# VDD 0.501057f
C3314 a_167_45260# a_n37_45144# 0.277898f
C3315 a_n3565_39304# a_n3690_39392# 0.247167f
C3316 a_n4318_37592# VDD 0.919667f
C3317 a_19443_46116# VDD 0.132317f
C3318 a_n1059_45260# a_18057_42282# 0.141112f
C3319 a_13259_45724# a_16922_45042# 0.401687f
C3320 a_526_44458# a_742_44458# 0.54618f
C3321 a_7499_43078# a_5111_44636# 0.753731f
C3322 VDAC_P C3_P_btm 6.90991f
C3323 a_n4334_37440# VDD 0.385859f
C3324 a_n2293_46634# a_n2312_38680# 0.131017f
C3325 a_n1741_47186# a_765_45546# 0.536367f
C3326 a_n1613_43370# a_4651_46660# 0.686447f
C3327 a_3537_45260# VDD 3.9063f
C3328 a_n1059_45260# a_18494_42460# 0.187733f
C3329 a_5807_45002# a_2324_44458# 0.232399f
C3330 a_15227_44166# a_19466_46812# 0.310201f
C3331 a_2982_43646# a_5742_30871# 0.196805f
C3332 a_9290_44172# a_5534_30871# 0.472376f
C3333 a_10157_44484# a_10334_44484# 0.159555f
C3334 a_4791_45118# a_3232_43370# 0.268929f
C3335 a_n1853_46287# a_n1736_46482# 0.170096f
C3336 a_9625_46129# a_9823_46155# 0.321686f
C3337 a_n1151_42308# a_6709_45028# 0.286957f
C3338 a_1049_43396# VDD 0.196328f
C3339 a_14539_43914# a_15493_43940# 0.625897f
C3340 a_20107_42308# a_7174_31319# 0.175129f
C3341 a_n2833_47464# a_n2497_47436# 0.217831f
C3342 a_22223_46124# VDD 0.300745f
C3343 a_4791_45118# a_4905_42826# 0.516502f
C3344 a_1273_38525# VDD 3.23397f
C3345 a_3754_38470# a_3726_37500# 0.554457f
C3346 VDAC_Ni a_5088_37509# 1.70462f
C3347 a_n3565_37414# a_n4064_37440# 0.230258f
C3348 a_16327_47482# a_19339_43156# 0.346029f
C3349 a_n443_42852# a_5891_43370# 0.175668f
C3350 a_n1613_43370# a_n1076_46494# 0.232314f
C3351 a_n743_46660# a_765_45546# 0.148721f
C3352 a_8701_44490# VDD 0.164475f
C3353 a_685_42968# a_791_42968# 0.13675f
C3354 a_n1991_46122# a_n1423_46090# 0.175891f
C3355 a_n2293_42282# a_1755_42282# 0.875855f
C3356 a_n1613_43370# VDD 4.75085f
C3357 a_4646_46812# a_3537_45260# 0.361823f
C3358 a_n746_45260# a_n356_44636# 0.418585f
C3359 a_9290_44172# a_n443_42852# 0.483812f
C3360 a_15227_44166# a_16147_45260# 0.282941f
C3361 a_n1533_42852# VDD 0.142813f
C3362 a_n2293_46098# VDD 1.7963f
C3363 a_8049_45260# a_19963_31679# 0.2062f
C3364 a_n2497_47436# a_n2293_46634# 0.174929f
C3365 a_4958_30871# C9_P_btm 0.209166f
C3366 a_10227_46804# a_13507_46334# 0.120657f
C3367 a_22485_38105# a_22613_38993# 0.253409f
C3368 a_2684_37794# VDAC_Pi 0.133177f
C3369 a_n97_42460# a_3626_43646# 0.394673f
C3370 a_19479_31679# a_19963_31679# 0.104687f
C3371 a_3357_43084# a_22591_45572# 0.181818f
C3372 a_13661_43548# a_13667_43396# 0.168674f
C3373 a_526_44458# a_n2661_43922# 0.154533f
C3374 C5_P_btm VIN_P 0.502041f
C3375 C7_N_btm C10_N_btm 1.39624f
C3376 C8_N_btm C9_N_btm 39.4538f
C3377 C5_N_btm VDD 0.267489f
C3378 C8_P_btm VREF_GND 2.58605f
C3379 C9_P_btm VCM 6.06251f
C3380 C7_P_btm VREF 1.818f
C3381 a_10227_46804# a_20623_46660# 0.156341f
C3382 a_n443_46116# a_n901_46420# 0.367344f
C3383 a_3422_30871# a_13258_32519# 0.410904f
C3384 a_n443_42852# a_10807_43548# 0.173997f
C3385 a_5205_44484# a_5343_44458# 0.129692f
C3386 a_10249_46116# a_10355_46116# 0.182836f
C3387 a_4361_42308# a_4921_42308# 0.472085f
C3388 a_2675_43914# VDD 0.200923f
C3389 a_n1925_42282# a_n2293_42282# 0.234055f
C3390 a_4791_45118# VDD 3.05095f
C3391 a_5755_42308# a_5932_42308# 0.196877f
C3392 a_n2956_39304# a_n3565_39304# 0.307358f
C3393 a_16292_46812# VDD 0.123916f
C3394 a_13259_45724# a_13163_45724# 0.166368f
C3395 a_n1736_42282# VDD 0.227152f
C3396 a_4915_47217# a_6151_47436# 0.783303f
C3397 a_n913_45002# a_17303_42282# 1.81467f
C3398 a_3090_45724# a_7542_44172# 0.137368f
C3399 a_8199_44636# a_5891_43370# 0.399007f
C3400 VDAC_P C4_P_btm 13.8049f
C3401 a_8530_39574# RST_Z 0.431385f
C3402 a_n881_46662# a_3877_44458# 0.142507f
C3403 a_n1613_43370# a_4646_46812# 1.38979f
C3404 a_n4209_37414# VDD 0.817366f
C3405 a_1568_43370# a_1847_42826# 0.153113f
C3406 a_3429_45260# VDD 0.142923f
C3407 a_1414_42308# a_1067_42314# 0.100434f
C3408 a_n1059_45260# a_18184_42460# 0.52106f
C3409 a_n863_45724# a_175_44278# 0.113317f
C3410 a_10227_46804# a_10586_45546# 0.306536f
C3411 a_n2129_44697# a_n2012_44484# 0.172424f
C3412 a_13747_46662# a_15765_45572# 0.5661f
C3413 a_n2497_47436# a_626_44172# 0.249352f
C3414 a_8199_44636# a_9290_44172# 0.516297f
C3415 a_9625_46129# a_9569_46155# 0.204034f
C3416 a_3483_46348# a_2324_44458# 0.668551f
C3417 a_3090_45724# a_n2661_45546# 0.561435f
C3418 a_1209_43370# VDD 0.191694f
C3419 a_768_44030# a_n699_43396# 1.37533f
C3420 a_16327_47482# a_9313_44734# 0.169217f
C3421 a_10903_43370# a_10907_45822# 0.199567f
C3422 a_18184_42460# a_19987_42826# 0.208392f
C3423 a_6945_45028# VDD 1.30257f
C3424 a_n913_45002# a_2713_42308# 0.291963f
C3425 a_13661_43548# a_15493_43396# 0.491785f
C3426 a_n881_46662# a_8128_46384# 0.206292f
C3427 a_4791_45118# a_4646_46812# 0.485113f
C3428 a_n4209_39590# VIN_P 0.105382f
C3429 a_n4064_40160# VCM 0.121302f
C3430 VDAC_Ni a_4338_37500# 0.640521f
C3431 a_7754_38636# a_5088_37509# 0.288061f
C3432 a_n4334_37440# a_n4064_37440# 0.448688f
C3433 a_n3690_37440# a_n3420_37440# 0.431074f
C3434 a_n3565_37414# a_n2946_37690# 0.407439f
C3435 a_n4209_37414# a_n2302_37690# 0.407594f
C3436 a_21811_47423# a_20916_46384# 0.109084f
C3437 a_10227_46804# a_n743_46660# 0.134234f
C3438 a_19319_43548# a_4190_30871# 0.188868f
C3439 a_16327_47482# a_18599_43230# 0.182696f
C3440 a_3537_45260# a_4927_45028# 0.216859f
C3441 a_15861_45028# a_16922_45042# 0.259169f
C3442 a_584_46384# a_n1925_42282# 0.194054f
C3443 a_n1613_43370# a_n901_46420# 0.406381f
C3444 a_n237_47217# a_5066_45546# 1.48406f
C3445 a_n3674_39768# a_n4064_39616# 0.464693f
C3446 a_8103_44636# VDD 0.124028f
C3447 a_n863_45724# a_n97_42460# 0.581863f
C3448 a_n2157_46122# a_n1641_46494# 0.105995f
C3449 a_8270_45546# a_5066_45546# 0.189476f
C3450 a_n2293_42282# a_1606_42308# 0.192228f
C3451 a_3877_44458# a_3537_45260# 0.12249f
C3452 a_2107_46812# a_9482_43914# 0.109711f
C3453 a_22365_46825# EN_OFFSET_CAL 0.195393f
C3454 a_n2472_46090# VDD 0.224658f
C3455 a_6151_47436# a_n881_46662# 1.58776f
C3456 a_14456_42282# VDD 0.265543f
C3457 a_22485_38105# a_22581_37893# 0.902394f
C3458 a_6812_45938# VDD 0.132317f
C3459 a_n863_45724# a_742_44458# 0.629795f
C3460 a_10227_46804# a_20841_46902# 0.164019f
C3461 a_18479_47436# a_20411_46873# 0.192791f
C3462 C6_P_btm VIN_P 0.391898f
C3463 C7_N_btm C9_N_btm 0.22201f
C3464 C6_N_btm C10_N_btm 0.895671f
C3465 C4_N_btm VDD 0.265463f
C3466 C8_P_btm VREF 3.6701f
C3467 C9_P_btm VREF_GND 5.18245f
C3468 C10_P_btm VCM 10.5945f
C3469 a_5111_44636# a_5883_43914# 0.281106f
C3470 a_3232_43370# a_6298_44484# 0.256727f
C3471 a_n357_42282# a_19862_44208# 0.138067f
C3472 a_16327_47482# a_2711_45572# 0.101699f
C3473 a_895_43940# VDD 0.318652f
C3474 a_n2293_46634# a_3357_43084# 0.963711f
C3475 a_n913_45002# a_10796_42968# 0.545674f
C3476 a_15559_46634# VDD 0.301657f
C3477 a_n3674_38216# VDD 0.309006f
C3478 a_4791_45118# a_6545_47178# 0.112353f
C3479 a_3422_30871# a_4190_30871# 12.909901f
C3480 a_2711_45572# a_14537_43396# 0.249285f
C3481 a_3090_45724# a_7281_43914# 0.170855f
C3482 a_n2661_46634# a_n1925_46634# 4.75867f
C3483 VDAC_P C5_P_btm 27.6071f
C3484 a_8530_39574# VDD 0.346613f
C3485 a_n2109_47186# a_765_45546# 0.126431f
C3486 a_n1613_43370# a_3877_44458# 1.43013f
C3487 a_3065_45002# VDD 0.501045f
C3488 a_11823_42460# a_n2293_43922# 0.494696f
C3489 a_n2017_45002# a_18184_42460# 0.205351f
C3490 a_7229_43940# a_n2293_42834# 0.148023f
C3491 a_n743_46660# a_8016_46348# 0.155955f
C3492 a_11823_42460# a_n97_42460# 0.324041f
C3493 a_8199_44636# a_10355_46116# 0.176325f
C3494 a_18597_46090# a_3357_43084# 0.160577f
C3495 a_458_43396# VDD 0.431902f
C3496 a_3067_47026# VDD 0.132018f
C3497 a_768_44030# a_4223_44672# 0.136643f
C3498 a_10227_46804# a_5891_43370# 0.2393f
C3499 a_21137_46414# VDD 0.219745f
C3500 a_n4064_40160# VREF_GND 0.493568f
C3501 VDAC_Ni a_3726_37500# 1.5261f
C3502 a_n4209_37414# a_n4064_37440# 0.265895f
C3503 a_n3565_37414# a_n3420_37440# 0.307576f
C3504 a_4883_46098# a_20916_46384# 0.471396f
C3505 a_16327_47482# a_18817_42826# 0.215236f
C3506 a_3537_45260# a_5111_44636# 1.36722f
C3507 a_8696_44636# a_16922_45042# 0.10244f
C3508 a_n863_45724# a_n2661_43922# 0.115404f
C3509 a_584_46384# a_526_44458# 0.458472f
C3510 a_n1613_43370# a_n1641_46494# 0.152421f
C3511 a_12861_44030# a_2324_44458# 0.95556f
C3512 a_10227_46804# a_9290_44172# 0.918064f
C3513 a_6298_44484# VDD 1.21616f
C3514 a_13059_46348# a_13759_46122# 0.249771f
C3515 a_n1853_46287# a_n1991_46122# 0.737461f
C3516 a_19692_46634# a_6945_45028# 0.669658f
C3517 a_4190_30871# a_7174_31319# 0.153555f
C3518 a_3065_45002# a_3080_42308# 0.171466f
C3519 a_13507_46334# a_11827_44484# 0.384415f
C3520 a_22223_46124# a_20205_31679# 0.160234f
C3521 a_11415_45002# a_11823_42460# 0.349238f
C3522 a_1115_44172# a_1241_43940# 0.143754f
C3523 a_10193_42453# a_13575_42558# 0.175489f
C3524 a_n2840_46090# VDD 0.295278f
C3525 a_12861_44030# a_19862_44208# 0.721035f
C3526 a_9290_44172# a_1307_43914# 0.122831f
C3527 a_n4064_37984# a_n2302_37984# 0.250408f
C3528 a_13575_42558# VDD 0.182133f
C3529 a_6151_47436# a_n1613_43370# 0.548675f
C3530 a_n1151_42308# a_12549_44172# 0.466584f
C3531 a_2479_44172# a_2905_42968# 0.163227f
C3532 a_n97_42460# a_2982_43646# 0.180648f
C3533 a_18597_46090# a_19123_46287# 0.188676f
C3534 C7_P_btm VIN_P 1.52449f
C3535 C7_N_btm C8_N_btm 31.072699f
C3536 C5_N_btm C10_N_btm 0.51798f
C3537 C6_N_btm C9_N_btm 0.165353f
C3538 C3_N_btm VDD 0.26836f
C3539 a_2063_45854# a_167_45260# 0.359284f
C3540 C9_P_btm VREF 7.369471f
C3541 C10_P_btm VREF_GND 10.3207f
C3542 a_20301_43646# a_20556_43646# 0.114664f
C3543 a_5649_42852# a_5379_42460# 0.35554f
C3544 a_2479_44172# VDD 0.431428f
C3545 a_13720_44458# a_13857_44734# 0.126609f
C3546 a_4007_47204# VDD 0.41212f
C3547 a_768_44030# a_413_45260# 0.182253f
C3548 a_n1613_43370# a_5111_44636# 0.601769f
C3549 a_n2956_39304# a_n4209_39304# 0.328727f
C3550 a_15368_46634# VDD 0.324877f
C3551 a_4646_46812# a_6298_44484# 1.65052f
C3552 a_16327_47482# a_20512_43084# 0.118893f
C3553 a_4185_45028# a_n913_45002# 0.855072f
C3554 a_13259_45724# a_11823_42460# 0.626941f
C3555 a_n4209_39304# a_n3565_39304# 6.82668f
C3556 a_n2104_42282# VDD 0.280329f
C3557 a_5937_45572# a_6109_44484# 0.163331f
C3558 a_2711_45572# a_14180_45002# 0.147337f
C3559 a_8016_46348# a_5891_43370# 0.183035f
C3560 a_n2661_46634# a_n2312_38680# 0.106815f
C3561 VDAC_P C6_P_btm 55.214397f
C3562 a_7754_38470# VDD 0.302129f
C3563 a_15681_43442# a_15781_43660# 0.167615f
C3564 a_2680_45002# VDD 0.145087f
C3565 a_18834_46812# a_15227_44166# 0.231715f
C3566 a_15279_43071# a_5342_30871# 0.214197f
C3567 a_3537_45260# a_3905_42865# 0.258917f
C3568 a_9290_44172# a_13635_43156# 0.394766f
C3569 a_4791_45118# a_5111_44636# 1.11355f
C3570 a_n229_43646# VDD 0.278436f
C3571 COMP_P a_n1329_42308# 0.232443f
C3572 a_19511_42282# a_7174_31319# 0.240861f
C3573 a_1467_44172# a_1427_43646# 0.104539f
C3574 a_13661_43548# a_18451_43940# 0.129334f
C3575 a_584_46384# a_3626_43646# 0.195961f
C3576 a_12549_44172# a_15493_43940# 0.932577f
C3577 a_n4315_30879# VCM 0.473529f
C3578 a_1666_39587# VDD 3.12922f
C3579 a_n3565_37414# a_n3690_37440# 0.247968f
C3580 a_21496_47436# a_20916_46384# 0.113102f
C3581 a_2382_45260# a_3232_43370# 0.239776f
C3582 a_4574_45260# a_4558_45348# 0.19344f
C3583 a_16327_47482# a_18249_42858# 0.315855f
C3584 a_9049_44484# a_8701_44490# 0.100038f
C3585 a_7499_43078# a_5883_43914# 0.100372f
C3586 a_6151_47436# a_6945_45028# 0.335681f
C3587 a_11599_46634# a_13925_46122# 0.549622f
C3588 a_n1613_43370# a_n1423_46090# 0.15966f
C3589 a_5518_44484# VDD 0.40715f
C3590 a_n913_45002# a_11967_42832# 0.156551f
C3591 a_11599_46634# a_15599_45572# 0.26676f
C3592 a_19692_46634# a_21137_46414# 0.242332f
C3593 a_n2157_46122# a_n1991_46122# 0.614266f
C3594 a_14815_43914# a_14673_44172# 0.173231f
C3595 a_3877_44458# a_3065_45002# 0.287919f
C3596 a_5891_43370# a_8791_43396# 0.194389f
C3597 a_768_44030# a_644_44056# 0.177755f
C3598 a_22485_38105# a_22527_39145# 0.984424f
C3599 a_5815_47464# a_n1613_43370# 0.360237f
C3600 a_13070_42354# VDD 0.18656f
C3601 a_18479_47436# a_19386_47436# 0.219411f
C3602 a_18780_47178# a_18597_46090# 0.175179f
C3603 a_13661_43548# a_9145_43396# 0.135139f
C3604 a_2711_45572# a_18494_42460# 0.1183f
C3605 a_n2293_46098# a_3905_42865# 0.237656f
C3606 C5_N_btm C9_N_btm 0.150576f
C3607 C4_N_btm C10_N_btm 0.703336f
C3608 C6_N_btm C8_N_btm 0.163943f
C3609 C2_N_btm VDD 0.268945f
C3610 C10_P_btm VREF 14.773f
C3611 C8_P_btm VIN_P 0.907642f
C3612 a_5205_44484# a_4223_44672# 0.235572f
C3613 a_3232_43370# a_5343_44458# 0.654021f
C3614 a_n1925_46634# a_8034_45724# 0.206805f
C3615 a_2127_44172# VDD 0.138239f
C3616 a_3815_47204# VDD 0.260661f
C3617 a_14537_43396# a_14955_43940# 0.104291f
C3618 a_22612_30879# a_20447_31679# 0.107874f
C3619 a_10809_44734# a_22959_46124# 0.172346f
C3620 a_8953_45546# a_8049_45260# 0.156816f
C3621 a_4921_42308# a_5932_42308# 0.194195f
C3622 a_n1794_35242# a_5742_30871# 1.85829f
C3623 a_14976_45028# VDD 0.484864f
C3624 a_3218_45724# a_3175_45822# 0.132424f
C3625 a_n2293_46098# a_5147_45002# 0.211057f
C3626 a_5937_45572# a_3357_43084# 0.257963f
C3627 a_4791_45118# a_3905_42865# 0.208831f
C3628 a_n4209_39304# a_n4334_39392# 0.253307f
C3629 a_n443_46116# a_5129_47502# 0.10632f
C3630 a_n4318_38216# VDD 0.538766f
C3631 a_18051_46116# VDD 0.189782f
C3632 a_7499_43078# a_3537_45260# 0.586701f
C3633 a_1823_45246# a_n2661_43922# 0.441151f
C3634 a_5807_45002# a_2107_46812# 1.5594f
C3635 a_n2472_46634# a_n2293_46634# 0.163804f
C3636 VDAC_P C7_P_btm 0.11042p
C3637 a_3754_38470# RST_Z 0.203816f
C3638 a_2382_45260# VDD 1.6285f
C3639 a_n97_42460# a_7227_42852# 0.117893f
C3640 a_n237_47217# a_1848_45724# 0.232571f
C3641 a_5534_30871# a_5342_30871# 11.128201f
C3642 a_15433_44458# VDD 0.201121f
C3643 a_3537_45260# a_3600_43914# 0.157156f
C3644 a_n2472_46090# a_n2956_38680# 0.157373f
C3645 a_4791_45118# a_5147_45002# 0.10845f
C3646 a_18479_47436# a_3357_43084# 0.292061f
C3647 a_3080_42308# C2_N_btm 0.108823f
C3648 a_3524_46660# VDD 0.278519f
C3649 a_18989_43940# a_18451_43940# 0.114286f
C3650 a_n2661_43922# a_n3674_39768# 0.152656f
C3651 a_19900_46494# VDD 0.279179f
C3652 a_n755_45592# a_n913_45002# 0.347782f
C3653 a_n1151_42308# a_n1557_42282# 0.214486f
C3654 a_n4209_37414# a_n3420_37440# 0.245806f
C3655 a_13507_46334# a_20916_46384# 0.123008f
C3656 a_n4315_30879# VREF_GND 0.168163f
C3657 a_n971_45724# a_7577_46660# 0.523694f
C3658 a_1169_39587# VDD 0.531695f
C3659 a_3537_45260# a_4558_45348# 0.236111f
C3660 a_n881_46662# a_n1853_46287# 0.229188f
C3661 a_11599_46634# a_13759_46122# 0.262969f
C3662 a_5343_44458# VDD 0.49245f
C3663 a_n1059_45260# a_11967_42832# 0.627158f
C3664 a_n2293_46634# a_n443_42852# 2.09483f
C3665 a_n1613_43370# a_7499_43078# 0.324998f
C3666 a_19692_46634# a_20708_46348# 0.318388f
C3667 a_n2157_46122# a_n1853_46287# 0.617317f
C3668 a_n357_42282# a_21356_42826# 0.156735f
C3669 a_12861_44030# a_15493_43396# 0.254093f
C3670 a_22485_38105# a_22589_40055# 0.212168f
C3671 a_4915_47217# a_n881_46662# 1.23372f
C3672 a_12563_42308# VDD 0.254292f
C3673 a_n1151_42308# a_11309_47204# 0.546434f
C3674 a_18479_47436# a_18597_46090# 0.473843f
C3675 a_2479_44172# a_1847_42826# 0.141223f
C3676 a_2437_43646# a_3357_43084# 0.424652f
C3677 a_22223_45572# a_19479_31679# 0.155323f
C3678 a_2711_45572# a_18184_42460# 0.367034f
C3679 a_12465_44636# a_13059_46348# 0.163448f
C3680 a_10227_46804# a_20107_46660# 0.312495f
C3681 C6_N_btm C7_N_btm 26.0771f
C3682 C5_N_btm C8_N_btm 0.145019f
C3683 C3_N_btm C10_N_btm 0.321945f
C3684 C4_N_btm C9_N_btm 0.154834f
C3685 C1_N_btm VDD 0.264503f
C3686 C9_P_btm VIN_P 1.82823f
C3687 a_4190_30871# a_743_42282# 0.18536f
C3688 a_453_43940# VDD 0.225569f
C3689 a_3785_47178# VDD 0.387755f
C3690 a_18494_42460# a_20512_43084# 0.115057f
C3691 a_12465_44636# a_13556_45296# 0.248126f
C3692 a_2324_44458# a_526_44458# 0.279023f
C3693 a_5937_45572# a_8049_45260# 0.103218f
C3694 a_3090_45724# VDD 2.05725f
C3695 a_2889_44172# a_2998_44172# 0.179664f
C3696 a_3218_45724# a_2711_45572# 0.1731f
C3697 a_4646_46812# a_5343_44458# 0.24395f
C3698 a_6755_46942# a_11691_44458# 0.192426f
C3699 a_n2472_42282# VDD 0.278905f
C3700 a_n443_46116# a_4915_47217# 0.395101f
C3701 a_4791_45118# a_5129_47502# 0.240381f
C3702 a_1823_45246# a_n2661_42834# 0.174801f
C3703 a_n2472_46634# a_n2442_46660# 0.155358f
C3704 a_3754_38470# VDD 2.52245f
C3705 VDAC_P C8_P_btm 0.220914p
C3706 a_2274_45254# VDD 0.256655f
C3707 a_n97_42460# a_5755_42852# 0.149651f
C3708 a_n2661_46098# a_1176_45822# 0.144277f
C3709 a_2107_46812# a_3483_46348# 0.100707f
C3710 a_14815_43914# VDD 0.307386f
C3711 a_3232_43370# a_1414_42308# 0.248035f
C3712 a_5937_45572# a_8953_45546# 0.3871f
C3713 a_3699_46634# VDD 0.347281f
C3714 a_n2661_42834# a_n3674_39768# 0.150968f
C3715 a_768_44030# a_742_44458# 0.216263f
C3716 a_9290_44172# a_10907_45822# 0.262972f
C3717 a_19647_42308# a_13258_32519# 0.153411f
C3718 a_20075_46420# VDD 0.347847f
C3719 a_n755_45592# a_n1059_45260# 0.53237f
C3720 a_n357_42282# a_n913_45002# 0.309845f
C3721 a_n443_46116# a_1568_43370# 0.584982f
C3722 a_3483_46348# a_n2661_44458# 1.44355f
C3723 a_12549_44172# a_11341_43940# 0.406618f
C3724 a_n1151_42308# a_4955_46873# 0.261025f
C3725 a_n4315_30879# VREF 1.73216f
C3726 a_n356_44636# a_6123_31319# 0.169259f
C3727 a_16327_47482# a_18083_42858# 0.591108f
C3728 a_3537_45260# a_4574_45260# 0.234297f
C3729 a_11599_46634# a_13351_46090# 0.105205f
C3730 a_4646_46812# a_3090_45724# 0.199722f
C3731 a_n1613_43370# a_n1853_46287# 0.354256f
C3732 a_4743_44484# VDD 0.266843f
C3733 a_n3674_39768# a_n3565_39590# 0.128683f
C3734 a_13507_46334# a_18907_42674# 0.202065f
C3735 a_18597_46090# a_19511_42282# 0.156698f
C3736 a_15227_44166# a_6945_45028# 0.548194f
C3737 a_3877_44458# a_2382_45260# 0.395451f
C3738 a_11453_44696# a_17719_45144# 0.105851f
C3739 a_3090_45724# a_18479_45785# 0.259218f
C3740 a_11415_45002# a_11652_45724# 0.128811f
C3741 a_8953_45546# a_n443_42852# 0.134632f
C3742 a_21076_30879# VDD 1.17053f
C3743 a_3090_45724# a_10057_43914# 0.230475f
C3744 a_2324_44458# a_8953_45002# 1.65784f
C3745 a_n3420_37984# a_n4064_37984# 8.18485f
C3746 a_n443_46116# a_n881_46662# 0.114922f
C3747 a_4915_47217# a_n1613_43370# 0.195064f
C3748 a_11633_42558# VDD 0.193501f
C3749 C5_N_btm C7_N_btm 0.151416f
C3750 C2_N_btm C10_N_btm 0.327137f
C3751 C3_N_btm C9_N_btm 0.137552f
C3752 C4_N_btm C8_N_btm 0.145646f
C3753 C0_N_btm VDD 1.02806f
C3754 C10_P_btm VIN_P 3.66034f
C3755 a_n2661_46634# a_6755_46942# 1.40968f
C3756 a_12861_44030# a_18280_46660# 0.140921f
C3757 a_5111_44636# a_5518_44484# 0.124556f
C3758 a_768_44030# a_13259_45724# 0.315247f
C3759 a_1414_42308# VDD 0.657887f
C3760 a_17730_32519# VREF_GND 0.241027f
C3761 a_11823_42460# a_14205_43396# 0.176571f
C3762 a_13076_44458# a_13213_44734# 0.126609f
C3763 a_3381_47502# VDD 0.197761f
C3764 a_4791_45118# a_n2661_43370# 0.408007f
C3765 a_12281_43396# VDD 0.341026f
C3766 a_4921_42308# a_5755_42308# 0.175841f
C3767 a_15009_46634# VDD 0.205396f
C3768 a_2675_43914# a_2998_44172# 0.173844f
C3769 a_768_44030# a_n2661_43922# 1.9176f
C3770 a_12549_44172# a_n2293_43922# 0.194293f
C3771 a_4791_45118# a_4915_47217# 0.226891f
C3772 a_2063_45854# a_9863_47436# 0.12173f
C3773 a_n3674_38680# VDD 0.503323f
C3774 a_n784_42308# C0_N_btm 0.281635f
C3775 a_12741_44636# a_14673_44172# 0.178572f
C3776 VDAC_P C9_P_btm 0.441881p
C3777 a_1667_45002# VDD 0.315476f
C3778 a_n237_47217# a_n755_45592# 0.286948f
C3779 a_n2840_46090# a_n2956_39304# 0.158668f
C3780 a_10227_46804# a_3357_43084# 0.305304f
C3781 a_8199_44636# a_8953_45546# 0.71291f
C3782 a_17538_32519# VREF_GND 0.117023f
C3783 a_2959_46660# VDD 0.19762f
C3784 a_n1613_43370# a_5883_43914# 0.352323f
C3785 a_19335_46494# VDD 0.198512f
C3786 a_n357_42282# a_n1059_45260# 7.3759f
C3787 a_1609_45822# a_2437_43646# 0.189329f
C3788 a_12741_44636# a_12607_44458# 0.134974f
C3789 a_12549_44172# a_21115_43940# 0.211261f
C3790 a_n4209_37414# a_n3565_37414# 6.90997f
C3791 a_16327_47482# a_n743_46660# 0.53683f
C3792 a_n1613_43370# a_n881_46662# 1.06426f
C3793 a_n971_45724# a_7411_46660# 0.567031f
C3794 a_10227_46804# a_5342_30871# 0.163388f
C3795 a_3357_43084# a_1307_43914# 0.197864f
C3796 a_n881_46662# a_n2293_46098# 0.291354f
C3797 a_4915_47217# a_6945_45028# 0.207881f
C3798 a_n1613_43370# a_n2157_46122# 0.296124f
C3799 a_3877_44458# a_3090_45724# 0.23348f
C3800 a_n699_43396# VDD 0.922998f
C3801 a_18114_32519# VCM 0.121302f
C3802 a_13059_46348# a_10903_43370# 0.11738f
C3803 a_n743_46660# a_n356_45724# 0.223429f
C3804 a_12861_44030# a_15903_45785# 0.156145f
C3805 a_22959_43948# VDD 0.297936f
C3806 SMPL_ON_N VIN_N 0.546477f
C3807 a_n2293_46634# a_1307_43914# 0.184387f
C3808 a_3090_45724# a_18175_45572# 0.130163f
C3809 a_n4318_38680# VDD 0.417422f
C3810 a_13575_42558# a_14113_42308# 0.11418f
C3811 a_22959_46660# VDD 0.299681f
C3812 a_10193_42453# a_11551_42558# 0.228057f
C3813 a_2324_44458# a_8191_45002# 0.120399f
C3814 a_n3420_37984# a_n2946_37984# 0.238664f
C3815 a_4791_45118# a_n881_46662# 0.429542f
C3816 a_n443_46116# a_n1613_43370# 0.410263f
C3817 a_12861_44030# a_11453_44696# 0.173308f
C3818 a_11551_42558# VDD 0.192086f
C3819 a_15493_43396# a_15743_43084# 0.517624f
C3820 a_2437_43646# a_22223_45572# 0.165664f
C3821 a_n443_46116# a_n2293_46098# 0.251135f
C3822 a_19998_35138# VIN_N 0.37444f
C3823 C4_N_btm C7_N_btm 0.145303f
C3824 C1_N_btm C10_N_btm 0.31753f
C3825 C2_N_btm C9_N_btm 0.141891f
C3826 C3_N_btm C8_N_btm 0.134581f
C3827 a_584_46384# a_1138_42852# 0.491749f
C3828 C5_N_btm C6_N_btm 22.305399f
C3829 EN_VIN_BSTR_N VCM 0.927954f
C3830 a_5111_44636# a_5343_44458# 0.477401f
C3831 a_12549_44172# a_13259_45724# 0.110646f
C3832 a_n1151_42308# a_10193_42453# 0.238612f
C3833 a_1467_44172# VDD 0.391994f
C3834 a_11823_42460# a_14358_43442# 0.122636f
C3835 a_n1151_42308# VDD 2.57238f
C3836 a_21076_30879# a_20692_30879# 0.117886f
C3837 a_6945_45028# a_10809_44734# 0.953135f
C3838 a_768_44030# a_n2661_42834# 4.99505f
C3839 a_4791_45118# a_n443_46116# 0.115639f
C3840 a_n2840_42282# VDD 0.294987f
C3841 a_7227_45028# a_6709_45028# 0.115677f
C3842 VDAC_P C10_P_btm 0.883474p
C3843 a_n2956_39768# a_n2442_46660# 6.5214f
C3844 VDAC_Ni VDD 0.288547f
C3845 a_22629_38406# a_22629_37990# 0.32625f
C3846 a_10227_46804# a_6755_46942# 0.778648f
C3847 a_327_44734# VDD 0.667364f
C3848 a_413_45260# RST_Z 0.199496f
C3849 a_3065_45002# a_n2661_43370# 0.356646f
C3850 a_4185_45028# a_20974_43370# 0.184625f
C3851 a_n1151_42308# a_n784_42308# 0.154055f
C3852 a_n746_45260# a_n755_45592# 0.172774f
C3853 a_n881_46662# a_6945_45028# 0.239384f
C3854 a_13857_44734# VDD 0.18416f
C3855 a_14543_43071# a_5534_30871# 0.196814f
C3856 a_2382_45260# a_3905_42865# 0.291572f
C3857 a_4791_45118# a_3537_45260# 0.33264f
C3858 a_8199_44636# a_5937_45572# 0.573373f
C3859 a_8016_46348# a_9625_46129# 0.128435f
C3860 a_n1809_43762# VDD 0.142403f
C3861 a_n1736_42282# a_n4318_37592# 0.153911f
C3862 a_n3674_39304# a_n4064_39072# 0.539144f
C3863 a_3177_46902# VDD 0.200982f
C3864 a_n4318_37592# a_n4209_37414# 0.105251f
C3865 a_133_42852# VDD 0.184203f
C3866 a_n913_45002# a_1755_42282# 0.169955f
C3867 a_19553_46090# VDD 0.204238f
C3868 a_n2293_45546# a_n967_45348# 0.119714f
C3869 a_n357_42282# a_n2017_45002# 0.580077f
C3870 a_12549_44172# a_20935_43940# 0.110704f
C3871 a_n2302_39866# VDD 0.361509f
C3872 a_12465_44636# a_13661_43548# 0.106973f
C3873 a_n4209_37414# a_n4334_37440# 0.253282f
C3874 a_n4315_30879# VIN_P 0.187185f
C3875 a_n1151_42308# a_4646_46812# 0.330834f
C3876 a_3429_45260# a_3537_45260# 0.138977f
C3877 a_10467_46802# a_6755_46942# 0.256039f
C3878 a_11599_46634# a_12005_46116# 0.27095f
C3879 a_4883_46098# a_4704_46090# 0.1774f
C3880 a_4223_44672# VDD 2.99073f
C3881 a_18114_32519# VREF_GND 0.493553f
C3882 a_10193_42453# a_15493_43940# 0.597095f
C3883 a_15227_44166# a_20708_46348# 0.106656f
C3884 a_13661_43548# a_2711_45572# 0.552383f
C3885 a_15493_43940# VDD 1.4617f
C3886 a_9313_44734# a_11967_42832# 0.216837f
C3887 a_4185_45028# a_2711_45572# 0.102913f
C3888 a_11415_45002# a_11322_45546# 0.527707f
C3889 a_4791_45118# a_8701_44490# 0.138973f
C3890 a_13507_46334# a_18494_42460# 0.234442f
C3891 a_3483_46348# a_4099_45572# 0.15767f
C3892 a_8034_45724# a_8049_45260# 0.141057f
C3893 a_n3674_39304# VDD 0.587205f
C3894 a_n3674_38680# a_n3420_39072# 0.172947f
C3895 a_13575_42558# a_13657_42558# 0.171361f
C3896 a_16922_45042# a_20749_43396# 0.106779f
C3897 a_12741_44636# VDD 0.988199f
C3898 a_10193_42453# a_5742_30871# 0.303452f
C3899 a_10903_43370# a_9482_43914# 1.20611f
C3900 a_22485_38105# a_22589_40599# 0.132855f
C3901 a_n3565_38216# a_n4064_37984# 0.342209f
C3902 a_4791_45118# a_n1613_43370# 0.223884f
C3903 a_584_46384# a_768_44030# 0.105366f
C3904 a_5934_30871# VCM 0.121361f
C3905 a_n1151_42308# a_9804_47204# 0.108722f
C3906 a_5742_30871# VDD 0.557144f
C3907 a_18143_47464# a_18479_47436# 0.238309f
C3908 a_n97_42460# a_n1557_42282# 0.149645f
C3909 a_1209_43370# a_1049_43396# 0.194938f
C3910 a_526_44458# a_3363_44484# 0.119556f
C3911 a_17715_44484# a_17517_44484# 0.163303f
C3912 a_13259_45724# a_13076_44458# 0.188498f
C3913 a_13059_46348# a_13483_43940# 0.124566f
C3914 a_4791_45118# a_n2293_46098# 0.411939f
C3915 C3_N_btm C7_N_btm 0.134911f
C3916 C0_N_btm C10_N_btm 0.365593f
C3917 C1_N_btm C9_N_btm 0.132506f
C3918 C2_N_btm C8_N_btm 0.138777f
C3919 C4_N_btm C6_N_btm 0.143514f
C3920 EN_VIN_BSTR_N VREF_GND 0.857366f
C3921 a_n2293_42834# VDD 0.853754f
C3922 a_21259_43561# a_4190_30871# 0.198353f
C3923 a_3537_45260# a_8103_44636# 0.140404f
C3924 a_12891_46348# a_13259_45724# 1.04614f
C3925 a_17339_46660# a_18285_46348# 0.184197f
C3926 a_1115_44172# VDD 0.165092f
C3927 a_4361_42308# a_3823_42558# 0.114877f
C3928 a_11823_42460# a_14579_43548# 0.106967f
C3929 a_3160_47472# VDD 0.256092f
C3930 a_765_45546# a_n443_42852# 0.232932f
C3931 a_6945_45028# a_22223_46124# 0.17119f
C3932 a_n784_42308# a_5742_30871# 0.550812f
C3933 a_13607_46688# VDD 0.209568f
C3934 a_n1761_44111# a_n1644_44306# 0.170098f
C3935 a_n443_46116# a_895_43940# 0.163929f
C3936 a_16375_45002# a_10193_42453# 0.125364f
C3937 a_4700_47436# a_n443_46116# 0.255594f
C3938 a_16375_45002# VDD 1.14948f
C3939 a_10227_46804# a_10249_46116# 0.137273f
C3940 CAL_P a_22629_37990# 0.205295f
C3941 a_413_45260# VDD 1.203f
C3942 a_n971_45724# a_n755_45592# 0.347347f
C3943 a_2382_45260# a_3600_43914# 0.158274f
C3944 a_14035_46660# a_14180_46482# 0.157972f
C3945 a_n3674_38216# a_n4318_37592# 2.7294f
C3946 a_n4318_38680# a_n3420_39072# 0.310238f
C3947 a_2609_46660# VDD 0.312974f
C3948 a_19279_43940# a_21398_44850# 0.183186f
C3949 a_4646_46812# a_n2293_42834# 0.152973f
C3950 a_18985_46122# VDD 0.253642f
C3951 a_15143_45578# a_15037_45618# 0.13675f
C3952 a_n755_45592# a_n2293_45010# 0.159033f
C3953 a_n4064_39616# VDD 1.6861f
C3954 a_12465_44636# a_5807_45002# 0.59474f
C3955 a_3065_45002# a_3537_45260# 0.162384f
C3956 a_10227_46804# a_5534_30871# 0.304847f
C3957 a_10623_46897# a_10554_47026# 0.209641f
C3958 a_10428_46928# a_6755_46942# 0.155315f
C3959 a_10467_46802# a_10249_46116# 0.12624f
C3960 a_4791_45118# a_6945_45028# 0.493927f
C3961 a_11599_46634# a_10903_43370# 0.439916f
C3962 a_n2661_46634# a_765_45546# 1.82448f
C3963 a_n4318_39768# a_n4209_39590# 0.105246f
C3964 a_2779_44458# VDD 0.38604f
C3965 a_526_44458# a_9803_43646# 0.170855f
C3966 a_n2472_46090# a_n2293_46098# 0.176709f
C3967 a_14035_46660# a_13925_46122# 0.207108f
C3968 a_n2293_42282# a_n1794_35242# 0.18361f
C3969 a_22223_43948# VDD 0.254313f
C3970 a_5649_42852# a_4958_30871# 0.293366f
C3971 a_13291_42460# a_14635_42282# 0.111986f
C3972 a_n913_45002# a_3539_42460# 0.359316f
C3973 a_13507_46334# a_18184_42460# 0.505552f
C3974 a_n13_43084# VDD 0.260551f
C3975 a_20820_30879# VDD 0.719562f
C3976 a_526_44458# a_n913_45002# 0.250864f
C3977 a_5937_45572# a_1307_43914# 0.101589f
C3978 a_n1151_42308# a_8128_46384# 0.328697f
C3979 a_n4334_38304# a_n4064_37984# 0.410244f
C3980 a_n3690_38304# a_n3420_37984# 0.414894f
C3981 a_n3565_38216# a_n2946_37984# 0.411006f
C3982 a_n4209_38216# a_n2302_37984# 0.407312f
C3983 a_2684_37794# a_2113_38308# 0.468006f
C3984 a_13717_47436# SMPL_ON_N 0.132417f
C3985 a_11323_42473# VDD 0.205172f
C3986 a_10227_46804# a_18479_47436# 1.40697f
C3987 a_11599_46634# a_4883_46098# 0.261488f
C3988 a_19692_46634# a_15493_43940# 0.16692f
C3989 a_13507_46334# a_13059_46348# 0.192049f
C3990 C2_N_btm C7_N_btm 0.138288f
C3991 C0_dummy_N_btm C10_N_btm 0.749362f
C3992 C0_N_btm C9_N_btm 0.146135f
C3993 C1_N_btm C8_N_btm 0.129306f
C3994 C3_N_btm C6_N_btm 0.133742f
C3995 C4_N_btm C5_N_btm 18.6196f
C3996 C0_P_btm VDD 1.02806f
C3997 a_n971_45724# a_3483_46348# 0.211534f
C3998 a_n743_46660# a_5066_45546# 0.124676f
C3999 a_2063_45854# a_11322_45546# 0.105268f
C4000 a_644_44056# VDD 0.147321f
C4001 a_14543_43071# a_13291_42460# 0.107887f
C4002 a_3232_43370# a_11341_43940# 0.112367f
C4003 a_11823_42460# a_13667_43396# 0.107673f
C4004 a_1431_47204# DATA[1] 0.334099f
C4005 a_2905_45572# VDD 1.22598f
C4006 a_3090_45724# a_7499_43078# 0.23734f
C4007 a_5379_42460# a_5932_42308# 0.761308f
C4008 a_12816_46660# VDD 0.293798f
C4009 a_11967_42832# a_15682_43940# 1.63211f
C4010 a_6755_46942# a_11827_44484# 0.529579f
C4011 a_n443_46116# a_2479_44172# 0.732848f
C4012 a_n755_45592# a_2711_45572# 0.168218f
C4013 a_11415_45002# a_6171_45002# 1.05801f
C4014 a_16327_47482# a_3422_30871# 0.220296f
C4015 a_4700_47436# a_4791_45118# 0.31818f
C4016 a_20753_42852# VDD 0.193909f
C4017 a_n784_42308# C0_P_btm 0.281635f
C4018 a_11415_45002# a_14673_44172# 0.229077f
C4019 a_10227_46804# a_10554_47026# 0.166977f
C4020 a_n37_45144# VDD 0.138f
C4021 a_n971_45724# a_n357_42282# 0.271282f
C4022 a_584_46384# a_n2661_45546# 0.100439f
C4023 a_3090_45724# a_15227_44166# 0.428743f
C4024 a_n746_45260# a_310_45028# 0.378188f
C4025 a_13213_44734# VDD 0.184239f
C4026 a_10227_46804# a_2437_43646# 0.150025f
C4027 a_17701_42308# a_17531_42308# 0.109201f
C4028 a_104_43370# VDD 0.252393f
C4029 a_n1059_45260# a_15743_43084# 0.101833f
C4030 a_2443_46660# VDD 0.413663f
C4031 a_11967_42832# a_20512_43084# 0.106819f
C4032 a_3090_45724# a_4558_45348# 0.147318f
C4033 a_18819_46122# VDD 0.453432f
C4034 a_20692_30879# a_413_45260# 0.111034f
C4035 a_n2946_39866# VDD 0.393552f
C4036 a_20894_47436# a_20843_47204# 0.134298f
C4037 a_16223_45938# VDD 0.132317f
C4038 a_2437_43646# a_1307_43914# 0.160142f
C4039 a_n357_42282# a_9313_44734# 5.02008f
C4040 a_n237_47217# a_n1925_42282# 0.109762f
C4041 a_10428_46928# a_10249_46116# 0.704177f
C4042 a_12465_44636# a_3483_46348# 0.210833f
C4043 a_10227_46804# a_8199_44636# 0.460391f
C4044 a_949_44458# VDD 1.2275f
C4045 a_13507_46334# a_17303_42282# 1.68549f
C4046 a_4185_45028# a_5649_42852# 8.049951f
C4047 a_14035_46660# a_13759_46122# 0.162408f
C4048 a_11341_43940# VDD 1.23655f
C4049 a_n913_45002# a_3626_43646# 0.104422f
C4050 a_3232_43370# a_n97_42460# 0.113391f
C4051 a_3483_46348# a_2711_45572# 0.167588f
C4052 a_n1076_43230# VDD 0.292942f
C4053 COMP_P a_1169_39587# 0.388738f
C4054 a_21076_30879# C8_N_btm 0.384801f
C4055 a_22591_46660# VDD 0.251892f
C4056 a_2063_45854# a_11309_47204# 0.141276f
C4057 a_n4209_38216# a_n4064_37984# 0.19304f
C4058 a_n3565_38216# a_n3420_37984# 0.238595f
C4059 a_6123_31319# VCM 0.144585f
C4060 a_13717_47436# a_22731_47423# 0.109987f
C4061 a_10723_42308# VDD 0.223902f
C4062 a_10227_46804# a_18143_47464# 0.112443f
C4063 a_n97_42460# a_4905_42826# 0.147727f
C4064 a_13259_45724# a_12607_44458# 0.132105f
C4065 C1_N_btm C7_N_btm 0.128479f
C4066 C0_dummy_N_btm C9_N_btm 0.111645f
C4067 C0_N_btm C8_N_btm 0.146541f
C4068 a_584_46384# a_805_46414# 0.135394f
C4069 C2_N_btm C6_N_btm 0.137206f
C4070 C3_N_btm C5_N_btm 0.135528f
C4071 C1_P_btm VDD 0.264503f
C4072 EN_VIN_BSTR_N VIN_N 1.41696f
C4073 a_n2109_47186# a_5164_46348# 0.603312f
C4074 EN_VIN_BSTR_P VCM 0.929382f
C4075 a_5111_44636# a_4223_44672# 0.418299f
C4076 a_17339_46660# a_765_45546# 0.244447f
C4077 a_175_44278# VDD 0.20887f
C4078 a_20820_30879# a_20692_30879# 8.973741f
C4079 a_8199_44636# a_8034_45724# 0.127067f
C4080 a_10341_43396# VDD 0.401264f
C4081 a_5379_42460# a_6171_42473# 0.110293f
C4082 a_12991_46634# VDD 0.357655f
C4083 a_n913_45002# a_8037_42858# 0.316376f
C4084 a_n443_46116# a_2127_44172# 0.196411f
C4085 a_3090_45724# a_n2661_43370# 0.101361f
C4086 a_1666_39587# a_1273_38525# 0.277775f
C4087 a_n3420_39616# a_n4064_39072# 6.32746f
C4088 a_n2840_46634# a_n2661_46634# 0.180867f
C4089 a_10227_46804# a_10623_46897# 0.180903f
C4090 a_5111_44636# a_n2293_42834# 0.110286f
C4091 a_n1151_42308# a_n961_42308# 0.109068f
C4092 a_n2293_43922# VDD 0.735266f
C4093 a_10193_42453# a_n97_42460# 0.304653f
C4094 a_8016_46348# a_8199_44636# 0.33718f
C4095 a_n4318_38216# a_n4318_37592# 0.139499f
C4096 a_n97_42460# VDD 3.61113f
C4097 a_n2661_46098# VDD 0.979859f
C4098 a_17957_46116# VDD 0.138777f
C4099 a_11341_43940# a_14021_43940# 3.06514f
C4100 a_742_44458# a_2905_42968# 0.15065f
C4101 a_n2956_38216# a_n2956_37592# 0.103811f
C4102 a_n863_45724# a_n913_45002# 0.565852f
C4103 a_n3420_39616# VDD 0.568506f
C4104 a_4883_46098# a_5807_45002# 1.76125f
C4105 a_n97_42460# a_16137_43396# 0.134668f
C4106 a_n2293_43922# a_n784_42308# 1.67292f
C4107 a_10227_46804# a_13460_43230# 0.243111f
C4108 a_2382_45260# a_3537_45260# 0.250657f
C4109 a_3483_46348# a_15682_43940# 0.261013f
C4110 a_7715_46873# a_7832_46660# 0.157972f
C4111 a_12861_44030# a_12594_46348# 0.43362f
C4112 a_n237_47217# a_526_44458# 0.198088f
C4113 a_10428_46928# a_10554_47026# 0.181217f
C4114 a_10467_46802# a_10623_46897# 0.107482f
C4115 a_742_44458# VDD 1.3845f
C4116 a_3232_43370# a_n2661_43922# 0.197944f
C4117 a_11827_44484# a_11691_44458# 0.881979f
C4118 a_12465_44636# a_13249_42308# 0.541909f
C4119 a_21115_43940# VDD 0.145936f
C4120 a_n1794_35242# a_n4209_39590# 0.12484f
C4121 a_n901_43156# VDD 0.475947f
C4122 a_11415_45002# VDD 1.84504f
C4123 a_5891_43370# a_6293_42852# 0.107308f
C4124 a_10193_42453# a_10533_42308# 0.101629f
C4125 a_16375_45002# a_16147_45260# 1.01554f
C4126 a_3090_45724# a_5883_43914# 0.132458f
C4127 a_n3565_38216# a_n3690_38304# 0.247167f
C4128 a_12861_44030# a_12465_44636# 0.242761f
C4129 a_10533_42308# VDD 0.216201f
C4130 a_11599_46634# a_13507_46334# 0.259318f
C4131 a_11967_42832# a_17333_42852# 0.14149f
C4132 a_n97_42460# a_3080_42308# 0.353977f
C4133 a_14021_43940# a_10341_43396# 1.5617f
C4134 EN_VIN_BSTR_P VREF_GND 0.857366f
C4135 C0_N_btm C7_N_btm 0.140846f
C4136 C0_dummy_N_btm C8_N_btm 0.234177f
C4137 a_584_46384# a_472_46348# 0.31609f
C4138 C1_N_btm C6_N_btm 0.127656f
C4139 C3_N_btm C4_N_btm 9.61674f
C4140 C2_N_btm C5_N_btm 0.13795f
C4141 C2_P_btm VDD 0.268945f
C4142 a_11530_34132# VIN_N 1.547f
C4143 a_n881_46662# a_3090_45724# 0.107805f
C4144 a_3537_45260# a_5343_44458# 0.378482f
C4145 a_n1925_46634# a_5066_45546# 0.195997f
C4146 a_12861_44030# a_2711_45572# 0.104124f
C4147 a_n984_44318# VDD 0.281427f
C4148 a_8975_43940# a_n2661_43922# 0.11532f
C4149 a_2553_47502# VDD 0.150286f
C4150 a_9885_43646# VDD 0.190473f
C4151 a_12251_46660# VDD 0.195617f
C4152 a_2479_44172# a_895_43940# 0.318312f
C4153 a_1414_42308# a_2998_44172# 0.447595f
C4154 a_n2472_43914# a_n3674_39768# 0.162742f
C4155 a_13259_45724# a_10193_42453# 0.284945f
C4156 a_n1741_47186# a_11599_46634# 0.164599f
C4157 a_13259_45724# VDD 2.41738f
C4158 a_11823_42460# a_n913_45002# 0.281323f
C4159 a_n2840_46634# a_n2956_39768# 0.156182f
C4160 a_10227_46804# a_10467_46802# 0.678578f
C4161 a_22537_39537# a_22629_37990# 0.490939f
C4162 a_n1613_43370# a_3524_46660# 0.28004f
C4163 a_n467_45028# VDD 0.385804f
C4164 a_n1151_42308# a_n1329_42308# 0.167748f
C4165 a_12549_44172# a_2324_44458# 0.506903f
C4166 a_n971_45724# a_n1099_45572# 0.508925f
C4167 a_n97_42460# a_15764_42576# 0.174403f
C4168 a_n2661_43922# VDD 0.611934f
C4169 a_13635_43156# a_13460_43230# 0.234322f
C4170 a_16327_47482# a_3357_43084# 0.114502f
C4171 a_3483_46348# a_10903_43370# 0.404121f
C4172 a_8016_46348# a_8349_46414# 0.232167f
C4173 a_n3674_39304# a_n3565_39304# 0.128699f
C4174 a_3080_42308# C2_P_btm 0.108823f
C4175 a_n2104_42282# a_n3674_38216# 0.155459f
C4176 a_n447_43370# VDD 0.204801f
C4177 a_1799_45572# VDD 0.381212f
C4178 a_3090_45724# a_3537_45260# 0.198803f
C4179 a_1467_44172# a_1756_43548# 0.100052f
C4180 a_18189_46348# VDD 0.211855f
C4181 en_comp a_n1794_35242# 2.31448f
C4182 a_12549_44172# a_19862_44208# 0.262561f
C4183 a_n2956_38216# a_n2810_45028# 5.73989f
C4184 a_n863_45724# a_n1059_45260# 0.162875f
C4185 a_11599_46634# a_n743_46660# 0.248412f
C4186 a_19787_47423# a_19594_46812# 0.108653f
C4187 a_n3690_39616# VDD 0.358567f
C4188 a_7754_38470# a_8530_39574# 0.143675f
C4189 a_9313_45822# a_2107_46812# 0.298046f
C4190 a_17478_45572# VDD 0.411207f
C4191 a_2680_45002# a_3065_45002# 0.13328f
C4192 a_10227_46804# a_13635_43156# 0.320228f
C4193 a_3483_46348# a_14955_43940# 0.242667f
C4194 a_10428_46928# a_10623_46897# 0.21686f
C4195 a_4883_46098# a_3483_46348# 0.813604f
C4196 a_13507_46334# a_4185_45028# 0.479559f
C4197 a_n452_44636# VDD 0.112149f
C4198 a_n3674_39768# a_n4064_40160# 0.139482f
C4199 a_15743_43084# a_19339_43156# 0.128224f
C4200 a_3232_43370# a_n2661_42834# 0.127534f
C4201 a_20935_43940# VDD 0.184334f
C4202 a_2747_46873# VDD 0.626468f
C4203 a_12465_44636# CLK 0.795478f
C4204 a_n913_45002# a_2982_43646# 0.498826f
C4205 a_n699_43396# a_2998_44172# 0.127437f
C4206 a_20202_43084# a_10193_42453# 0.296862f
C4207 a_2063_45854# a_8975_43940# 0.149528f
C4208 a_n1641_43230# VDD 0.203991f
C4209 a_20202_43084# VDD 0.987622f
C4210 a_2324_44458# a_5205_44484# 0.523531f
C4211 a_10903_43370# a_11963_45334# 0.209081f
C4212 a_9290_44172# a_9482_43914# 0.135239f
C4213 a_16327_47482# a_18597_46090# 1.28053f
C4214 a_17591_47464# a_10227_46804# 0.292864f
C4215 a_11967_42832# a_18083_42858# 0.472348f
C4216 a_7499_43078# a_n2293_42834# 0.352878f
C4217 C0_dummy_N_btm C7_N_btm 0.119061f
C4218 a_584_46384# a_376_46348# 0.232754f
C4219 C0_N_btm C6_N_btm 0.139059f
C4220 C1_N_btm C5_N_btm 0.127408f
C4221 C2_N_btm C4_N_btm 7.72909f
C4222 C3_P_btm VDD 0.26836f
C4223 a_n237_47217# a_167_45260# 0.280171f
C4224 a_5837_45028# VDD 0.191549f
C4225 a_n443_42852# a_n2661_42282# 0.133617f
C4226 a_15227_44166# a_12741_44636# 0.250453f
C4227 a_2063_45854# a_10193_42453# 0.114552f
C4228 a_3090_45724# a_n2293_46098# 0.642755f
C4229 a_n809_44244# VDD 0.47719f
C4230 a_18184_42460# a_3422_30871# 0.649102f
C4231 a_11823_42460# a_9145_43396# 0.146085f
C4232 a_2063_45854# VDD 3.60498f
C4233 a_8016_46348# a_8034_45724# 0.254614f
C4234 a_14955_43396# VDD 0.401358f
C4235 a_12469_46902# VDD 0.203316f
C4236 a_n755_45592# a_6123_31319# 0.199766f
C4237 a_2127_44172# a_895_43940# 0.132679f
C4238 a_1414_42308# a_2889_44172# 0.128883f
C4239 a_n443_46116# a_1414_42308# 0.18376f
C4240 a_n1151_42308# a_4915_47217# 0.1374f
C4241 a_n971_45724# a_n1435_47204# 2.23698f
C4242 a_n3420_39616# a_n3420_39072# 0.115485f
C4243 a_14383_46116# VDD 0.132317f
C4244 a_n356_44636# a_5342_30871# 0.133551f
C4245 a_11823_42460# a_n1059_45260# 0.100641f
C4246 a_4791_45118# a_3090_45724# 0.206257f
C4247 a_n1613_43370# a_3699_46634# 0.344308f
C4248 a_5691_45260# a_5837_45028# 0.171361f
C4249 a_16327_47482# a_8049_45260# 0.605463f
C4250 a_11813_46116# a_12156_46660# 0.157972f
C4251 a_n2661_42834# VDD 1.00348f
C4252 a_12545_42858# a_5534_30871# 0.17182f
C4253 a_n357_42282# a_8685_43396# 0.319118f
C4254 a_15227_44166# a_16375_45002# 0.117865f
C4255 a_584_46384# a_3232_43370# 0.277433f
C4256 a_n4318_38216# a_n3674_38216# 2.91597f
C4257 a_n1352_43396# VDD 0.288329f
C4258 a_10903_43370# a_13249_42308# 0.211356f
C4259 a_12594_46348# a_13527_45546# 0.100424f
C4260 a_6755_46942# a_14537_43396# 0.120241f
C4261 a_n2293_42282# VDD 0.464485f
C4262 a_17715_44484# VDD 0.526119f
C4263 a_742_44458# a_1847_42826# 0.372436f
C4264 a_9313_44734# a_15743_43084# 1.48048f
C4265 a_n3674_39768# a_n4318_39304# 2.75695f
C4266 a_10193_42453# a_15861_45028# 0.432483f
C4267 a_n863_45724# a_n2017_45002# 0.111825f
C4268 a_n3565_39590# VDD 1.26315f
C4269 a_7754_40130# a_11206_38545# 0.736866f
C4270 a_13507_46334# a_5807_45002# 1.64614f
C4271 a_15861_45028# VDD 0.690795f
C4272 a_2382_45260# a_3065_45002# 0.632538f
C4273 a_10227_46804# a_12895_43230# 0.152365f
C4274 a_3483_46348# a_13483_43940# 0.194464f
C4275 a_n971_45724# a_526_44458# 0.21769f
C4276 a_10428_46928# a_10467_46802# 0.820079f
C4277 a_n1151_42308# a_10809_44734# 0.334692f
C4278 a_12861_44030# a_10903_43370# 0.378457f
C4279 a_n1352_44484# VDD 0.276725f
C4280 a_n4318_39768# a_n4064_40160# 0.293052f
C4281 a_626_44172# a_n356_44636# 0.249281f
C4282 a_15227_44166# a_18985_46122# 0.287996f
C4283 a_n2438_43548# a_n755_45592# 0.213107f
C4284 a_4190_30871# a_19332_42282# 0.154377f
C4285 a_20623_43914# VDD 0.258478f
C4286 a_5111_44636# a_n97_42460# 0.211832f
C4287 a_16327_47482# a_20193_45348# 0.359904f
C4288 a_4791_45118# a_4743_44484# 0.165321f
C4289 a_n1423_42826# VDD 0.211036f
C4290 a_22365_46825# VDD 0.193587f
C4291 a_9885_42558# VDD 0.18767f
C4292 a_2063_45854# a_9804_47204# 0.249806f
C4293 a_n1151_42308# a_n881_46662# 1.41446f
C4294 w_1575_34946# EN_VIN_BSTR_P 3.97882f
C4295 a_8696_44636# a_3232_43370# 0.169534f
C4296 C0_dummy_N_btm C6_N_btm 0.1194f
C4297 C2_N_btm C3_N_btm 5.99608f
C4298 C0_N_btm C5_N_btm 0.138093f
C4299 C1_N_btm C4_N_btm 0.128167f
C4300 C4_P_btm VDD 0.265463f
C4301 a_n746_45260# a_167_45260# 0.234425f
C4302 a_5093_45028# VDD 0.168437f
C4303 a_3080_42308# a_n2293_42282# 0.122474f
C4304 a_19692_46634# a_20202_43084# 0.172738f
C4305 a_n2661_46098# a_n2956_38680# 0.123968f
C4306 a_n1549_44318# VDD 0.200608f
C4307 a_584_46384# VDD 2.50905f
C4308 a_327_47204# DATA[0] 0.353891f
C4309 a_15095_43370# VDD 0.169652f
C4310 COMP_P a_5742_30871# 0.109332f
C4311 a_n2840_43914# a_n4318_39768# 0.170372f
C4312 a_11901_46660# VDD 0.57548f
C4313 a_2127_44172# a_2479_44172# 0.168988f
C4314 a_453_43940# a_895_43940# 0.420851f
C4315 a_1414_42308# a_2675_43914# 0.305556f
C4316 a_3815_47204# a_4007_47204# 0.224415f
C4317 a_14097_32519# VDD 0.284675f
C4318 a_22537_39537# a_22629_38406# 0.198762f
C4319 a_5807_45002# a_n743_46660# 0.669712f
C4320 a_10227_46804# a_10150_46912# 0.236747f
C4321 a_n1613_43370# a_2959_46660# 0.187029f
C4322 a_21513_45002# a_21359_45002# 0.289039f
C4323 a_413_45260# a_n2661_43370# 1.31746f
C4324 a_n746_45260# a_n863_45724# 0.664707f
C4325 a_5343_44458# a_6298_44484# 0.128602f
C4326 a_4223_44672# a_5883_43914# 0.967973f
C4327 a_9290_44172# a_10835_43094# 0.172486f
C4328 a_413_45260# a_2998_44172# 0.161528f
C4329 a_3357_43084# a_3499_42826# 0.134316f
C4330 a_7920_46348# a_8016_46348# 0.318386f
C4331 a_n1177_43370# VDD 0.354704f
C4332 a_3090_45724# a_3065_45002# 0.475346f
C4333 a_526_44458# a_2711_45572# 0.392618f
C4334 a_19332_42282# a_19511_42282# 0.174683f
C4335 a_22959_42860# VDD 0.30747f
C4336 a_17583_46090# VDD 0.23578f
C4337 a_9028_43914# a_9165_43940# 0.126609f
C4338 a_10193_42453# a_8696_44636# 0.225102f
C4339 a_7754_40130# VDAC_P 0.334598f
C4340 VDAC_Pi a_6886_37412# 0.259481f
C4341 a_n4334_39616# VDD 0.385881f
C4342 a_8696_44636# VDD 1.12228f
C4343 a_10227_46804# a_13113_42826# 0.159547f
C4344 a_10150_46912# a_10467_46802# 0.102355f
C4345 a_n1177_44458# VDD 0.347966f
C4346 a_13249_42308# a_13483_43940# 0.193724f
C4347 a_11827_44484# a_22223_45036# 0.179208f
C4348 a_15227_44166# a_18819_46122# 0.288885f
C4349 a_20365_43914# VDD 0.261299f
C4350 a_n2312_40392# CLK_DATA 0.213071f
C4351 a_16327_47482# a_11691_44458# 0.536141f
C4352 a_n1991_42858# VDD 0.575656f
C4353 a_18494_42460# a_743_42282# 0.476713f
C4354 a_20820_30879# C7_N_btm 0.184297f
C4355 a_10809_44734# a_413_45260# 0.333257f
C4356 a_2324_44458# a_6171_45002# 2.73828f
C4357 a_5742_30871# C6_N_btm 0.170624f
C4358 a_n4209_38216# a_n3565_38216# 6.80743f
C4359 a_16327_47482# a_18479_47436# 0.723416f
C4360 a_n1151_42308# a_n1613_43370# 1.19311f
C4361 a_7227_45028# VDD 0.501104f
C4362 w_1575_34946# a_n1057_35174# 37.7491f
C4363 a_16327_47482# a_4190_30871# 0.335014f
C4364 EN_VIN_BSTR_P VIN_P 1.41696f
C4365 C1_N_btm C3_N_btm 8.06688f
C4366 C0_dummy_N_btm C5_N_btm 0.11375f
C4367 C0_N_btm C4_N_btm 0.138331f
C4368 C5_P_btm VDD 0.267489f
C4369 a_n237_47217# a_1823_45246# 0.370766f
C4370 a_5009_45028# VDD 0.151712f
C4371 a_3422_30871# a_4958_30871# 0.101017f
C4372 a_3537_45260# a_4223_44672# 0.1907f
C4373 a_n1331_43914# VDD 0.203823f
C4374 a_3422_30871# VCM 1.12142f
C4375 a_n2312_38680# a_n2302_38778# 0.161815f
C4376 SMPL_ON_P VIN_P 0.546737f
C4377 a_n785_47204# DATA[0] 0.598846f
C4378 a_14205_43396# VDD 0.311811f
C4379 a_11813_46116# VDD 0.434656f
C4380 a_1414_42308# a_895_43940# 0.208524f
C4381 a_18189_46348# a_16147_45260# 0.129202f
C4382 a_1169_39587# a_1666_39587# 0.105143f
C4383 a_3785_47178# a_4007_47204# 0.106797f
C4384 a_n1151_42308# a_4791_45118# 1.16458f
C4385 a_2063_45854# a_6151_47436# 0.448977f
C4386 a_22400_42852# VDD 0.888056f
C4387 a_20512_43084# a_15743_43084# 0.761578f
C4388 a_13661_43548# a_19319_43548# 0.189089f
C4389 VDAC_N EN_VIN_BSTR_N 0.341739f
C4390 a_10227_46804# a_9863_46634# 0.278164f
C4391 a_22581_37893# a_22629_37990# 0.333805f
C4392 a_n1613_43370# a_3177_46902# 0.209276f
C4393 a_n967_45348# VDD 0.556063f
C4394 en_comp RST_Z 4.35406f
C4395 a_4927_45028# a_5093_45028# 0.143754f
C4396 a_3537_45260# a_n2293_42834# 0.195818f
C4397 a_n971_45724# a_n863_45724# 0.199707f
C4398 a_3090_45724# a_15368_46634# 0.440843f
C4399 a_n97_42460# a_14113_42308# 0.356407f
C4400 a_12545_42858# a_13460_43230# 0.118423f
C4401 a_12379_42858# a_5534_30871# 0.128429f
C4402 a_7499_43078# a_n97_42460# 0.212833f
C4403 a_413_45260# a_2889_44172# 0.127135f
C4404 a_20820_30879# a_10809_44734# 0.234047f
C4405 a_n443_46116# a_413_45260# 0.369976f
C4406 a_4646_46812# a_7227_45028# 0.305597f
C4407 a_n1917_43396# VDD 0.204644f
C4408 a_n1059_45260# a_17499_43370# 0.385066f
C4409 a_19279_43940# a_18579_44172# 0.372064f
C4410 a_2324_44458# a_8746_45002# 0.34917f
C4411 a_22223_42860# VDD 0.250812f
C4412 a_4958_30871# a_7174_31319# 0.107892f
C4413 a_15682_46116# VDD 1.25004f
C4414 a_n2293_46098# a_4223_44672# 0.422068f
C4415 a_n2109_47186# a_5257_43370# 0.153164f
C4416 a_7754_40130# a_8912_37509# 1.81084f
C4417 a_n443_46116# a_2609_46660# 0.349838f
C4418 VDAC_Pi a_5700_37509# 2.20213f
C4419 a_n4209_39590# VDD 2.06918f
C4420 a_18494_42460# a_13258_32519# 0.298557f
C4421 a_16680_45572# VDD 0.275078f
C4422 a_n443_42852# a_n356_44636# 0.262144f
C4423 a_10150_46912# a_10428_46928# 0.118759f
C4424 a_n2293_46634# a_13059_46348# 0.207934f
C4425 a_n1917_44484# VDD 0.186988f
C4426 a_18494_42460# a_20193_45348# 0.116597f
C4427 a_20269_44172# VDD 0.169009f
C4428 a_n4318_40392# a_n4318_39768# 2.73673f
C4429 a_4791_45118# a_4223_44672# 0.399086f
C4430 a_n1613_43370# a_n2293_42834# 0.123758f
C4431 a_n1853_43023# VDD 0.370563f
C4432 a_18184_42460# a_743_42282# 0.126294f
C4433 a_7499_43078# a_10533_42308# 0.225871f
C4434 a_526_44458# a_n2661_45010# 0.703081f
C4435 a_12861_44030# a_12429_44172# 0.108591f
C4436 a_2324_44458# a_3232_43370# 0.410727f
C4437 a_n4209_38216# a_n4334_38304# 0.253307f
C4438 a_12861_44030# a_13507_46334# 0.315418f
C4439 a_5932_42308# VCM 0.146001f
C4440 a_6598_45938# VDD 0.204705f
C4441 a_15493_43396# a_16409_43396# 0.566182f
C4442 w_1575_34946# a_n1696_35090# 0.799782f
C4443 a_4185_45028# a_3422_30871# 0.176529f
C4444 a_n1057_35174# VIN_P 1.547f
C4445 a_11599_46634# a_20107_46660# 0.266678f
C4446 C0_dummy_N_btm C4_N_btm 0.113156f
C4447 C1_N_btm C2_N_btm 5.24136f
C4448 C0_N_btm C3_N_btm 0.409238f
C4449 C6_P_btm VDD 0.210613f
C4450 a_2809_45028# VDD 0.189682f
C4451 a_n1899_43946# VDD 0.475205f
C4452 a_3422_30871# VREF_GND 0.10463f
C4453 a_n237_47217# DATA[1] 0.139838f
C4454 a_n2312_38680# a_n4064_38528# 0.22404f
C4455 a_1431_47204# VDD 0.423871f
C4456 a_8953_45546# a_5066_45546# 0.191859f
C4457 a_14358_43442# VDD 0.170277f
C4458 a_11735_46660# VDD 0.407307f
C4459 a_1414_42308# a_2479_44172# 0.110442f
C4460 a_742_44458# a_1756_43548# 0.152145f
C4461 a_3785_47178# a_3815_47204# 0.270823f
C4462 a_2905_45572# a_n443_46116# 0.14923f
C4463 a_n1605_47204# a_n1435_47204# 0.110832f
C4464 a_15861_45028# a_16147_45260# 0.146279f
C4465 VDAC_P EN_VIN_BSTR_P 0.340512f
C4466 a_5807_45002# a_n1925_46634# 0.933976f
C4467 a_21588_30879# a_22612_30879# 7.53611f
C4468 a_n1613_43370# a_2609_46660# 0.631348f
C4469 en_comp VDD 4.30454f
C4470 a_6755_46942# a_13059_46348# 0.239671f
C4471 a_n971_45724# a_n1079_45724# 0.150623f
C4472 a_n746_45260# a_n2293_45546# 0.404324f
C4473 a_3090_45724# a_14976_45028# 0.730613f
C4474 a_3626_43646# a_5934_30871# 0.192998f
C4475 a_10617_44484# VDD 0.141193f
C4476 a_13113_42826# a_12895_43230# 0.209641f
C4477 a_n2312_39304# a_n2302_39072# 0.130454f
C4478 a_9290_44172# a_10083_42826# 0.136441f
C4479 a_3483_46348# a_9290_44172# 0.207611f
C4480 a_15227_44166# a_13259_45724# 0.916975f
C4481 a_n1699_43638# VDD 0.210236f
C4482 a_n2472_42282# a_n4318_38216# 0.157105f
C4483 a_11967_42832# a_3422_30871# 0.139082f
C4484 a_6755_46942# a_13556_45296# 0.103107f
C4485 a_19321_45002# a_20193_45348# 0.489018f
C4486 a_22165_42308# VDD 0.336187f
C4487 a_2324_44458# VDD 2.73366f
C4488 VDAC_Pi a_5088_37509# 0.391059f
C4489 a_18479_47436# a_19594_46812# 0.108004f
C4490 a_19386_47436# a_13747_46662# 0.145228f
C4491 a_7754_40130# VDAC_N 0.434929f
C4492 a_n971_45724# a_6540_46812# 0.31827f
C4493 a_12861_44030# a_n743_46660# 0.100542f
C4494 a_n2293_43922# COMP_P 0.151768f
C4495 a_16855_45546# VDD 0.339227f
C4496 a_n357_42282# a_5891_43370# 0.304889f
C4497 a_2274_45254# a_2382_45260# 0.130215f
C4498 a_12549_44172# a_17639_46660# 0.129285f
C4499 a_n1699_44726# VDD 0.198612f
C4500 a_n743_46660# a_310_45028# 0.143623f
C4501 a_12465_44636# a_11823_42460# 0.127538f
C4502 a_19862_44208# VDD 0.588967f
C4503 a_4185_45028# a_5932_42308# 0.118319f
C4504 en_comp a_3080_42308# 1.2852f
C4505 a_9290_44172# a_n357_42282# 0.138435f
C4506 a_n2157_42858# VDD 0.424058f
C4507 a_18494_42460# a_4190_30871# 0.242908f
C4508 a_10193_42453# a_9803_42558# 0.20198f
C4509 a_9803_42558# VDD 0.253745f
C4510 a_16327_47482# a_10227_46804# 0.630403f
C4511 a_16763_47508# a_16588_47582# 0.233657f
C4512 a_6667_45809# VDD 0.195842f
C4513 a_3699_46634# a_3524_46660# 0.233657f
C4514 a_n971_45724# a_1823_45246# 0.514159f
C4515 C0_N_btm C2_N_btm 0.827449f
C4516 C7_P_btm VDD 0.121904f
C4517 a_4915_47217# a_11415_45002# 0.134061f
C4518 a_2063_45854# a_7499_43078# 0.478913f
C4519 a_n1761_44111# VDD 0.620042f
C4520 a_9482_43914# a_9672_43914# 0.122568f
C4521 a_1239_47204# VDD 0.278979f
C4522 a_5937_45572# a_5066_45546# 0.419426f
C4523 a_20075_46420# a_19900_46494# 0.233657f
C4524 a_1606_42308# a_6123_31319# 1.43958f
C4525 a_14579_43548# VDD 0.278225f
C4526 a_742_44458# a_1568_43370# 0.525694f
C4527 a_10586_45546# CLK 0.125859f
C4528 a_12839_46116# VDD 0.347766f
C4529 a_8696_44636# a_16147_45260# 0.284694f
C4530 a_n1613_43370# a_2443_46660# 0.917984f
C4531 a_22527_39145# a_22629_37990# 0.172129f
C4532 a_22581_37893# a_22629_38406# 0.236891f
C4533 a_n2956_37592# VDD 1.25966f
C4534 a_15415_45028# a_15595_45028# 0.185422f
C4535 a_n2661_46098# a_n2157_46122# 0.227082f
C4536 a_12379_42858# a_13460_43230# 0.102325f
C4537 a_12545_42858# a_12895_43230# 0.215953f
C4538 a_n2661_43370# a_n2661_43922# 0.13591f
C4539 a_11415_45002# a_10809_44734# 0.140489f
C4540 a_n2267_43396# VDD 0.570924f
C4541 a_5342_30871# a_4958_30871# 10.9366f
C4542 a_n3674_38680# a_n4318_38216# 2.82961f
C4543 a_491_47026# VDD 0.132552f
C4544 a_21671_42860# VDD 0.229963f
C4545 a_5342_30871# VCM 0.325566f
C4546 a_14840_46494# VDD 0.275785f
C4547 a_n863_45724# a_n2661_45010# 0.345234f
C4548 a_n443_46116# a_n97_42460# 0.131756f
C4549 a_n2293_45546# a_n2293_45010# 0.257189f
C4550 VDAC_Pi a_4338_37500# 1.92369f
C4551 a_18597_46090# a_13747_46662# 0.391702f
C4552 a_18479_47436# a_19321_45002# 0.262984f
C4553 a_7754_39964# a_5088_37509# 0.392826f
C4554 a_n443_46116# a_n2661_46098# 0.198865f
C4555 a_16115_45572# VDD 0.194492f
C4556 a_n1613_43370# a_n1076_43230# 0.224215f
C4557 a_2711_45572# a_14539_43914# 0.199754f
C4558 a_10227_46804# a_12379_42858# 0.298444f
C4559 a_9863_46634# a_10150_46912# 0.233657f
C4560 a_13747_46662# a_19123_46287# 0.191545f
C4561 a_n2267_44484# VDD 0.289888f
C4562 a_n743_46660# a_n1099_45572# 0.108295f
C4563 a_15227_44166# a_17715_44484# 0.385336f
C4564 a_19478_44306# VDD 0.127794f
C4565 a_3537_45260# a_n97_42460# 0.74108f
C4566 a_n2312_39304# VDD 0.587668f
C4567 a_n357_42282# a_16795_42852# 0.180926f
C4568 a_15227_44166# a_15861_45028# 0.208121f
C4569 a_1823_45246# a_2711_45572# 0.262616f
C4570 a_n2472_42826# VDD 0.229608f
C4571 a_n1794_35242# a_n4315_30879# 0.129428f
C4572 a_18184_42460# a_4190_30871# 0.630738f
C4573 a_11599_46634# a_18597_46090# 0.191253f
C4574 a_9223_42460# VDD 0.205797f
C4575 a_16327_47482# a_17591_47464# 0.339529f
C4576 a_6511_45714# VDD 0.405279f
C4577 a_n97_42460# a_1049_43396# 0.195034f
C4578 a_13507_46334# a_15743_43084# 0.158635f
C4579 a_13747_46662# a_6755_46942# 0.316914f
C4580 a_n1550_35608# VIN_P 0.37444f
C4581 C8_P_btm VDD 0.19922f
C4582 C0_dummy_N_btm C2_N_btm 7.14548f
C4583 C0_N_btm C1_N_btm 11.2332f
C4584 SMPL_ON_N a_n1794_35242# 0.150516f
C4585 a_13556_45296# a_11691_44458# 0.399095f
C4586 a_16388_46812# a_765_45546# 0.164902f
C4587 a_13747_46662# a_8049_45260# 0.208778f
C4588 a_6151_47436# a_6598_45938# 0.173467f
C4589 w_1575_34946# a_3422_30871# 1.88476f
C4590 a_n2438_43548# a_526_44458# 0.107408f
C4591 a_3877_44458# a_2324_44458# 0.153319f
C4592 a_n881_46662# a_13259_45724# 0.507296f
C4593 a_n2065_43946# VDD 0.4213f
C4594 a_12281_43396# a_12563_42308# 0.173003f
C4595 a_10440_44484# a_10617_44484# 0.134298f
C4596 a_1209_47178# VDD 0.38145f
C4597 a_8199_44636# a_5066_45546# 0.178583f
C4598 a_13667_43396# VDD 0.402378f
C4599 a_10768_47026# VDD 0.132317f
C4600 a_644_44056# a_895_43940# 0.106452f
C4601 a_1414_42308# a_453_43940# 0.248504f
C4602 a_5891_43370# a_9127_43156# 0.457718f
C4603 a_n1613_43370# a_n2661_46098# 1.40554f
C4604 a_22589_40055# a_22629_37990# 0.234448f
C4605 a_11599_46634# a_6755_46942# 0.321942f
C4606 a_n2810_45028# VDD 0.526631f
C4607 a_n2293_46098# a_n97_42460# 0.333817f
C4608 a_n357_42282# a_3422_30871# 0.122733f
C4609 a_15009_46634# a_3090_45724# 0.154981f
C4610 a_11599_46634# a_8049_45260# 0.14064f
C4611 a_n2497_47436# a_n755_45592# 0.45034f
C4612 a_3422_30871# CAL_N 0.236929f
C4613 a_3626_43646# a_6123_31319# 0.109715f
C4614 a_2982_43646# a_5934_30871# 0.178f
C4615 a_12545_42858# a_13113_42826# 0.178024f
C4616 a_n2661_43370# a_n2661_42834# 0.306215f
C4617 a_n881_46662# a_17478_45572# 0.11503f
C4618 a_4646_46812# a_6511_45714# 0.421269f
C4619 a_n2129_43609# VDD 0.400674f
C4620 a_14539_43914# a_15682_43940# 0.161926f
C4621 a_n2661_42834# a_2998_44172# 0.790177f
C4622 a_12594_46348# a_11962_45724# 0.177228f
C4623 a_19321_45002# a_19113_45348# 0.147788f
C4624 a_10903_43370# a_11823_42460# 1.16382f
C4625 a_21195_42852# VDD 0.285496f
C4626 a_n2017_45002# a_n1794_35242# 0.111641f
C4627 a_15015_46420# VDD 0.337162f
C4628 a_n967_45348# a_n961_42308# 0.174237f
C4629 a_9290_44172# CLK 0.151406f
C4630 a_7499_43078# a_8696_44636# 0.155392f
C4631 VDAC_Pi a_3726_37500# 1.17174f
C4632 a_n2302_40160# VDD 0.428934f
C4633 a_18597_46090# a_13661_43548# 0.266647f
C4634 a_7754_38636# a_7754_38470# 0.296258f
C4635 a_n2810_45028# a_n2302_37690# 0.162246f
C4636 a_16333_45814# VDD 0.201203f
C4637 a_n1613_43370# a_n901_43156# 0.281398f
C4638 a_13661_43548# a_743_42282# 0.132115f
C4639 a_2711_45572# a_16112_44458# 0.183744f
C4640 a_2063_45854# a_10809_44734# 0.169005f
C4641 a_7411_46660# a_6755_46942# 0.265786f
C4642 a_n2129_44697# VDD 1.4165f
C4643 a_3232_43370# a_3363_44484# 0.103472f
C4644 a_21101_45002# a_21359_45002# 0.22264f
C4645 a_15493_43396# VDD 2.34659f
C4646 a_4190_30871# a_17303_42282# 0.279034f
C4647 a_n2312_40392# VDD 0.947797f
C4648 a_5257_43370# a_3357_43084# 0.894879f
C4649 a_15227_44166# a_8696_44636# 0.203885f
C4650 a_16327_47482# a_11827_44484# 0.107078f
C4651 a_n2840_42826# VDD 0.302305f
C4652 a_9290_44172# a_10951_45334# 0.136064f
C4653 a_3483_46348# a_1423_45028# 0.110369f
C4654 a_n1613_43370# a_n984_44318# 0.245331f
C4655 a_8791_42308# VDD 0.226318f
C4656 a_2063_45854# a_n881_46662# 0.612456f
C4657 a_16327_47482# a_16588_47582# 0.276601f
C4658 a_21381_43940# a_2982_43646# 0.236232f
C4659 a_6472_45840# VDD 0.257073f
C4660 a_10809_44734# a_n2661_42834# 0.14417f
C4661 a_20273_45572# a_3357_43084# 0.358383f
C4662 C9_P_btm VDD 0.345685f
C4663 C0_dummy_N_btm C1_N_btm 1.24905f
C4664 a_n2661_42282# a_5379_42460# 0.121051f
C4665 a_9482_43914# a_11691_44458# 0.616964f
C4666 a_16388_46812# a_17339_46660# 0.24887f
C4667 a_6151_47436# a_6667_45809# 0.1609f
C4668 a_12891_46348# a_12638_46436# 0.13727f
C4669 a_n2472_43914# VDD 0.236691f
C4670 a_1307_43914# a_3499_42826# 0.532672f
C4671 a_5883_43914# a_n2661_42834# 0.106812f
C4672 a_327_47204# VDD 0.367528f
C4673 a_n971_45724# DATA[0] 0.213213f
C4674 a_11453_44696# a_6171_45002# 1.39146f
C4675 a_3823_42558# a_3905_42558# 0.171361f
C4676 a_10695_43548# VDD 0.201247f
C4677 a_n1613_43370# a_n2661_43922# 0.113996f
C4678 a_584_46384# a_2998_44172# 0.181241f
C4679 a_18707_42852# VDD 0.132317f
C4680 a_2063_45854# a_n443_46116# 0.177177f
C4681 a_n3565_39590# a_n4209_39304# 5.4667f
C4682 a_22527_39145# a_22629_38406# 0.123152f
C4683 a_n1761_44111# a_n473_42460# 0.110251f
C4684 a_n745_45366# VDD 0.20887f
C4685 a_2982_43646# a_5649_42852# 0.205161f
C4686 a_12379_42858# a_12895_43230# 0.109156f
C4687 a_n699_43396# a_4743_44484# 0.235328f
C4688 a_4223_44672# a_5343_44458# 0.229803f
C4689 a_18479_45785# a_15493_43396# 0.235084f
C4690 a_413_45260# a_2127_44172# 0.104737f
C4691 a_n881_46662# a_15861_45028# 0.153795f
C4692 a_4646_46812# a_6472_45840# 0.129446f
C4693 a_n2433_43396# VDD 0.416276f
C4694 a_17517_44484# a_22591_44484# 0.196232f
C4695 a_1983_46706# VDD 0.119964f
C4696 a_2324_44458# a_9049_44484# 0.102942f
C4697 a_21356_42826# VDD 0.225688f
C4698 a_14275_46494# VDD 0.196859f
C4699 a_15493_43396# a_14021_43940# 0.139192f
C4700 a_n4064_40160# VDD 2.37273f
C4701 a_12465_44636# a_768_44030# 0.120859f
C4702 a_10227_46804# a_19321_45002# 0.111029f
C4703 a_18780_47178# a_13661_43548# 0.153988f
C4704 VDAC_Ni a_3754_38470# 0.911632f
C4705 a_n2810_45028# a_n4064_37440# 0.22413f
C4706 a_15765_45572# VDD 0.249471f
C4707 a_n2956_37592# a_n2946_37690# 0.148852f
C4708 a_19319_43548# a_19268_43646# 0.17076f
C4709 a_6293_42852# a_6452_43396# 0.157972f
C4710 a_7287_43370# a_7112_43396# 0.234322f
C4711 a_n1613_43370# a_n1641_43230# 0.152896f
C4712 a_8696_44636# a_n2661_43370# 0.674122f
C4713 a_10227_46804# a_10922_42852# 0.159426f
C4714 a_n2433_44484# VDD 0.40658f
C4715 a_n2293_42834# a_5343_44458# 0.165923f
C4716 a_768_44030# a_2711_45572# 0.529995f
C4717 a_22959_46660# a_21076_30879# 0.165603f
C4718 a_19328_44172# VDD 0.263964f
C4719 a_4190_30871# a_4958_30871# 11.510201f
C4720 a_22959_47212# VDD 0.245964f
C4721 a_n913_45002# a_4905_42826# 0.101072f
C4722 a_n699_43396# a_1414_42308# 0.104607f
C4723 a_5066_45546# a_8034_45724# 0.242476f
C4724 a_4190_30871# VCM 1.23535f
C4725 a_11551_42558# a_11633_42558# 0.171361f
C4726 a_n357_42282# a_20712_42282# 0.173926f
C4727 a_10057_43914# a_10695_43548# 0.148476f
C4728 a_3090_45724# a_4223_44672# 0.269823f
C4729 a_8199_44636# a_9482_43914# 0.276776f
C4730 a_9290_44172# a_10775_45002# 0.215292f
C4731 a_n1613_43370# a_n809_44244# 0.291484f
C4732 a_8685_42308# VDD 0.286875f
C4733 a_584_46384# a_n881_46662# 0.286501f
C4734 a_16327_47482# a_16763_47508# 0.338544f
C4735 a_6194_45824# VDD 0.274689f
C4736 a_20107_45572# a_3357_43084# 0.308463f
C4737 a_16327_47482# a_16823_43084# 0.535969f
C4738 a_526_44458# a_5891_43370# 1.12739f
C4739 a_3090_45724# a_15493_43940# 0.255251f
C4740 a_2609_46660# a_3524_46660# 0.118759f
C4741 a_5807_45002# a_6755_46942# 1.47519f
C4742 a_2063_45854# a_n2293_46098# 0.994164f
C4743 C10_P_btm VDD 2.40001f
C4744 a_10227_46804# a_13059_46348# 0.656528f
C4745 C0_dummy_N_btm C0_N_btm 7.97415f
C4746 a_3232_43370# a_n2661_44458# 0.468391f
C4747 a_5807_45002# a_8049_45260# 1.37423f
C4748 a_6151_47436# a_6511_45714# 0.3215f
C4749 a_n4318_38680# a_n3674_38680# 3.04229f
C4750 a_n2840_43914# VDD 0.304745f
C4751 a_n2312_38680# a_n3565_38502# 0.134976f
C4752 a_18184_42460# a_18579_44172# 0.161593f
C4753 a_n755_45592# a_743_42282# 0.160592f
C4754 a_n785_47204# VDD 0.452945f
C4755 a_9290_44172# a_526_44458# 0.200352f
C4756 a_18985_46122# a_19900_46494# 0.118759f
C4757 a_11453_44696# a_3232_43370# 0.132496f
C4758 a_9803_43646# VDD 0.261557f
C4759 a_1467_44172# a_1414_42308# 0.335735f
C4760 a_1115_44172# a_453_43940# 0.150214f
C4761 a_16327_47482# a_19279_43940# 0.446333f
C4762 a_n1613_43370# a_n2661_42834# 0.112184f
C4763 a_10809_44734# a_8696_44636# 0.117876f
C4764 a_584_46384# a_n443_46116# 0.496286f
C4765 a_n1794_35242# a_18194_35068# 0.466445f
C4766 a_10193_42453# a_n913_45002# 0.562004f
C4767 a_n1613_43370# a_n1352_43396# 0.244933f
C4768 a_n755_45592# a_626_44172# 0.100613f
C4769 a_22537_40625# a_22629_37990# 0.130478f
C4770 a_22589_40055# a_22629_38406# 0.1922f
C4771 a_3626_43646# a_4361_42308# 5.20633f
C4772 a_n913_45002# VDD 9.190901f
C4773 a_n2661_46098# a_n2840_46090# 0.170439f
C4774 a_n2293_46634# a_3483_46348# 0.157275f
C4775 a_n97_42460# a_13575_42558# 0.179828f
C4776 a_2982_43646# a_6123_31319# 0.163265f
C4777 a_12089_42308# a_12545_42858# 0.261463f
C4778 a_3422_30871# VDAC_P 0.476125f
C4779 a_584_46384# a_3537_45260# 0.108506f
C4780 a_n881_46662# a_8696_44636# 0.178516f
C4781 a_n2840_42282# a_n3674_38680# 0.154001f
C4782 a_n4318_39304# VDD 0.643395f
C4783 a_22400_42852# COMP_P 0.595635f
C4784 a_2107_46812# VDD 0.350275f
C4785 a_17517_44484# a_22485_44484# 0.110643f
C4786 a_n356_44636# a_n2661_42282# 2.54767f
C4787 a_3090_45724# a_413_45260# 0.135828f
C4788 a_13661_43548# a_11691_44458# 0.263889f
C4789 a_n1613_43370# a_n1352_44484# 0.232498f
C4790 a_10903_43370# a_11962_45724# 0.357882f
C4791 a_20922_43172# VDD 0.192467f
C4792 a_14493_46090# VDD 0.203567f
C4793 a_n2017_45002# a_n3674_37592# 0.241068f
C4794 a_2479_44172# a_n97_42460# 0.196935f
C4795 a_584_46384# a_1049_43396# 0.148494f
C4796 a_n4334_40480# VDD 0.390668f
C4797 a_15903_45785# VDD 0.291109f
C4798 a_n2956_37592# a_n3420_37440# 0.233174f
C4799 a_n1613_43370# a_n1423_42826# 0.15981f
C4800 a_13661_43548# a_4190_30871# 0.147163f
C4801 a_3483_46348# a_9672_43914# 0.125466f
C4802 a_10227_46804# a_10991_42826# 0.152133f
C4803 a_n2661_44458# VDD 1.06317f
C4804 a_10193_42453# a_18451_43940# 0.20167f
C4805 a_4185_45028# a_4190_30871# 0.16524f
C4806 a_21005_45260# a_21101_45002# 0.419086f
C4807 a_15227_44166# a_2324_44458# 0.190521f
C4808 a_12549_44172# a_2711_45572# 2.05236f
C4809 a_18451_43940# VDD 0.172318f
C4810 a_11453_44696# VDD 3.75355f
C4811 SMPL_ON_N RST_Z 2.43362f
C4812 a_4190_30871# VREF_GND 0.105109f
C4813 a_17364_32525# VDD 0.511443f
C4814 a_7499_43078# a_9803_42558# 0.158876f
C4815 a_n1613_43370# a_n1549_44318# 0.16289f
C4816 a_15507_47210# a_10227_46804# 0.23187f
C4817 a_8325_42308# VDD 0.313956f
C4818 a_15673_47210# a_16588_47582# 0.125324f
C4819 a_n3420_38528# a_n4064_37984# 7.35343f
C4820 a_16327_47482# a_16023_47582# 0.159305f
C4821 a_5907_45546# VDD 0.390381f
C4822 a_21753_35634# VDD 0.527767f
C4823 a_3177_46902# a_2959_46660# 0.209641f
C4824 a_2443_46660# a_3524_46660# 0.102325f
C4825 a_11599_46634# a_765_45546# 0.332797f
C4826 a_5257_43370# a_5937_45572# 0.262028f
C4827 a_18597_46090# a_n357_42282# 0.250702f
C4828 a_n3674_39304# a_n3674_38680# 0.17962f
C4829 a_19237_31679# VDD 0.746417f
C4830 a_19778_44110# a_18579_44172# 0.268475f
C4831 a_n23_47502# VDD 0.152616f
C4832 a_19553_46090# a_19335_46494# 0.209641f
C4833 a_18819_46122# a_19900_46494# 0.102355f
C4834 a_9145_43396# VDD 2.43736f
C4835 a_5267_42460# a_5379_42460# 0.156424f
C4836 a_1115_44172# a_1414_42308# 0.134389f
C4837 a_n913_45002# a_2075_43172# 0.175893f
C4838 a_16327_47482# a_20766_44850# 0.17113f
C4839 a_n356_45724# a_n23_45546# 0.360492f
C4840 a_21076_30879# a_413_45260# 0.141502f
C4841 a_n2661_45546# a_2711_45572# 0.359276f
C4842 a_n755_45592# a_1609_45822# 0.12055f
C4843 a_n1741_47186# a_9313_45822# 0.102019f
C4844 a_5891_43370# a_8037_42858# 0.12253f
C4845 a_10193_42453# a_n1059_45260# 0.440111f
C4846 a_n1613_43370# a_n1177_43370# 0.325171f
C4847 a_n357_42282# a_626_44172# 0.551369f
C4848 a_22581_37893# a_22537_39537# 1.00904f
C4849 a_22613_38993# a_22889_38993# 0.237336f
C4850 a_7754_39632# VDD 0.205733f
C4851 a_n1059_45260# VDD 4.75361f
C4852 en_comp a_n2661_43370# 0.164814f
C4853 a_n2312_39304# a_n2956_39304# 6.38528f
C4854 a_12379_42858# a_12545_42858# 0.810394f
C4855 a_413_45260# a_1414_42308# 0.12534f
C4856 a_4223_44672# a_n699_43396# 0.217586f
C4857 a_n2312_39304# a_n3565_39304# 0.104981f
C4858 a_3483_46348# a_8953_45546# 0.133493f
C4859 a_n2840_43370# VDD 0.246858f
C4860 a_10193_42453# a_19987_42826# 0.164153f
C4861 a_n1059_45260# a_16137_43396# 0.438785f
C4862 a_948_46660# VDD 0.278482f
C4863 a_20679_44626# a_19279_43940# 0.279785f
C4864 a_20835_44721# a_20766_44850# 0.209641f
C4865 a_5807_45002# a_11691_44458# 0.117249f
C4866 a_n1613_43370# a_n1177_44458# 0.332209f
C4867 a_18057_42282# a_18214_42558# 0.18824f
C4868 a_19987_42826# VDD 0.588466f
C4869 en_comp COMP_P 1.91962f
C4870 a_15493_43940# a_22959_43948# 0.182001f
C4871 a_13925_46122# VDD 0.251868f
C4872 a_10227_46804# a_13747_46662# 0.16398f
C4873 a_n4315_30879# VDD 4.0486f
C4874 a_13258_32519# VIN_N 0.143165f
C4875 a_15599_45572# VDD 0.390565f
C4876 a_8667_46634# a_8492_46660# 0.233657f
C4877 a_n3674_39304# a_n4318_38680# 2.92578f
C4878 a_n4318_40392# VDD 0.573389f
C4879 a_10193_42453# a_18326_43940# 0.130866f
C4880 a_12741_44636# a_22959_46660# 0.17409f
C4881 a_20820_30879# a_21076_30879# 8.6867f
C4882 a_18326_43940# VDD 0.129408f
C4883 a_n2293_42282# a_n3674_38216# 0.111055f
C4884 SMPL_ON_N VDD 0.497819f
C4885 a_22959_43396# VDD 0.303237f
C4886 a_1606_42308# a_7174_31319# 2.41314f
C4887 a_10057_43914# a_9145_43396# 0.121499f
C4888 a_n1613_43370# a_n1331_43914# 0.16678f
C4889 a_8270_45546# a_8975_43940# 0.207334f
C4890 a_8016_46348# a_9482_43914# 0.293982f
C4891 a_7227_45028# a_7230_45938# 0.170618f
C4892 a_13059_46348# a_11827_44484# 0.495367f
C4893 a_11599_46634# a_10227_46804# 0.60865f
C4894 a_2112_39137# a_2113_38308# 0.478223f
C4895 a_16241_47178# a_16023_47582# 0.209641f
C4896 a_5263_45724# VDD 0.202719f
C4897 a_19998_35138# VDD 0.320029f
C4898 a_2609_46660# a_2959_46660# 0.216095f
C4899 C3_P_btm C3_N_btm 2.90911f
C4900 a_11599_46634# a_17339_46660# 0.131185f
C4901 a_413_45260# a_n699_43396# 0.100762f
C4902 a_4791_45118# a_7227_45028# 0.288276f
C4903 a_6151_47436# a_6194_45824# 0.227219f
C4904 a_22959_44484# VDD 0.303517f
C4905 a_18494_42460# a_19279_43940# 0.137363f
C4906 a_n237_47217# VDD 4.05131f
C4907 a_n356_44636# a_n23_44458# 0.220577f
C4908 a_18985_46122# a_19335_46494# 0.210876f
C4909 a_n1613_43370# a_n967_45348# 0.213625f
C4910 a_1606_42308# a_5932_42308# 0.111585f
C4911 a_n913_45002# a_1847_42826# 0.294312f
C4912 a_1115_44172# a_1467_44172# 0.115277f
C4913 a_8270_45546# VDD 1.26092f
C4914 a_175_44278# a_453_43940# 0.112594f
C4915 a_16327_47482# a_20835_44721# 0.157393f
C4916 a_n755_45592# a_n443_42852# 0.469263f
C4917 a_3160_47472# a_n1151_42308# 0.357683f
C4918 a_2905_45572# a_3381_47502# 0.208262f
C4919 a_5891_43370# a_7765_42852# 0.168516f
C4920 a_n1613_43370# a_n1917_43396# 0.153085f
C4921 a_n755_45592# a_375_42282# 0.366231f
C4922 a_12861_44030# a_6755_46942# 0.376009f
C4923 a_2747_46873# a_2864_46660# 0.174836f
C4924 a_22581_37893# a_22889_38993# 0.112329f
C4925 a_11599_46634# a_10467_46802# 0.261176f
C4926 a_2982_43646# a_4361_42308# 0.545077f
C4927 a_3357_43084# CLK 2.63944f
C4928 a_n2017_45002# VDD 3.8321f
C4929 a_n2438_43548# a_1138_42852# 0.646257f
C4930 a_12549_44172# a_10903_43370# 0.792848f
C4931 a_12861_44030# a_8049_45260# 0.109405f
C4932 a_12379_42858# a_12089_42308# 0.16885f
C4933 a_3422_30871# VDAC_N 0.480156f
C4934 a_3483_46348# a_5937_45572# 0.767636f
C4935 a_n1151_42308# a_413_45260# 0.135643f
C4936 a_5111_44636# a_9803_43646# 0.118936f
C4937 a_n2017_45002# a_16137_43396# 0.63011f
C4938 a_1123_46634# VDD 0.469393f
C4939 a_20640_44752# a_19279_43940# 0.22152f
C4940 a_19615_44636# a_18579_44172# 0.158449f
C4941 a_9290_44172# a_11823_42460# 0.864145f
C4942 a_n1613_43370# a_n1917_44484# 0.153277f
C4943 a_18727_42674# a_18907_42674# 0.185422f
C4944 a_19164_43230# VDD 0.278643f
C4945 a_13759_46122# VDD 0.399995f
C4946 a_4185_45028# a_22959_45036# 0.17601f
C4947 a_526_44458# a_1423_45028# 0.133656f
C4948 a_584_46384# a_458_43396# 0.196763f
C4949 a_n4209_39304# C7_P_btm 0.184297f
C4950 a_14021_43940# a_22959_43396# 0.191956f
C4951 a_n2956_37592# a_n3565_37414# 0.304738f
C4952 a_6197_43396# a_7112_43396# 0.118423f
C4953 a_10227_46804# a_10835_43094# 0.295543f
C4954 a_n1613_43370# a_n1853_43023# 0.423772f
C4955 a_413_45260# a_327_44734# 0.195096f
C4956 a_13661_43548# a_17339_46660# 0.599051f
C4957 a_5807_45002# a_765_45546# 0.103324f
C4958 a_15743_43084# a_15567_42826# 0.215954f
C4959 a_n2840_44458# VDD 0.247948f
C4960 a_5649_42852# a_5111_42852# 0.110096f
C4961 a_1823_45246# a_4361_42308# 0.11884f
C4962 a_18079_43940# VDD 0.162408f
C4963 a_22731_47423# VDD 0.196667f
C4964 a_21811_47423# SINGLE_ENDED 0.215228f
C4965 a_13661_43548# a_1307_43914# 0.396211f
C4966 a_12861_44030# a_20193_45348# 0.680394f
C4967 a_n2661_46634# a_13017_45260# 0.123713f
C4968 a_14209_32519# VDD 0.284433f
C4969 a_13661_43548# a_18579_44172# 0.229269f
C4970 a_15673_47210# a_16023_47582# 0.228897f
C4971 a_14955_47212# a_10227_46804# 0.175517f
C4972 a_n3420_38528# a_n3420_37984# 0.113087f
C4973 a_15507_47210# a_16588_47582# 0.102325f
C4974 a_16241_47178# a_16327_47482# 0.185907f
C4975 a_4099_45572# VDD 0.296272f
C4976 a_n2956_37592# a_n4209_39304# 0.102982f
C4977 a_12861_44030# a_18285_46348# 0.247326f
C4978 a_2609_46660# a_3177_46902# 0.17072f
C4979 a_2443_46660# a_2959_46660# 0.110816f
C4980 a_19250_35138# VDD 0.323729f
C4981 a_3090_45724# a_11415_45002# 0.16525f
C4982 a_6151_47436# a_5907_45546# 0.274247f
C4983 a_12089_42308# a_12800_43218# 0.15794f
C4984 a_17730_32519# VDD 0.289738f
C4985 a_n746_45260# VDD 1.41433f
C4986 a_7499_43078# a_10695_43548# 0.124597f
C4987 a_18184_42460# a_19279_43940# 0.132218f
C4988 a_18985_46122# a_19553_46090# 0.16939f
C4989 a_18819_46122# a_19335_46494# 0.108964f
C4990 a_n699_43396# a_104_43370# 0.21575f
C4991 a_12465_44636# a_14673_44172# 0.101564f
C4992 a_16327_47482# a_20679_44626# 0.318301f
C4993 a_10227_46804# a_11967_42832# 0.461417f
C4994 a_10586_45546# a_11962_45724# 0.137051f
C4995 a_n357_42282# a_n443_42852# 0.763015f
C4996 a_n4064_39616# a_n2302_39866# 0.239588f
C4997 a_n2661_42282# a_6293_42852# 0.16527f
C4998 a_14539_43914# a_17595_43084# 0.141972f
C4999 a_2711_45572# a_6171_45002# 0.457554f
C5000 a_n1613_43370# a_n1699_43638# 0.160308f
C5001 a_n357_42282# a_375_42282# 0.142311f
C5002 a_17339_46660# a_11967_42832# 0.493072f
C5003 a_7754_39964# RST_Z 0.843939f
C5004 a_22581_37893# a_22613_38993# 0.275268f
C5005 a_22527_39145# a_22537_39537# 0.351623f
C5006 VDAC_Pi VDD 0.591846f
C5007 a_n2109_45247# VDD 0.266396f
C5008 a_14180_45002# a_14537_43396# 0.143922f
C5009 a_12891_46348# a_10903_43370# 0.132903f
C5010 a_n13_43084# a_133_42852# 0.171361f
C5011 a_n2312_39304# a_n4209_39304# 0.19527f
C5012 a_5164_46348# a_5497_46414# 0.203417f
C5013 a_3483_46348# a_8199_44636# 1.81719f
C5014 a_3090_45724# a_13259_45724# 0.261789f
C5015 a_2107_46812# a_9049_44484# 0.240008f
C5016 a_3160_47472# a_413_45260# 0.208121f
C5017 a_n1435_47204# a_3357_43084# 1.08491f
C5018 a_17538_32519# VDD 0.352239f
C5019 a_22612_30879# VCM 0.473529f
C5020 a_383_46660# VDD 0.198466f
C5021 a_20679_44626# a_20835_44721# 0.105995f
C5022 a_20640_44752# a_20766_44850# 0.17072f
C5023 a_13249_42308# a_5534_30871# 0.215947f
C5024 a_11967_42832# a_18579_44172# 0.158329f
C5025 a_10903_43370# a_11322_45546# 0.313957f
C5026 a_12465_44636# a_12607_44458# 0.186652f
C5027 a_n1613_43370# a_n1699_44726# 0.166123f
C5028 a_19339_43156# VDD 0.338297f
C5029 a_n2293_43922# a_12281_43396# 0.147288f
C5030 a_13351_46090# VDD 0.238036f
C5031 a_1414_42308# a_n97_42460# 0.196768f
C5032 a_22485_38105# VDD 1.31335f
C5033 a_10227_46804# a_5807_45002# 0.262866f
C5034 a_n2810_45028# a_n3565_37414# 0.135518f
C5035 a_18494_42460# a_18907_42674# 0.11494f
C5036 a_6765_43638# a_6547_43396# 0.209641f
C5037 a_10227_46804# a_10518_42984# 0.225803f
C5038 a_n1613_43370# a_n2157_42858# 0.303592f
C5039 a_4791_45118# a_2324_44458# 0.19212f
C5040 a_19721_31679# VDD 0.521155f
C5041 a_3232_43370# a_9313_44734# 0.11426f
C5042 a_20820_30879# a_12741_44636# 0.103478f
C5043 a_n881_46662# a_6511_45714# 0.149116f
C5044 a_17973_43940# VDD 0.265874f
C5045 a_22223_47212# VDD 0.236555f
C5046 a_4883_46098# SINGLE_ENDED 0.1664f
C5047 a_12861_44030# a_11691_44458# 0.196929f
C5048 a_3090_45724# a_17478_45572# 0.128299f
C5049 a_22591_43396# VDD 0.280354f
C5050 a_11323_42473# a_5742_30871# 0.198522f
C5051 a_16922_45042# a_743_42282# 0.120316f
C5052 a_20731_47026# VDD 0.132317f
C5053 a_n1613_43370# a_n1761_44111# 0.148121f
C5054 a_167_45260# a_1423_45028# 0.123079f
C5055 a_15673_47210# a_16327_47482# 0.206019f
C5056 a_n237_47217# a_8128_46384# 0.113499f
C5057 a_3175_45822# VDD 0.193907f
C5058 a_18194_35068# VDD 2.24958f
C5059 C0_P_btm C0_dummy_P_btm 7.97415f
C5060 a_n2293_46634# a_526_44458# 0.579444f
C5061 a_22591_44484# VDD 0.223346f
C5062 a_n971_45724# VDD 4.911799f
C5063 SMPL_ON_P CLK_DATA 0.200962f
C5064 a_8975_43940# a_9313_44734# 0.391938f
C5065 a_765_45546# a_n357_42282# 0.209746f
C5066 a_2324_44458# a_6945_45028# 0.183081f
C5067 a_n699_43396# a_n97_42460# 0.152094f
C5068 a_n1059_45260# a_791_42968# 0.122941f
C5069 a_310_45028# a_n443_42852# 0.376934f
C5070 a_2905_45572# a_3160_47472# 0.54473f
C5071 a_n237_47217# a_6151_47436# 0.360224f
C5072 a_5891_43370# a_7227_42852# 0.129383f
C5073 a_n863_45724# a_1423_45028# 0.113534f
C5074 a_7499_43078# a_n913_45002# 0.548687f
C5075 a_7754_39964# VDD 0.848281f
C5076 a_6151_47436# a_8270_45546# 0.142873f
C5077 CAL_N a_22629_38406# 0.204616f
C5078 a_n2293_45010# VDD 1.885f
C5079 SMPL_ON_P a_n1794_35242# 6.11493f
C5080 a_n2497_47436# a_n863_45724# 0.337007f
C5081 a_9313_44734# VDD 0.389068f
C5082 a_5164_46348# a_5204_45822# 0.132894f
C5083 a_584_46384# a_2382_45260# 0.185451f
C5084 a_2905_45572# a_413_45260# 0.124898f
C5085 a_16327_47482# a_21188_45572# 0.227468f
C5086 a_20974_43370# VDD 0.550101f
C5087 a_22612_30879# VREF_GND 0.168163f
C5088 a_21588_30879# VCM 0.179761f
C5089 a_601_46902# VDD 0.204253f
C5090 a_20640_44752# a_20835_44721# 0.20669f
C5091 a_13661_43548# a_11827_44484# 0.120515f
C5092 a_18599_43230# VDD 0.197104f
C5093 a_11341_43940# a_15493_43940# 0.216602f
C5094 a_12594_46348# VDD 1.03351f
C5095 a_1467_44172# a_n97_42460# 0.190191f
C5096 a_3422_30871# a_2982_43646# 0.140944f
C5097 a_12549_44172# a_12429_44172# 0.137881f
C5098 a_526_44458# a_626_44172# 0.180416f
C5099 a_3090_45724# a_n2661_42834# 0.164804f
C5100 a_13507_46334# a_12549_44172# 0.363125f
C5101 a_7754_38968# a_3754_38470# 0.209356f
C5102 a_n971_45724# a_4646_46812# 0.303249f
C5103 a_16327_47482# a_19321_45002# 0.925259f
C5104 a_6031_43396# a_7112_43396# 0.101963f
C5105 a_6197_43396# a_6547_43396# 0.216095f
C5106 a_n2956_37592# a_n4209_37414# 0.145558f
C5107 a_10227_46804# a_10083_42826# 0.292997f
C5108 a_7577_46660# a_8492_46660# 0.118423f
C5109 a_18114_32519# VDD 0.550506f
C5110 a_16922_45042# a_20193_45348# 0.328274f
C5111 a_3090_45724# a_17715_44484# 0.108364f
C5112 a_n881_46662# a_6472_45840# 0.179318f
C5113 a_17737_43940# VDD 0.285511f
C5114 a_n2293_42282# a_n2472_42282# 0.163758f
C5115 a_12465_44636# VDD 0.773277f
C5116 a_16327_47482# a_18184_42460# 0.168018f
C5117 a_13661_43548# a_15595_45028# 0.214904f
C5118 a_3090_45724# a_15861_45028# 0.125763f
C5119 a_13887_32519# VDD 0.424101f
C5120 a_10723_42308# a_5742_30871# 0.185564f
C5121 a_n1613_43370# a_n2065_43946# 0.30437f
C5122 a_2711_45572# a_10193_42453# 0.218272f
C5123 a_15673_47210# a_16241_47178# 0.183195f
C5124 a_15507_47210# a_16023_47582# 0.109156f
C5125 a_8515_42308# VDD 0.194691f
C5126 a_12861_44030# a_18143_47464# 0.394543f
C5127 a_n4064_40160# a_n3565_37414# 4.2965f
C5128 a_2711_45572# VDD 1.22011f
C5129 a_2443_46660# a_2609_46660# 0.579196f
C5130 a_11453_44696# a_15227_44166# 0.979188f
C5131 a_12861_44030# a_765_45546# 0.190301f
C5132 EN_VIN_BSTR_N VDD 1.20174f
C5133 C1_P_btm C0_dummy_P_btm 1.24905f
C5134 a_10227_46804# a_n357_42282# 0.103631f
C5135 a_16388_46812# a_16721_46634# 0.222024f
C5136 a_22485_44484# VDD 0.258874f
C5137 a_10057_43914# a_9313_44734# 0.139382f
C5138 a_n881_46662# a_n745_45366# 0.152998f
C5139 a_5204_45822# a_5066_45546# 0.402457f
C5140 a_18819_46122# a_18985_46122# 0.749955f
C5141 a_n1059_45260# a_685_42968# 0.103646f
C5142 a_16327_47482# a_20362_44736# 0.213851f
C5143 a_584_46384# a_453_43940# 0.125447f
C5144 a_13059_46348# a_14537_43396# 0.30244f
C5145 a_10586_45546# a_11525_45546# 0.115475f
C5146 a_16877_42852# VDD 0.192454f
C5147 a_n971_45724# a_6545_47178# 0.295443f
C5148 a_2952_47436# a_3160_47472# 0.192116f
C5149 a_5891_43370# a_5755_42852# 0.160849f
C5150 a_14021_43940# a_20974_43370# 0.893848f
C5151 a_12741_44636# a_n2293_43922# 0.114756f
C5152 a_7499_43078# a_n1059_45260# 0.277353f
C5153 a_2324_44458# a_6298_44484# 0.315008f
C5154 a_n1613_43370# a_n2129_43609# 0.44294f
C5155 CAL_N CAL_P 5.92093f
C5156 a_22589_40055# a_22889_38993# 0.19183f
C5157 a_22527_39145# a_22613_38993# 0.12129f
C5158 a_2437_43646# CLK 0.101524f
C5159 a_2982_43646# a_21487_43396# 0.169809f
C5160 a_3626_43646# a_743_42282# 0.147999f
C5161 a_n2472_45002# VDD 0.217954f
C5162 a_13556_45296# a_14537_43396# 0.590856f
C5163 a_768_44030# a_9290_44172# 0.189655f
C5164 a_n97_42460# a_5742_30871# 0.259664f
C5165 a_n881_46662# a_15765_45572# 0.58719f
C5166 a_n1151_42308# a_n467_45028# 0.406349f
C5167 a_5068_46348# a_5204_45822# 0.20685f
C5168 a_16327_47482# a_21363_45546# 0.276554f
C5169 a_14401_32519# VDD 0.562673f
C5170 a_n3674_39304# a_n3420_39616# 0.152699f
C5171 a_22612_30879# VREF 1.73216f
C5172 a_5891_43370# a_7845_44172# 0.119969f
C5173 a_33_46660# VDD 0.272723f
C5174 a_20640_44752# a_20679_44626# 0.582607f
C5175 a_n2293_42834# a_n97_42460# 0.17628f
C5176 a_19321_45002# a_20567_45036# 0.205038f
C5177 a_18817_42826# VDD 0.204624f
C5178 a_11341_43940# a_22223_43948# 0.175191f
C5179 a_8199_44636# CLK 0.231904f
C5180 a_12005_46116# VDD 0.518463f
C5181 a_3754_38802# VDAC_Ni 0.301032f
C5182 a_n971_45724# a_3877_44458# 0.927248f
C5183 a_6197_43396# a_6765_43638# 0.17072f
C5184 a_14033_45822# VDD 0.195067f
C5185 a_4185_45028# a_n2661_42282# 0.833759f
C5186 a_8145_46902# a_7927_46660# 0.209641f
C5187 a_n2661_43370# a_n2661_44458# 1.0558f
C5188 a_16922_45042# a_11691_44458# 0.428229f
C5189 a_19778_44110# a_21005_45260# 0.135527f
C5190 a_22591_46660# a_20820_30879# 0.166885f
C5191 a_11415_45002# a_12741_44636# 1.07921f
C5192 a_n2293_46634# a_n863_45724# 0.157683f
C5193 a_15682_43940# VDD 1.22657f
C5194 a_21811_47423# VDD 0.201359f
C5195 a_13507_46334# SINGLE_ENDED 0.111959f
C5196 a_167_45260# a_2277_45546# 0.214157f
C5197 a_n1151_42308# a_n452_44636# 0.238824f
C5198 a_13661_43548# a_15415_45028# 0.133591f
C5199 a_22223_43396# VDD 0.279195f
C5200 a_22000_46634# VDD 0.257047f
C5201 a_16922_45042# a_4190_30871# 0.353708f
C5202 a_8199_44636# a_10951_45334# 0.237774f
C5203 a_10903_43370# a_3232_43370# 0.114259f
C5204 a_5934_30871# VDD 0.431427f
C5205 a_15507_47210# a_16327_47482# 0.425757f
C5206 a_n1741_47186# a_12891_46348# 0.107238f
C5207 a_12861_44030# a_10227_46804# 0.291378f
C5208 a_12861_44030# a_17339_46660# 1.25428f
C5209 a_11530_34132# VDD 0.362849f
C5210 C1_P_btm C0_P_btm 11.2332f
C5211 C2_P_btm C0_dummy_P_btm 7.14548f
C5212 a_15743_43084# a_4190_30871# 0.290729f
C5213 a_16751_45260# a_17023_45118# 0.13675f
C5214 a_5257_43370# a_6419_46155# 0.186651f
C5215 a_17730_32519# C9_N_btm 0.215899f
C5216 a_20512_43084# VDD 0.317257f
C5217 a_n4318_39304# a_n4209_39304# 0.135369f
C5218 a_n815_47178# VDD 0.380339f
C5219 a_n699_43396# a_n2661_42834# 0.131393f
C5220 a_12741_44636# a_13259_45724# 0.113445f
C5221 a_n784_42308# a_5934_30871# 0.142087f
C5222 a_10586_45546# a_11322_45546# 0.220166f
C5223 a_16327_47482# a_20159_44458# 0.270426f
C5224 a_12861_44030# a_18579_44172# 0.221909f
C5225 a_584_46384# a_1414_42308# 0.321387f
C5226 a_n3420_39616# a_n4064_39616# 6.66063f
C5227 a_16245_42852# VDD 0.205729f
C5228 a_2952_47436# a_2905_45572# 0.318161f
C5229 a_n971_45724# a_6151_47436# 0.29974f
C5230 a_2063_45854# a_n1151_42308# 0.425035f
C5231 a_n1794_35242# a_n1696_35090# 0.462414f
C5232 a_18579_44172# a_19700_43370# 0.175511f
C5233 a_n2661_42834# a_n4318_38680# 0.102282f
C5234 a_n1613_43370# a_n2433_43396# 0.299968f
C5235 a_2324_44458# a_5518_44484# 0.112753f
C5236 a_22537_40625# a_22537_39537# 0.604835f
C5237 a_n881_46662# a_2107_46812# 0.138703f
C5238 a_11206_38545# CAL_P 0.234643f
C5239 a_7754_40130# VDD 13.6809f
C5240 a_19321_45002# a_19594_46812# 0.267862f
C5241 a_n97_42460# a_n13_43084# 0.13246f
C5242 a_n356_44636# a_17303_42282# 0.10316f
C5243 a_n2661_45010# VDD 0.842431f
C5244 a_n2497_47436# a_n2293_45546# 0.307373f
C5245 a_12991_46634# a_12816_46660# 0.233657f
C5246 a_11453_44696# a_10809_44734# 0.274367f
C5247 a_3080_42308# a_5934_30871# 1.27306f
C5248 a_n755_45592# a_8147_43396# 0.134231f
C5249 a_n971_45724# a_5111_44636# 0.381443f
C5250 a_n1435_47204# a_2437_43646# 0.191468f
C5251 a_5068_46348# a_5164_46348# 0.31819f
C5252 a_16327_47482# a_20623_45572# 0.168593f
C5253 a_21381_43940# VDD 0.344882f
C5254 a_21588_30879# VREF 0.860047f
C5255 a_171_46873# VDD 0.539781f
C5256 a_20362_44736# a_20679_44626# 0.102355f
C5257 a_n2661_43370# a_n2840_43370# 0.172532f
C5258 a_22612_30879# VIN_N 0.19035f
C5259 a_10903_43370# a_10193_42453# 0.402091f
C5260 a_n1613_43370# a_n2433_44484# 0.29864f
C5261 a_13259_45724# a_16375_45002# 0.60955f
C5262 a_526_44458# a_n443_42852# 2.06448f
C5263 a_18249_42858# VDD 0.250132f
C5264 a_10903_43370# VDD 2.60588f
C5265 a_16763_47508# a_5807_45002# 0.127783f
C5266 a_16327_47482# a_13747_46662# 0.128159f
C5267 a_6031_43396# a_6547_43396# 0.105995f
C5268 a_18184_42460# a_18057_42282# 0.19301f
C5269 a_n913_45002# a_3537_45260# 0.148413f
C5270 a_n143_45144# a_n37_45144# 0.13675f
C5271 a_7411_46660# a_8492_46660# 0.102325f
C5272 a_7577_46660# a_7927_46660# 0.206455f
C5273 a_18114_32519# C10_N_btm 0.460005f
C5274 a_7229_43940# a_7640_43914# 0.177622f
C5275 a_18184_42460# a_18494_42460# 1.31047f
C5276 a_20202_43084# a_12741_44636# 0.22243f
C5277 a_14955_43940# VDD 0.253201f
C5278 a_4883_46098# VDD 1.12729f
C5279 a_4185_45028# a_5379_42460# 0.189676f
C5280 a_11823_42460# a_743_42282# 0.147603f
C5281 a_18287_44626# a_18579_44172# 0.107662f
C5282 a_10227_46804# CLK 0.207445f
C5283 a_167_45260# a_1609_45822# 0.141505f
C5284 a_13661_43548# a_14797_45144# 0.116989f
C5285 a_584_46384# a_n699_43396# 0.632931f
C5286 a_18189_46348# a_16375_45002# 0.165328f
C5287 a_5649_42852# VDD 0.438443f
C5288 a_21188_46660# VDD 0.284105f
C5289 a_16922_45042# a_21259_43561# 0.108631f
C5290 a_15811_47375# a_15673_47210# 0.281607f
C5291 a_11599_46634# a_16327_47482# 0.526398f
C5292 a_7963_42308# VDD 0.266057f
C5293 a_11341_43940# a_10341_43396# 0.289072f
C5294 w_11334_34010# a_n1794_35242# 3.10971f
C5295 a_n2497_47436# a_1138_42852# 0.144386f
C5296 EN_VIN_BSTR_N C10_N_btm 0.320569f
C5297 a_n217_35174# VDD 0.296751f
C5298 C2_P_btm C0_P_btm 0.827449f
C5299 a_2982_43646# a_5342_30871# 0.178973f
C5300 a_16751_45260# a_16922_45042# 0.12103f
C5301 SMPL_ON_N COMP_P 2.13481f
C5302 a_5257_43370# a_6165_46155# 0.11382f
C5303 a_10341_42308# a_11554_42852# 0.170124f
C5304 a_3626_43646# a_19647_42308# 0.170024f
C5305 a_n1605_47204# VDD 0.20224f
C5306 a_n881_46662# a_n1059_45260# 0.121542f
C5307 a_n1613_43370# a_n913_45002# 0.686014f
C5308 a_765_45546# a_380_45546# 0.141908f
C5309 a_8685_43396# VDD 0.261626f
C5310 a_3218_45724# a_3316_45546# 0.162813f
C5311 a_n863_45724# a_1609_45822# 0.117311f
C5312 a_10586_45546# a_10490_45724# 0.235237f
C5313 a_n3420_39616# a_n2946_39866# 0.236674f
C5314 a_18597_46090# a_2982_43646# 0.239147f
C5315 a_19692_46634# a_20512_43084# 0.387138f
C5316 a_2324_44458# a_5343_44458# 0.255488f
C5317 a_22589_40055# a_22581_37893# 0.461959f
C5318 a_22589_40599# a_22537_39537# 0.380009f
C5319 a_2747_46873# a_2609_46660# 0.347674f
C5320 a_n356_44636# a_4958_30871# 0.46356f
C5321 a_n2840_45002# VDD 0.289706f
C5322 a_13556_45296# a_13777_45326# 0.101558f
C5323 a_n2293_46634# a_1823_45246# 0.230429f
C5324 a_n2293_42834# a_n2661_42834# 0.202366f
C5325 a_742_44458# a_949_44458# 0.185221f
C5326 a_4791_45118# a_n913_45002# 0.254334f
C5327 a_n881_46662# a_15599_45572# 0.601034f
C5328 a_16327_47482# a_20841_45814# 0.161808f
C5329 a_19741_43940# VDD 0.153579f
C5330 a_n133_46660# VDD 0.483405f
C5331 a_20362_44736# a_20640_44752# 0.118759f
C5332 a_21588_30879# VIN_N 0.106594f
C5333 a_3483_46348# a_10907_45822# 0.140023f
C5334 a_17333_42852# VDD 0.525529f
C5335 a_7754_38968# a_7754_38636# 0.296258f
C5336 a_n4064_39072# EN_VIN_BSTR_P 1.00234f
C5337 a_16327_47482# a_13661_43548# 0.132061f
C5338 a_6293_42852# a_6197_43396# 0.213423f
C5339 a_n97_42460# a_10341_43396# 0.917198f
C5340 a_n1059_45260# a_3537_45260# 0.162323f
C5341 a_7577_46660# a_8145_46902# 0.170059f
C5342 a_n901_43156# a_n1076_43230# 0.234322f
C5343 a_n1853_43023# a_n1736_43218# 0.183149f
C5344 a_3090_45724# a_2324_44458# 0.684819f
C5345 a_11415_45002# a_22591_46660# 0.172844f
C5346 a_n881_46662# a_5263_45724# 0.180025f
C5347 a_13483_43940# VDD 0.219591f
C5348 a_21496_47436# VDD 0.198362f
C5349 a_n743_46660# a_6171_45002# 0.140224f
C5350 a_167_45260# a_n443_42852# 0.246952f
C5351 a_12861_44030# a_11827_44484# 0.466435f
C5352 a_13661_43548# a_14537_43396# 0.505634f
C5353 a_13678_32519# VDD 0.454512f
C5354 a_10533_42308# a_10723_42308# 0.23663f
C5355 a_n2293_43922# a_n97_42460# 0.136247f
C5356 a_21363_46634# VDD 0.357368f
C5357 a_12549_44172# a_3422_30871# 0.148646f
C5358 a_5937_45572# a_8191_45002# 0.180306f
C5359 a_8270_45546# a_5883_43914# 0.20967f
C5360 a_8199_44636# a_8953_45002# 0.12099f
C5361 a_6123_31319# VDD 0.533328f
C5362 a_n237_47217# a_n881_46662# 0.958566f
C5363 a_15507_47210# a_15673_47210# 0.81159f
C5364 a_21363_45546# a_21188_45572# 0.233657f
C5365 EN_VIN_BSTR_N C9_N_btm 0.226529f
C5366 EN_VIN_BSTR_P VDD 0.922997f
C5367 C2_P_btm C1_P_btm 5.24136f
C5368 C3_P_btm C0_P_btm 0.409238f
C5369 C4_P_btm C0_dummy_P_btm 0.113156f
C5370 a_17339_46660# a_15743_43084# 0.450316f
C5371 a_n971_45724# a_7499_43078# 0.857375f
C5372 a_3626_43646# a_19511_42282# 0.182478f
C5373 SMPL_ON_P VDD 0.613663f
C5374 a_8270_45546# a_8162_45546# 0.170838f
C5375 a_n1613_43370# a_n1059_45260# 0.202724f
C5376 a_n784_42308# a_6123_31319# 0.144274f
C5377 a_8035_47026# VDD 0.132317f
C5378 a_13059_46348# a_13556_45296# 0.274813f
C5379 a_16327_47482# a_11967_42832# 0.241578f
C5380 a_n863_45724# a_n443_42852# 0.556081f
C5381 a_584_46384# a_1115_44172# 0.174981f
C5382 a_15597_42852# VDD 0.239357f
C5383 a_n3565_39590# a_n4064_39616# 0.231239f
C5384 a_n237_47217# a_n443_46116# 0.110841f
C5385 a_n2293_45546# a_626_44172# 0.150062f
C5386 a_4185_45028# a_n356_44636# 1.54308f
C5387 a_n863_45724# a_375_42282# 0.451905f
C5388 a_2747_46873# a_2443_46660# 0.129886f
C5389 a_n1613_43370# a_948_46660# 0.281392f
C5390 a_3422_30871# a_n1794_35242# 0.828871f
C5391 a_9482_43914# a_13777_45326# 0.206086f
C5392 a_10796_42968# a_10341_42308# 0.65943f
C5393 a_10991_42826# a_10922_42852# 0.209641f
C5394 a_3626_43646# a_4921_42308# 0.431551f
C5395 a_3080_42308# a_6123_31319# 1.45722f
C5396 a_11691_44458# a_16979_44734# 0.12231f
C5397 a_584_46384# a_413_45260# 0.164383f
C5398 a_n1151_42308# a_n967_45348# 0.170453f
C5399 a_11823_42460# a_5534_30871# 0.511874f
C5400 a_n2438_43548# VDD 3.40589f
C5401 a_7640_43914# a_7542_44172# 0.20977f
C5402 a_19321_45002# a_19778_44110# 0.568668f
C5403 a_16327_47482# a_18989_43940# 0.100946f
C5404 a_12741_44636# a_8696_44636# 2.20704f
C5405 a_18083_42858# VDD 0.408512f
C5406 a_11133_46155# VDD 0.176249f
C5407 a_13483_43940# a_14021_43940# 0.109097f
C5408 a_526_44458# a_1307_43914# 0.467539f
C5409 a_22775_42308# VDD 0.426061f
C5410 a_16327_47482# a_5807_45002# 0.451783f
C5411 a_6031_43396# a_6197_43396# 0.581047f
C5412 a_n913_45002# a_3065_45002# 0.225034f
C5413 a_7411_46660# a_7927_46660# 0.105839f
C5414 a_9313_45822# a_5937_45572# 0.137696f
C5415 a_13259_45724# a_n97_42460# 0.182889f
C5416 a_19778_44110# a_18184_42460# 0.119002f
C5417 a_765_45546# a_167_45260# 0.276049f
C5418 a_12429_44172# VDD 0.169047f
C5419 a_13507_46334# VDD 1.4135f
C5420 a_1823_45246# a_1609_45822# 0.35471f
C5421 a_21855_43396# VDD 0.289066f
C5422 a_20623_46660# VDD 0.194217f
C5423 a_n443_42852# a_11823_42460# 0.356965f
C5424 a_8199_44636# a_8191_45002# 0.234072f
C5425 a_7227_42308# VDD 0.296912f
C5426 a_n3565_38502# a_n4209_38216# 5.84657f
C5427 a_n746_45260# a_n881_46662# 0.190303f
C5428 a_15507_47210# a_15811_47375# 0.170975f
C5429 a_11967_42832# a_12379_42858# 0.492977f
C5430 a_11599_46634# a_16388_46812# 0.24092f
C5431 a_n1057_35174# VDD 0.338357f
C5432 C5_P_btm C0_dummy_P_btm 0.11375f
C5433 C3_P_btm C1_P_btm 8.06688f
C5434 C4_P_btm C0_P_btm 0.138331f
C5435 a_n1741_47186# VDD 0.912651f
C5436 a_11415_45002# a_13259_45724# 0.505354f
C5437 a_15227_44166# a_2711_45572# 0.113396f
C5438 a_2713_42308# a_2903_42308# 0.23738f
C5439 a_5111_44636# a_5649_42852# 0.121004f
C5440 a_13059_46348# a_9482_43914# 0.448068f
C5441 a_n2293_45546# a_1609_45822# 0.159696f
C5442 a_12861_44030# a_19279_43940# 0.152657f
C5443 a_10586_45546# a_10193_42453# 0.380236f
C5444 a_n3690_39616# a_n3420_39616# 0.431154f
C5445 a_n3565_39590# a_n2946_39866# 0.406088f
C5446 a_n4209_39590# a_n2302_39866# 0.406459f
C5447 a_n4334_39616# a_n4064_39616# 0.4504f
C5448 a_n237_47217# a_4791_45118# 0.10712f
C5449 a_10586_45546# VDD 0.582083f
C5450 a_22589_40055# a_22527_39145# 0.130029f
C5451 a_22537_40625# a_22581_37893# 0.656829f
C5452 a_n1613_43370# a_1123_46634# 0.358475f
C5453 a_768_44030# a_n2293_46634# 0.26984f
C5454 a_2982_43646# a_4190_30871# 0.3223f
C5455 a_9482_43914# a_13556_45296# 0.726155f
C5456 a_5205_44484# a_1423_45028# 0.821456f
C5457 a_11901_46660# a_12816_46660# 0.125324f
C5458 a_10796_42968# a_10922_42852# 0.170059f
C5459 a_10835_43094# a_10341_42308# 0.541777f
C5460 a_11691_44458# a_14539_43914# 0.268287f
C5461 a_n2661_46634# a_11823_42460# 0.331717f
C5462 a_n743_46660# a_10193_42453# 0.25279f
C5463 a_16327_47482# a_20107_45572# 0.674639f
C5464 a_11967_42832# a_20679_44626# 0.863531f
C5465 a_n743_46660# VDD 1.75634f
C5466 a_20159_44458# a_20362_44736# 0.233657f
C5467 a_22612_30879# EN_OFFSET_CAL 0.118817f
C5468 a_11189_46129# a_10193_42453# 0.123385f
C5469 a_13747_46662# a_18184_42460# 0.123281f
C5470 a_16327_47482# a_18374_44850# 0.16003f
C5471 a_17701_42308# VDD 0.243354f
C5472 a_4958_30871# a_17531_42308# 0.192941f
C5473 a_11189_46129# VDD 0.944289f
C5474 a_20935_43940# a_21115_43940# 0.185422f
C5475 a_21613_42308# VDD 0.27399f
C5476 a_n3420_39072# EN_VIN_BSTR_P 0.814814f
C5477 a_6031_43396# a_6293_42852# 0.163953f
C5478 a_12549_44172# a_20556_43646# 0.125209f
C5479 a_n755_45592# a_n356_44636# 2.42652f
C5480 a_13747_46662# a_13059_46348# 0.273684f
C5481 a_5807_45002# a_16721_46634# 0.112018f
C5482 a_7715_46873# a_7577_46660# 0.205227f
C5483 a_3232_43370# a_5891_43370# 0.137859f
C5484 a_11750_44172# VDD 0.131662f
C5485 a_10193_42453# a_4361_42308# 0.274131f
C5486 a_21177_47436# VDD 0.179587f
C5487 a_768_44030# a_626_44172# 0.186913f
C5488 a_1823_45246# a_n443_42852# 0.125287f
C5489 a_4361_42308# VDD 0.42717f
C5490 a_20841_46902# VDD 0.20446f
C5491 a_5937_45572# a_6709_45028# 0.629301f
C5492 a_6761_42308# VDD 0.259312f
C5493 a_5742_30871# C6_P_btm 0.170624f
C5494 a_n971_45724# a_n881_46662# 0.236696f
C5495 a_n746_45260# a_n1613_43370# 0.146842f
C5496 a_2553_47502# a_2747_46873# 0.14563f
C5497 a_11599_46634# a_15811_47375# 0.107881f
C5498 a_n2293_43922# a_n2293_42282# 0.19201f
C5499 a_2711_45572# a_n2661_43370# 0.112998f
C5500 a_3090_45724# a_15493_43396# 0.134629f
C5501 C3_P_btm C2_P_btm 5.99608f
C5502 C5_P_btm C0_P_btm 0.138093f
C5503 C4_P_btm C1_P_btm 0.128167f
C5504 a_13507_46334# a_19692_46634# 0.823157f
C5505 a_11599_46634# a_13059_46348# 0.371555f
C5506 EN_VIN_BSTR_N C7_N_btm 0.115875f
C5507 a_n1696_35090# VDD 2.24276f
C5508 C6_P_btm C0_dummy_P_btm 0.1194f
C5509 a_n2661_42282# a_1755_42282# 0.145244f
C5510 a_4915_47217# a_2711_45572# 0.265557f
C5511 a_16327_47482# a_n357_42282# 0.49929f
C5512 a_15227_44166# a_22000_46634# 0.154332f
C5513 a_5883_43914# a_9313_44734# 0.124999f
C5514 a_n2833_47464# CLK_DATA 0.331592f
C5515 a_n1920_47178# VDD 0.229556f
C5516 a_11823_42460# a_13291_42460# 0.257506f
C5517 a_n809_44244# a_n984_44318# 0.234322f
C5518 a_1823_45246# a_2437_43646# 0.324477f
C5519 a_n755_45592# a_3503_45724# 0.163919f
C5520 a_n1151_42308# a_n1761_44111# 0.642214f
C5521 a_n3565_39590# a_n3420_39616# 0.281955f
C5522 a_n971_45724# a_n443_46116# 0.129009f
C5523 a_n4209_39590# a_n4064_39616# 0.269818f
C5524 a_9290_44172# a_8975_43940# 0.114958f
C5525 a_n2293_45546# a_375_42282# 0.104283f
C5526 a_2324_44458# a_4223_44672# 0.56408f
C5527 a_22589_40599# a_22581_37893# 0.365664f
C5528 a_n1613_43370# a_383_46660# 0.182504f
C5529 a_9804_47204# a_n743_46660# 0.295465f
C5530 a_20447_31679# VDD 0.665793f
C5531 en_comp a_n2293_42834# 0.103485f
C5532 a_13348_45260# a_13556_45296# 0.189446f
C5533 a_n1925_42282# a_n2661_42282# 2.27741f
C5534 a_12469_46902# a_12251_46660# 0.209641f
C5535 a_10796_42968# a_10991_42826# 0.206455f
C5536 a_5891_43370# VDD 2.12137f
C5537 a_n971_45724# a_3537_45260# 0.266743f
C5538 a_18533_43940# VDD 0.182147f
C5539 a_11967_42832# a_20640_44752# 0.588649f
C5540 a_n1021_46688# VDD 0.226043f
C5541 a_9290_44172# a_10193_42453# 1.23123f
C5542 a_13747_46662# a_19778_44110# 0.670692f
C5543 a_16327_47482# a_18443_44721# 0.1665f
C5544 a_10903_43370# a_7499_43078# 0.888628f
C5545 a_17595_43084# VDD 0.168112f
C5546 a_4958_30871# a_17303_42282# 0.168656f
C5547 a_n2956_38216# a_n2946_37984# 0.150404f
C5548 a_9290_44172# VDD 2.74561f
C5549 a_19862_44208# a_15493_43940# 0.534481f
C5550 a_2324_44458# a_n2293_42834# 0.168086f
C5551 a_768_44030# a_9028_43914# 0.113848f
C5552 a_584_46384# a_n97_42460# 0.526796f
C5553 a_21887_42336# VDD 0.210392f
C5554 a_584_46384# a_n2661_46098# 0.17431f
C5555 a_12465_44636# a_n881_46662# 0.813228f
C5556 a_12549_44172# a_743_42282# 0.119701f
C5557 a_n357_42282# a_n356_44636# 0.308599f
C5558 a_7411_46660# a_7577_46660# 0.634781f
C5559 a_5807_45002# a_16388_46812# 0.235518f
C5560 a_13661_43548# a_13059_46348# 0.267127f
C5561 a_16547_43609# a_16414_43172# 0.143695f
C5562 a_n2472_42826# a_n4318_38680# 0.158196f
C5563 a_n1991_42858# a_n1076_43230# 0.123255f
C5564 a_n1853_43023# a_n13_43084# 0.109925f
C5565 w_11334_34010# VDD 1.9159f
C5566 a_10227_46804# a_11823_42460# 0.428745f
C5567 a_n881_46662# a_2711_45572# 0.170524f
C5568 a_n2293_46634# a_n2661_45546# 0.85166f
C5569 a_10807_43548# VDD 0.68049f
C5570 a_20990_47178# VDD 0.210484f
C5571 a_19787_47423# START 0.220891f
C5572 a_n2661_42834# a_n2661_43922# 0.841361f
C5573 a_15368_46634# a_15599_45572# 0.100853f
C5574 a_13661_43548# a_13556_45296# 0.559682f
C5575 a_1138_42852# a_n443_42852# 0.14758f
C5576 a_17715_44484# a_13259_45724# 0.391904f
C5577 VCM VSS 30.7148f
C5578 VREF_GND VSS 17.6497f
C5579 VREF VSS 8.8492f
C5580 VIN_N VSS 13.1487f
C5581 VIN_P VSS 13.1241f
C5582 CLK VSS 1.55797f
C5583 EN_OFFSET_CAL VSS 0.505642f
C5584 DATA[5] VSS 0.561058f
C5585 DATA[4] VSS 0.755679f
C5586 DATA[3] VSS 1.01838f
C5587 DATA[2] VSS 0.536983f
C5588 DATA[1] VSS 0.550109f
C5589 DATA[0] VSS 0.616231f
C5590 CLK_DATA VSS 0.488979f
C5591 SINGLE_ENDED VSS 0.60168f
C5592 START VSS 0.991673f
C5593 RST_Z VSS 11.362901f
C5594 VDD VSS 0.589075p
C5595 C10_N_btm VSS 0.210692p 
C5596 C9_N_btm VSS 79.926506f 
C5597 C8_N_btm VSS 45.547f 
C5598 C7_N_btm VSS 25.886099f 
C5599 C6_N_btm VSS 15.5273f 
C5600 C5_N_btm VSS 9.624539f 
C5601 C4_N_btm VSS 8.794849f 
C5602 C3_N_btm VSS 6.38289f 
C5603 C2_N_btm VSS 5.46028f 
C5604 C1_N_btm VSS 5.26099f 
C5605 C0_N_btm VSS 7.20283f 
C5606 C0_dummy_N_btm VSS 5.03035f 
C5607 C0_dummy_P_btm VSS 5.0181f 
C5608 C0_P_btm VSS 7.1984f 
C5609 C1_P_btm VSS 5.27428f 
C5610 C2_P_btm VSS 5.46972f 
C5611 C3_P_btm VSS 6.37616f 
C5612 C4_P_btm VSS 8.785789f 
C5613 C5_P_btm VSS 9.614769f 
C5614 C6_P_btm VSS 15.5172f 
C5615 C7_P_btm VSS 25.876501f 
C5616 C8_P_btm VSS 45.531998f 
C5617 C9_P_btm VSS 79.8995f 
C5618 C10_P_btm VSS 0.210676p 
C5619 a_21753_35634# VSS 0.728261f 
C5620 a_19998_35138# VSS 1.74918f 
C5621 a_19250_35138# VSS 1.6987f 
C5622 a_18194_35068# VSS 2.12114f 
C5623 EN_VIN_BSTR_N VSS 9.10061f 
C5624 a_11530_34132# VSS 14.0076f 
C5625 a_n217_35174# VSS 1.73474f 
C5626 EN_VIN_BSTR_P VSS 9.35043f 
C5627 a_n1057_35174# VSS 14.1073f 
C5628 a_n1696_35090# VSS 2.16403f 
C5629 a_n1550_35608# VSS 1.7497f 
C5630 a_n2002_35608# VSS 0.734464f 
C5631 a_22629_37990# VSS 0.468764f 
C5632 a_22629_38406# VSS 0.583873f 
C5633 CAL_P VSS 11.437099f 
C5634 a_22537_39537# VSS 2.60616f 
C5635 a_22889_38993# VSS 0.497542f 
C5636 a_22613_38993# VSS 0.357645f 
C5637 a_22581_37893# VSS 1.83807f 
C5638 a_22527_39145# VSS 2.28594f 
C5639 a_22589_40055# VSS 1.23689f 
C5640 a_22537_40625# VSS 1.5788f 
C5641 a_22589_40599# VSS 1.83268f 
C5642 CAL_N VSS 8.71062f 
C5643 a_11206_38545# VSS 0.713084f 
C5644 VDAC_P VSS 0.107582p 
C5645 a_8912_37509# VSS 3.72815f 
C5646 VDAC_N VSS 0.108181p 
C5647 a_6886_37412# VSS 3.84636f 
C5648 a_5700_37509# VSS 2.08109f 
C5649 a_5088_37509# VSS 2.72043f 
C5650 a_4338_37500# VSS 2.61032f 
C5651 a_3726_37500# VSS 4.48332f 
C5652 a_n2302_37690# VSS 0.513659f 
C5653 a_n4064_37440# VSS 1.7233f 
C5654 a_n2946_37690# VSS 0.517242f 
C5655 a_n3420_37440# VSS 5.23286f 
C5656 a_n3690_37440# VSS 0.548488f 
C5657 a_n3565_37414# VSS 3.1619f 
C5658 a_n4334_37440# VSS 0.561497f 
C5659 a_n4209_37414# VSS 3.16671f 
C5660 a_8530_39574# VSS 2.76228f 
C5661 a_7754_38470# VSS 3.24403f 
C5662 a_3754_38470# VSS 4.77654f 
C5663 VDAC_Ni VSS 2.86378f 
C5664 a_7754_38636# VSS 0.353706f 
C5665 a_3754_38802# VSS 0.390074f 
C5666 a_7754_38968# VSS 0.330037f 
C5667 a_3754_39134# VSS 0.401983f 
C5668 a_7754_39300# VSS 0.330682f 
C5669 a_3754_39466# VSS 0.401172f 
C5670 a_7754_39632# VSS 0.340942f 
C5671 VDAC_Pi VSS 3.50356f 
C5672 a_7754_39964# VSS 2.62481f 
C5673 a_7754_40130# VSS 2.84033f 
C5674 a_3754_39964# VSS 0.671366f 
C5675 a_2113_38308# VSS 2.64726f 
C5676 a_n2302_37984# VSS 0.483504f 
C5677 a_n4064_37984# VSS 1.65074f 
C5678 a_n2946_37984# VSS 0.485942f 
C5679 a_n3420_37984# VSS 1.75918f 
C5680 a_n3690_38304# VSS 0.517812f 
C5681 a_n3565_38216# VSS 1.49194f 
C5682 a_n4334_38304# VSS 0.529531f 
C5683 a_n4209_38216# VSS 3.03817f 
C5684 a_2684_37794# VSS 0.414596f 
C5685 a_1107_38525# VSS 0.6415f 
C5686 a_n2302_38778# VSS 0.483515f 
C5687 a_n4064_38528# VSS 1.69554f 
C5688 a_n2946_38778# VSS 0.485895f 
C5689 a_n3420_38528# VSS 2.03238f 
C5690 a_n3690_38528# VSS 0.516979f 
C5691 a_n3565_38502# VSS 1.56115f 
C5692 a_n4334_38528# VSS 0.529888f 
C5693 a_n4209_38502# VSS 3.02222f 
C5694 a_2112_39137# VSS 0.414404f 
C5695 comp_n VSS 0.572075f 
C5696 a_1666_39043# VSS 0.909399f 
C5697 a_1169_39043# VSS 0.615041f 
C5698 a_n2302_39072# VSS 0.483504f 
C5699 a_n4064_39072# VSS 1.71497f 
C5700 a_n2946_39072# VSS 0.486447f 
C5701 a_n3420_39072# VSS 2.21329f 
C5702 a_n3690_39392# VSS 0.517965f 
C5703 a_n3565_39304# VSS 1.46077f 
C5704 a_n4334_39392# VSS 0.529516f 
C5705 a_n4209_39304# VSS 3.25318f 
C5706 a_1273_38525# VSS 3.59416f 
C5707 a_1666_39587# VSS 1.1306f 
C5708 a_1169_39587# VSS 0.633906f 
C5709 a_n2302_39866# VSS 0.483537f 
C5710 a_n4064_39616# VSS 2.17927f 
C5711 a_n2946_39866# VSS 0.527929f 
C5712 a_n3420_39616# VSS 2.11278f 
C5713 a_n3690_39616# VSS 0.574329f 
C5714 a_n3565_39590# VSS 2.14063f 
C5715 a_n4334_39616# VSS 0.529903f 
C5716 a_n4209_39590# VSS 4.08248f 
C5717 a_n2302_40160# VSS 0.522244f 
C5718 a_n4064_40160# VSS 3.30536f 
C5719 a_n4334_40480# VSS 0.578721f 
C5720 a_n4315_30879# VSS 5.10714f 
C5721 a_22485_38105# VSS 1.90993f 
C5722 a_22775_42308# VSS 0.602116f 
C5723 a_21613_42308# VSS 0.725532f 
C5724 a_21887_42336# VSS 0.234022f 
C5725 a_21335_42336# VSS 0.259392f 
C5726 a_7174_31319# VSS 5.511971f 
C5727 a_20712_42282# VSS 0.349662f 
C5728 a_20107_42308# VSS 0.344464f 
C5729 a_13258_32519# VSS 6.35834f 
C5730 a_19647_42308# VSS 0.313304f 
C5731 a_19511_42282# VSS 0.751141f 
C5732 a_19332_42282# VSS 0.31505f 
C5733 a_18907_42674# VSS 0.209311f 
C5734 a_18727_42674# VSS 0.233526f 
C5735 a_18057_42282# VSS 0.370712f 
C5736 a_17531_42308# VSS 0.253358f 
C5737 a_17303_42282# VSS 1.19776f 
C5738 a_4958_30871# VSS 5.01459f 
C5739 a_17124_42282# VSS 0.332693f 
C5740 a_15890_42674# VSS 0.180637f 
C5741 a_15959_42545# VSS 0.263128f 
C5742 a_15803_42450# VSS 0.566963f 
C5743 a_15764_42576# VSS 0.298494f 
C5744 a_15486_42560# VSS 0.263746f 
C5745 a_15051_42282# VSS 0.790649f 
C5746 a_14113_42308# VSS 1.42448f 
C5747 a_14456_42282# VSS 0.33927f 
C5748 a_13575_42558# VSS 0.370369f 
C5749 a_13070_42354# VSS 0.222095f 
C5750 a_12563_42308# VSS 0.330976f 
C5751 a_11551_42558# VSS 0.372919f 
C5752 a_5742_30871# VSS 8.19336f 
C5753 a_11323_42473# VSS 0.253445f 
C5754 a_10723_42308# VSS 0.342975f 
C5755 a_10533_42308# VSS 0.310658f 
C5756 a_9803_42558# VSS 0.370474f 
C5757 a_9223_42460# VSS 0.236204f 
C5758 a_8791_42308# VSS 0.301f 
C5759 a_8685_42308# VSS 0.163732f 
C5760 a_8325_42308# VSS 0.316205f 
C5761 a_8515_42308# VSS 0.250762f 
C5762 a_5934_30871# VSS 5.17377f 
C5763 a_7963_42308# VSS 0.256292f 
C5764 a_6123_31319# VSS 5.02387f 
C5765 a_7227_42308# VSS 0.359705f 
C5766 a_6761_42308# VSS 0.447596f 
C5767 a_5932_42308# VSS 5.11988f 
C5768 a_6171_42473# VSS 0.257988f 
C5769 a_5755_42308# VSS 0.314735f 
C5770 a_4921_42308# VSS 0.511258f 
C5771 a_5379_42460# VSS 0.564806f 
C5772 a_5267_42460# VSS 0.204309f 
C5773 a_3823_42558# VSS 0.381485f 
C5774 a_3318_42354# VSS 0.238394f 
C5775 a_2903_42308# VSS 0.340659f 
C5776 a_2713_42308# VSS 0.31991f 
C5777 a_2351_42308# VSS 0.210162f 
C5778 a_2123_42473# VSS 0.21778f 
C5779 a_1755_42282# VSS 3.17706f 
C5780 a_1606_42308# VSS 5.25671f 
C5781 a_961_42354# VSS 0.215753f 
C5782 a_1184_42692# VSS 0.222827f 
C5783 a_1576_42282# VSS 0.327109f 
C5784 a_1067_42314# VSS 0.32917f 
C5785 a_n1794_35242# VSS 10.0162f 
C5786 a_564_42282# VSS 0.36802f 
C5787 a_n3674_37592# VSS 3.04613f 
C5788 a_n784_42308# VSS 6.50157f 
C5789 a_196_42282# VSS 0.343186f 
C5790 a_n473_42460# VSS 0.366068f 
C5791 a_n961_42308# VSS 0.328065f 
C5792 a_n1329_42308# VSS 0.30898f 
C5793 COMP_P VSS 10.9891f 
C5794 a_n4318_37592# VSS 1.00428f 
C5795 a_n1736_42282# VSS 0.320711f 
C5796 a_n3674_38216# VSS 1.68571f 
C5797 a_n2104_42282# VSS 0.346472f 
C5798 a_n4318_38216# VSS 0.964502f 
C5799 a_n2472_42282# VSS 0.335792f 
C5800 a_n3674_38680# VSS 0.881032f 
C5801 a_n2840_42282# VSS 0.343361f 
C5802 a_14097_32519# VSS 1.90783f 
C5803 a_22400_42852# VSS 1.97851f 
C5804 a_20256_43172# VSS 0.192089f 
C5805 a_14635_42282# VSS 0.336817f 
C5806 a_13291_42460# VSS 0.197331f 
C5807 a_n2293_42282# VSS 2.62914f 
C5808 a_22959_42860# VSS 0.34332f 
C5809 a_22223_42860# VSS 0.328988f 
C5810 a_22165_42308# VSS 0.354098f 
C5811 a_21671_42860# VSS 0.316857f 
C5812 a_21195_42852# VSS 0.277519f 
C5813 a_21356_42826# VSS 0.304166f 
C5814 a_20922_43172# VSS 0.266814f 
C5815 a_19987_42826# VSS 0.378798f 
C5816 a_19164_43230# VSS 0.264863f 
C5817 a_19339_43156# VSS 0.471496f 
C5818 a_18599_43230# VSS 0.266382f 
C5819 a_18817_42826# VSS 0.182139f 
C5820 a_18249_42858# VSS 0.302863f 
C5821 a_17333_42852# VSS 0.29982f 
C5822 a_18083_42858# VSS 0.578693f 
C5823 a_17701_42308# VSS 0.179963f 
C5824 a_17595_43084# VSS 0.205109f 
C5825 a_16795_42852# VSS 0.362281f 
C5826 a_16414_43172# VSS 0.270304f 
C5827 a_15567_42826# VSS 0.316627f 
C5828 a_5342_30871# VSS 4.18155f 
C5829 a_15279_43071# VSS 0.248252f 
C5830 a_5534_30871# VSS 4.58471f 
C5831 a_14543_43071# VSS 0.246071f 
C5832 a_13460_43230# VSS 0.259861f 
C5833 a_13635_43156# VSS 0.7696f 
C5834 a_12895_43230# VSS 0.250159f 
C5835 a_13113_42826# VSS 0.174096f 
C5836 a_12545_42858# VSS 0.287468f 
C5837 a_12089_42308# VSS 0.283874f 
C5838 a_12379_42858# VSS 0.549229f 
C5839 a_10341_42308# VSS 0.317389f 
C5840 a_10922_42852# VSS 0.176112f 
C5841 a_10991_42826# VSS 0.261283f 
C5842 a_10796_42968# VSS 0.29877f 
C5843 a_10835_43094# VSS 0.59174f 
C5844 a_10518_42984# VSS 0.260322f 
C5845 a_10083_42826# VSS 0.762957f 
C5846 a_8952_43230# VSS 0.261046f 
C5847 a_9127_43156# VSS 0.77314f 
C5848 a_8387_43230# VSS 0.255573f 
C5849 a_8605_42826# VSS 0.181157f 
C5850 a_8037_42858# VSS 0.293593f 
C5851 a_7765_42852# VSS 0.252651f 
C5852 a_7871_42858# VSS 0.503534f 
C5853 a_7227_42852# VSS 0.36607f 
C5854 a_5755_42852# VSS 0.383967f 
C5855 a_5111_42852# VSS 0.354197f 
C5856 a_4520_42826# VSS 0.334784f 
C5857 a_3935_42891# VSS 0.26911f 
C5858 a_3681_42891# VSS 0.301094f 
C5859 a_2905_42968# VSS 0.305424f 
C5860 a_2075_43172# VSS 0.537699f 
C5861 a_1847_42826# VSS 0.670072f 
C5862 a_791_42968# VSS 0.335942f 
C5863 a_685_42968# VSS 0.220885f 
C5864 a_n4318_38680# VSS 1.39087f 
C5865 a_n3674_39304# VSS 1.06639f 
C5866 a_n13_43084# VSS 0.368998f 
C5867 a_n1076_43230# VSS 0.263204f 
C5868 a_n901_43156# VSS 0.76245f 
C5869 a_n1641_43230# VSS 0.256397f 
C5870 a_n1423_42826# VSS 0.1805f 
C5871 a_n1991_42858# VSS 0.295941f 
C5872 a_n1853_43023# VSS 1.30078f 
C5873 a_n2157_42858# VSS 0.556569f 
C5874 a_n2472_42826# VSS 0.301801f 
C5875 a_n2840_42826# VSS 0.327636f 
C5876 a_20749_43396# VSS 0.253248f 
C5877 a_17364_32525# VSS 1.89103f 
C5878 a_22959_43396# VSS 0.345439f 
C5879 a_14209_32519# VSS 2.01016f 
C5880 a_22591_43396# VSS 0.335697f 
C5881 a_13887_32519# VSS 1.94312f 
C5882 a_22223_43396# VSS 0.333609f 
C5883 a_5649_42852# VSS 1.95364f 
C5884 a_13678_32519# VSS 2.06126f 
C5885 a_21855_43396# VSS 0.334538f 
C5886 a_4361_42308# VSS 1.30251f 
C5887 a_13467_32519# VSS 2.22551f 
C5888 a_19095_43396# VSS 0.132304f 
C5889 a_21487_43396# VSS 0.293844f 
C5890 a_743_42282# VSS 1.36822f 
C5891 a_4190_30871# VSS 7.379981f 
C5892 a_21259_43561# VSS 0.217667f 
C5893 a_16823_43084# VSS 1.23251f 
C5894 a_19700_43370# VSS 0.335707f 
C5895 a_19268_43646# VSS 0.242693f 
C5896 a_15743_43084# VSS 1.49489f 
C5897 a_18783_43370# VSS 0.360096f 
C5898 a_18525_43370# VSS 0.361236f 
C5899 a_18429_43548# VSS 0.222219f 
C5900 a_17324_43396# VSS 0.258017f 
C5901 a_17499_43370# VSS 0.762886f 
C5902 a_16759_43396# VSS 0.252915f 
C5903 a_16977_43638# VSS 0.178776f 
C5904 a_16409_43396# VSS 0.290743f 
C5905 a_16547_43609# VSS 0.561468f 
C5906 a_16243_43396# VSS 0.562369f 
C5907 a_16137_43396# VSS 0.635905f 
C5908 a_15781_43660# VSS 0.234761f 
C5909 a_15681_43442# VSS 0.20154f 
C5910 a_12281_43396# VSS 0.691406f 
C5911 a_10341_43396# VSS 0.796012f 
C5912 a_14955_43396# VSS 0.266041f 
C5913 a_15095_43370# VSS 0.436411f 
C5914 a_14205_43396# VSS 0.2933f 
C5915 a_14358_43442# VSS 0.198188f 
C5916 a_14579_43548# VSS 0.293668f 
C5917 a_13667_43396# VSS 0.265557f 
C5918 a_10695_43548# VSS 0.279385f 
C5919 a_9803_43646# VSS 0.371929f 
C5920 a_9145_43396# VSS 0.437647f 
C5921 a_8685_43396# VSS 1.0146f 
C5922 a_3457_43396# VSS 0.379621f 
C5923 a_2813_43396# VSS 0.412407f 
C5924 a_9396_43370# VSS 0.338475f 
C5925 a_8791_43396# VSS 0.235222f 
C5926 a_8147_43396# VSS 0.256103f 
C5927 a_7112_43396# VSS 0.256956f 
C5928 a_7287_43370# VSS 0.754599f 
C5929 a_6547_43396# VSS 0.253718f 
C5930 a_6765_43638# VSS 0.174622f 
C5931 a_6197_43396# VSS 0.290517f 
C5932 a_6293_42852# VSS 0.473619f 
C5933 a_6031_43396# VSS 0.541083f 
C5934 a_648_43396# VSS 0.231254f 
C5935 a_3539_42460# VSS 0.337918f 
C5936 a_3626_43646# VSS 1.9807f 
C5937 a_2982_43646# VSS 3.25953f 
C5938 a_n1557_42282# VSS 0.870257f 
C5939 a_4905_42826# VSS 0.781685f 
C5940 a_3080_42308# VSS 5.07266f 
C5941 a_4699_43561# VSS 0.267684f 
C5942 a_4235_43370# VSS 0.33553f 
C5943 a_4093_43548# VSS 0.320586f 
C5944 a_1756_43548# VSS 0.322408f 
C5945 a_1568_43370# VSS 0.63594f 
C5946 a_1049_43396# VSS 0.216408f 
C5947 a_1209_43370# VSS 0.281234f 
C5948 a_458_43396# VSS 0.252302f 
C5949 a_104_43370# VSS 0.297328f 
C5950 a_n97_42460# VSS 6.9914f 
C5951 a_n447_43370# VSS 0.269574f 
C5952 a_n1352_43396# VSS 0.260107f 
C5953 a_n1177_43370# VSS 0.478516f 
C5954 a_n1917_43396# VSS 0.258245f 
C5955 a_n1699_43638# VSS 0.175452f 
C5956 a_n2267_43396# VSS 0.297246f 
C5957 a_n2129_43609# VSS 1.07965f 
C5958 a_n2433_43396# VSS 0.56533f 
C5959 a_n4318_39304# VSS 0.959585f 
C5960 a_n2840_43370# VSS 0.316787f 
C5961 a_17538_32519# VSS 1.88845f 
C5962 a_20974_43370# VSS 0.458091f 
C5963 a_14401_32519# VSS 2.32028f 
C5964 a_21381_43940# VSS 0.358332f 
C5965 a_19319_43548# VSS 0.229395f 
C5966 a_14021_43940# VSS 0.387813f 
C5967 a_11173_44260# VSS 0.219946f 
C5968 a_10555_44260# VSS 0.346315f 
C5969 a_22959_43948# VSS 0.341565f 
C5970 a_15493_43940# VSS 0.460801f 
C5971 a_22223_43948# VSS 0.31992f 
C5972 a_11341_43940# VSS 0.365183f 
C5973 a_21115_43940# VSS 0.204633f 
C5974 a_20935_43940# VSS 0.222887f 
C5975 a_20623_43914# VSS 0.371294f 
C5976 a_20365_43914# VSS 0.359455f 
C5977 a_20269_44172# VSS 0.225063f 
C5978 a_19862_44208# VSS 0.562087f 
C5979 a_19478_44306# VSS 0.278384f 
C5980 a_15493_43396# VSS 0.277875f 
C5981 a_19328_44172# VSS 0.2031f 
C5982 a_18451_43940# VSS 0.377396f 
C5983 a_18326_43940# VSS 0.276559f 
C5984 a_18079_43940# VSS 0.21121f 
C5985 a_17973_43940# VSS 0.359917f 
C5986 a_17737_43940# VSS 0.386318f 
C5987 a_15682_43940# VSS 1.9643f 
C5988 a_14955_43940# VSS 0.365393f 
C5989 a_13483_43940# VSS 0.376442f 
C5990 a_12429_44172# VSS 0.389129f 
C5991 a_11750_44172# VSS 0.221782f 
C5992 a_10807_43548# VSS 0.451031f 
C5993 a_10949_43914# VSS 0.257331f 
C5994 a_10729_43914# VSS 0.34307f 
C5995 a_10405_44172# VSS 0.142993f 
C5996 a_9672_43914# VSS 0.323006f 
C5997 a_9028_43914# VSS 0.398016f 
C5998 a_8333_44056# VSS 0.331632f 
C5999 a_n2661_42282# VSS 1.51789f 
C6000 a_3499_42826# VSS 0.380221f 
C6001 a_n3674_39768# VSS 0.890487f 
C6002 a_n4318_39768# VSS 1.09976f 
C6003 a_7845_44172# VSS 0.239173f 
C6004 a_7542_44172# VSS 0.283767f 
C6005 a_7281_43914# VSS 0.271121f 
C6006 a_6453_43914# VSS 0.26639f 
C6007 a_5663_43940# VSS 0.488325f 
C6008 a_5495_43940# VSS 0.212229f 
C6009 a_5013_44260# VSS 0.279924f 
C6010 a_5244_44056# VSS 0.216368f 
C6011 a_3905_42865# VSS 0.9893f 
C6012 a_3600_43914# VSS 0.422049f 
C6013 a_2998_44172# VSS 0.503048f 
C6014 a_2889_44172# VSS 0.217034f 
C6015 a_2675_43914# VSS 0.2974f 
C6016 a_895_43940# VSS 0.237723f 
C6017 a_2479_44172# VSS 0.817462f 
C6018 a_2127_44172# VSS 0.517911f 
C6019 a_453_43940# VSS 0.285192f 
C6020 a_1414_42308# VSS 1.07452f 
C6021 a_1467_44172# VSS 0.187431f 
C6022 a_1115_44172# VSS 0.52592f 
C6023 a_644_44056# VSS 0.227493f 
C6024 a_175_44278# VSS 0.226801f 
C6025 a_n984_44318# VSS 0.27358f 
C6026 a_n809_44244# VSS 0.785904f 
C6027 a_n1549_44318# VSS 0.264547f 
C6028 a_n1331_43914# VSS 0.185087f 
C6029 a_n1899_43946# VSS 0.299008f 
C6030 a_n1761_44111# VSS 0.392075f 
C6031 a_n2065_43946# VSS 0.658803f 
C6032 a_n2472_43914# VSS 0.3103f 
C6033 a_n2840_43914# VSS 0.345355f 
C6034 a_19237_31679# VSS 1.4857f 
C6035 a_22959_44484# VSS 0.343897f 
C6036 a_17730_32519# VSS 2.45467f 
C6037 a_22591_44484# VSS 0.315361f 
C6038 a_22485_44484# VSS 0.590119f 
C6039 a_20512_43084# VSS 0.561552f 
C6040 a_22315_44484# VSS 0.238239f 
C6041 a_3422_30871# VSS 9.021831f 
C6042 a_18579_44172# VSS 0.812679f 
C6043 a_19279_43940# VSS 1.69633f 
C6044 a_20766_44850# VSS 0.177656f 
C6045 a_20835_44721# VSS 0.260406f 
C6046 a_20679_44626# VSS 0.58931f 
C6047 a_20640_44752# VSS 0.296084f 
C6048 a_20362_44736# VSS 0.255907f 
C6049 a_20159_44458# VSS 0.483669f 
C6050 a_19615_44636# VSS 0.238459f 
C6051 a_11967_42832# VSS 6.11191f 
C6052 a_17517_44484# VSS 0.244051f 
C6053 a_14673_44172# VSS 0.290001f 
C6054 a_11541_44484# VSS 0.139071f 
C6055 a_15433_44458# VSS 0.301508f 
C6056 a_14815_43914# VSS 0.445698f 
C6057 a_n2293_43922# VSS 3.31971f 
C6058 a_n2661_43922# VSS 1.51991f 
C6059 a_n2661_42834# VSS 1.20196f 
C6060 a_9159_44484# VSS 0.158168f 
C6061 a_10617_44484# VSS 0.119149f 
C6062 a_5708_44484# VSS 0.231649f 
C6063 a_3363_44484# VSS 0.27629f 
C6064 a_556_44484# VSS 0.201935f 
C6065 a_9313_44734# VSS 1.31461f 
C6066 a_5891_43370# VSS 2.82295f 
C6067 a_8375_44464# VSS 0.211867f 
C6068 a_7640_43914# VSS 0.542377f 
C6069 a_6109_44484# VSS 0.648821f 
C6070 a_n23_44458# VSS 0.278255f 
C6071 a_n356_44636# VSS 2.91333f 
C6072 a_18989_43940# VSS 0.423174f 
C6073 a_18374_44850# VSS 0.179731f 
C6074 a_18443_44721# VSS 0.253971f 
C6075 a_18287_44626# VSS 0.507939f 
C6076 a_18248_44752# VSS 0.294917f 
C6077 a_17970_44736# VSS 0.26161f 
C6078 a_17767_44458# VSS 0.474097f 
C6079 a_16979_44734# VSS 0.363013f 
C6080 a_14539_43914# VSS 1.18088f 
C6081 a_16112_44458# VSS 0.326339f 
C6082 a_15004_44636# VSS 0.254778f 
C6083 a_13720_44458# VSS 0.403209f 
C6084 a_13076_44458# VSS 0.38829f 
C6085 a_12883_44458# VSS 0.287544f 
C6086 a_12607_44458# VSS 0.499331f 
C6087 a_8975_43940# VSS 0.652857f 
C6088 a_10057_43914# VSS 0.654189f 
C6089 a_10440_44484# VSS 0.210149f 
C6090 a_10334_44484# VSS 0.210217f 
C6091 a_10157_44484# VSS 0.208916f 
C6092 a_9838_44484# VSS 0.276258f 
C6093 a_5883_43914# VSS 0.792825f 
C6094 a_8701_44490# VSS 0.358059f 
C6095 a_8103_44636# VSS 0.340824f 
C6096 a_6298_44484# VSS 1.93814f 
C6097 a_5518_44484# VSS 0.242995f 
C6098 a_5343_44458# VSS 1.28071f 
C6099 a_4743_44484# VSS 0.327178f 
C6100 a_n699_43396# VSS 1.82142f 
C6101 a_4223_44672# VSS 0.659279f 
C6102 a_2779_44458# VSS 0.532137f 
C6103 a_949_44458# VSS 1.97734f 
C6104 a_742_44458# VSS 1.02263f 
C6105 a_n452_44636# VSS 0.254732f 
C6106 a_n1352_44484# VSS 0.269853f 
C6107 a_n1177_44458# VSS 0.493891f 
C6108 a_n1917_44484# VSS 0.280038f 
C6109 a_n1699_44726# VSS 0.197478f 
C6110 a_n2267_44484# VSS 0.308908f 
C6111 a_n2129_44697# VSS 0.307327f 
C6112 a_n2433_44484# VSS 0.679598f 
C6113 a_n2661_44458# VSS 0.487677f 
C6114 a_n4318_40392# VSS 0.995833f 
C6115 a_n2840_44458# VSS 0.316322f 
C6116 a_19721_31679# VSS 1.61938f 
C6117 a_18114_32519# VSS 3.11986f 
C6118 a_20193_45348# VSS 1.70015f 
C6119 a_11691_44458# VSS 1.78467f 
C6120 a_19113_45348# VSS 0.367248f 
C6121 a_22959_45036# VSS 0.345334f 
C6122 a_22223_45036# VSS 0.354178f 
C6123 a_11827_44484# VSS 1.28091f 
C6124 a_21359_45002# VSS 0.397791f 
C6125 a_21101_45002# VSS 0.35202f 
C6126 a_21005_45260# VSS 0.212992f 
C6127 a_20567_45036# VSS 0.31908f 
C6128 a_18494_42460# VSS 1.15626f 
C6129 a_18184_42460# VSS 0.838573f 
C6130 a_19778_44110# VSS 0.599421f 
C6131 a_18911_45144# VSS 0.307008f 
C6132 a_18587_45118# VSS 0.214925f 
C6133 a_18315_45260# VSS 0.334834f 
C6134 a_17719_45144# VSS 0.331229f 
C6135 a_17613_45144# VSS 0.244364f 
C6136 a_17023_45118# VSS 0.20885f 
C6137 a_16922_45042# VSS 0.818675f 
C6138 a_n2661_43370# VSS 0.820606f 
C6139 a_8560_45348# VSS 0.185033f 
C6140 a_n2293_42834# VSS 1.1151f 
C6141 a_2304_45348# VSS 0.182367f 
C6142 a_1423_45028# VSS 0.980773f 
C6143 a_626_44172# VSS 0.67926f 
C6144 a_375_42282# VSS 0.447027f 
C6145 a_16751_45260# VSS 0.316547f 
C6146 a_1307_43914# VSS 2.30311f 
C6147 a_16019_45002# VSS 0.25377f 
C6148 a_15595_45028# VSS 0.214111f 
C6149 a_15415_45028# VSS 0.221991f 
C6150 a_14797_45144# VSS 0.249222f 
C6151 a_14537_43396# VSS 1.73146f 
C6152 a_14180_45002# VSS 0.327485f 
C6153 a_13777_45326# VSS 0.272936f 
C6154 a_13556_45296# VSS 1.01916f 
C6155 a_9482_43914# VSS 3.42654f 
C6156 a_13348_45260# VSS 0.243533f 
C6157 a_13159_45002# VSS 0.265737f 
C6158 a_13017_45260# VSS 0.362048f 
C6159 a_11963_45334# VSS 0.226884f 
C6160 a_11787_45002# VSS 0.212512f 
C6161 a_10951_45334# VSS 0.228638f 
C6162 a_10775_45002# VSS 0.204487f 
C6163 a_8953_45002# VSS 1.94941f 
C6164 a_8191_45002# VSS 0.325964f 
C6165 a_7705_45326# VSS 0.273009f 
C6166 a_6709_45028# VSS 0.354418f 
C6167 a_7229_43940# VSS 0.786182f 
C6168 a_7276_45260# VSS 0.251523f 
C6169 a_5205_44484# VSS 0.546179f 
C6170 a_6431_45366# VSS 0.233718f 
C6171 a_6171_45002# VSS 0.700605f 
C6172 a_3232_43370# VSS 2.99721f 
C6173 a_5691_45260# VSS 0.370273f 
C6174 a_4927_45028# VSS 0.520892f 
C6175 a_5111_44636# VSS 3.44603f 
C6176 a_5147_45002# VSS 0.803306f 
C6177 a_4558_45348# VSS 0.446148f 
C6178 a_4574_45260# VSS 0.208274f 
C6179 a_3537_45260# VSS 2.45782f 
C6180 a_3429_45260# VSS 0.274034f 
C6181 a_3065_45002# VSS 0.864786f 
C6182 a_2680_45002# VSS 0.321351f 
C6183 a_2382_45260# VSS 1.03422f 
C6184 a_2274_45254# VSS 0.187307f 
C6185 a_1667_45002# VSS 0.345429f 
C6186 a_327_44734# VSS 0.419171f 
C6187 a_413_45260# VSS 4.87522f 
C6188 a_n37_45144# VSS 0.321746f 
C6189 a_n143_45144# VSS 0.209896f 
C6190 a_n467_45028# VSS 0.311181f 
C6191 a_n967_45348# VSS 0.453992f 
C6192 en_comp VSS 7.84057f 
C6193 a_n2956_37592# VSS 2.90302f 
C6194 a_n2810_45028# VSS 1.52635f 
C6195 a_n745_45366# VSS 0.257282f 
C6196 a_n913_45002# VSS 5.04725f 
C6197 a_n1059_45260# VSS 2.30619f 
C6198 a_n2017_45002# VSS 1.09013f 
C6199 a_n2109_45247# VSS 0.252392f 
C6200 a_n2293_45010# VSS 0.614925f 
C6201 a_n2472_45002# VSS 0.298945f 
C6202 a_n2661_45010# VSS 0.839496f 
C6203 a_n2840_45002# VSS 0.340687f 
C6204 a_20447_31679# VSS 1.49249f 
C6205 a_22959_45572# VSS 0.34535f 
C6206 a_19963_31679# VSS 1.43879f 
C6207 a_22591_45572# VSS 0.363695f 
C6208 a_3357_43084# VSS 2.42707f 
C6209 a_19479_31679# VSS 1.67279f 
C6210 a_22223_45572# VSS 0.334964f 
C6211 a_2437_43646# VSS 6.25635f 
C6212 a_21513_45002# VSS 0.669089f 
C6213 a_21188_45572# VSS 0.284872f 
C6214 a_21363_45546# VSS 0.515994f 
C6215 a_20623_45572# VSS 0.256236f 
C6216 a_20841_45814# VSS 0.180037f 
C6217 a_20273_45572# VSS 0.288513f 
C6218 a_20107_45572# VSS 0.541125f 
C6219 a_17668_45572# VSS 0.217142f 
C6220 a_19256_45572# VSS 0.257674f 
C6221 a_19431_45546# VSS 0.487121f 
C6222 a_18691_45572# VSS 0.255356f 
C6223 a_18909_45814# VSS 0.178658f 
C6224 a_18341_45572# VSS 0.291608f 
C6225 a_18479_45785# VSS 1.15946f 
C6226 a_18175_45572# VSS 0.516981f 
C6227 a_16147_45260# VSS 0.506229f 
C6228 a_17478_45572# VSS 0.232341f 
C6229 a_15861_45028# VSS 0.449058f 
C6230 a_8696_44636# VSS 0.917254f 
C6231 a_16680_45572# VSS 0.258674f 
C6232 a_16855_45546# VSS 0.471485f 
C6233 a_16115_45572# VSS 0.253972f 
C6234 a_16333_45814# VSS 0.178165f 
C6235 a_15765_45572# VSS 0.291326f 
C6236 a_15903_45785# VSS 0.4164f 
C6237 a_15599_45572# VSS 0.50233f 
C6238 a_15037_45618# VSS 0.209713f 
C6239 a_11136_45572# VSS 0.17156f 
C6240 a_9159_45572# VSS 0.151638f 
C6241 a_8192_45572# VSS 0.17002f 
C6242 a_10907_45822# VSS 0.547001f 
C6243 a_15143_45578# VSS 0.315994f 
C6244 a_14495_45572# VSS 0.325874f 
C6245 a_13249_42308# VSS 1.08648f 
C6246 a_13904_45546# VSS 0.327907f 
C6247 a_13527_45546# VSS 0.245514f 
C6248 a_13163_45724# VSS 0.180841f 
C6249 a_12791_45546# VSS 0.237787f 
C6250 a_11823_42460# VSS 2.45644f 
C6251 a_12427_45724# VSS 0.190531f 
C6252 a_11962_45724# VSS 0.218739f 
C6253 a_11652_45724# VSS 0.258015f 
C6254 a_11525_45546# VSS 0.346102f 
C6255 a_11322_45546# VSS 0.62914f 
C6256 a_10490_45724# VSS 0.972668f 
C6257 a_8746_45002# VSS 0.547616f 
C6258 a_10193_42453# VSS 3.59848f 
C6259 a_10180_45724# VSS 0.281135f 
C6260 a_10053_45546# VSS 0.373668f 
C6261 a_9049_44484# VSS 0.249658f 
C6262 a_7499_43078# VSS 3.22587f 
C6263 a_8568_45546# VSS 0.317032f 
C6264 a_8162_45546# VSS 0.376225f 
C6265 a_4880_45572# VSS 0.182839f 
C6266 a_3775_45552# VSS 0.209244f 
C6267 a_7227_45028# VSS 0.439395f 
C6268 a_6598_45938# VSS 0.185967f 
C6269 a_6667_45809# VSS 0.264656f 
C6270 a_6511_45714# VSS 0.647716f 
C6271 a_6472_45840# VSS 0.310105f 
C6272 a_6194_45824# VSS 0.2717f 
C6273 a_5907_45546# VSS 0.592148f 
C6274 a_5263_45724# VSS 0.250928f 
C6275 a_4099_45572# VSS 0.33915f 
C6276 a_2711_45572# VSS 1.77517f 
C6277 a_2277_45546# VSS 0.303704f 
C6278 a_1609_45822# VSS 0.5528f 
C6279 a_n443_42852# VSS 4.64762f 
C6280 a_n23_45546# VSS 0.281189f 
C6281 a_n356_45724# VSS 0.32306f 
C6282 a_3503_45724# VSS 0.322319f 
C6283 a_3316_45546# VSS 0.336134f 
C6284 a_3218_45724# VSS 0.379893f 
C6285 a_2957_45546# VSS 0.276358f 
C6286 a_1848_45724# VSS 0.245258f 
C6287 a_997_45618# VSS 0.248122f 
C6288 a_n755_45592# VSS 5.8889f 
C6289 a_n357_42282# VSS 2.46134f 
C6290 a_310_45028# VSS 0.207165f 
C6291 a_n1099_45572# VSS 0.339525f 
C6292 a_380_45546# VSS 0.337145f 
C6293 a_n452_45724# VSS 0.253614f 
C6294 a_n863_45724# VSS 3.49288f 
C6295 a_n1079_45724# VSS 0.289271f 
C6296 a_n2293_45546# VSS 0.879703f 
C6297 a_n2956_38216# VSS 1.49846f 
C6298 a_n2472_45546# VSS 0.340801f 
C6299 a_n2661_45546# VSS 1.58481f 
C6300 a_n2810_45572# VSS 1.43198f 
C6301 a_n2840_45546# VSS 0.344757f 
C6302 a_20692_30879# VSS 1.6166f 
C6303 a_20205_31679# VSS 1.45868f 
C6304 a_16375_45002# VSS 1.44161f 
C6305 a_13259_45724# VSS 4.49032f 
C6306 a_12638_46436# VSS 0.162178f 
C6307 a_12379_46436# VSS 0.275423f 
C6308 a_10586_45546# VSS 0.542658f 
C6309 a_8049_45260# VSS 0.741927f 
C6310 a_8034_45724# VSS 0.299594f 
C6311 a_5066_45546# VSS 0.436834f 
C6312 a_n1925_42282# VSS 1.34109f 
C6313 a_526_44458# VSS 6.44493f 
C6314 a_n2956_38680# VSS 1.34225f 
C6315 a_n2956_39304# VSS 1.60721f 
C6316 a_22959_46124# VSS 0.345245f 
C6317 a_10809_44734# VSS 1.05002f 
C6318 a_22223_46124# VSS 0.354467f 
C6319 a_6945_45028# VSS 0.978274f 
C6320 a_21137_46414# VSS 0.340736f 
C6321 a_20708_46348# VSS 0.268156f 
C6322 a_19900_46494# VSS 0.26164f 
C6323 a_20075_46420# VSS 0.475201f 
C6324 a_19335_46494# VSS 0.260378f 
C6325 a_19553_46090# VSS 0.179968f 
C6326 a_18985_46122# VSS 0.297132f 
C6327 a_18819_46122# VSS 0.545109f 
C6328 a_17957_46116# VSS 0.309446f 
C6329 a_18189_46348# VSS 0.296366f 
C6330 a_17715_44484# VSS 0.55862f 
C6331 a_17583_46090# VSS 0.307562f 
C6332 a_15682_46116# VSS 1.96743f 
C6333 a_2324_44458# VSS 6.12227f 
C6334 a_14840_46494# VSS 0.263367f 
C6335 a_15015_46420# VSS 0.472948f 
C6336 a_14275_46494# VSS 0.258968f 
C6337 a_14493_46090# VSS 0.176122f 
C6338 a_13925_46122# VSS 0.294602f 
C6339 a_13759_46122# VSS 0.518292f 
C6340 a_13351_46090# VSS 0.304427f 
C6341 a_12594_46348# VSS 0.284494f 
C6342 a_12005_46116# VSS 0.381711f 
C6343 a_10903_43370# VSS 2.66576f 
C6344 a_11387_46155# VSS 0.260117f 
C6345 a_11133_46155# VSS 0.299642f 
C6346 a_11189_46129# VSS 0.32558f 
C6347 a_9290_44172# VSS 4.78398f 
C6348 a_10355_46116# VSS 0.290668f 
C6349 a_9823_46155# VSS 0.261206f 
C6350 a_9569_46155# VSS 0.304755f 
C6351 a_9625_46129# VSS 0.369694f 
C6352 a_8953_45546# VSS 1.00397f 
C6353 a_5937_45572# VSS 1.8333f 
C6354 a_8199_44636# VSS 2.29742f 
C6355 a_8349_46414# VSS 0.273442f 
C6356 a_8016_46348# VSS 0.539696f 
C6357 a_7920_46348# VSS 0.269852f 
C6358 a_6419_46155# VSS 0.273686f 
C6359 a_6165_46155# VSS 0.303989f 
C6360 a_5497_46414# VSS 0.304684f 
C6361 a_5204_45822# VSS 0.338817f 
C6362 a_5164_46348# VSS 0.419282f 
C6363 a_5068_46348# VSS 0.25855f 
C6364 a_4704_46090# VSS 0.296767f 
C6365 a_4419_46090# VSS 0.357571f 
C6366 a_4185_45028# VSS 2.50496f 
C6367 a_3699_46348# VSS 0.226584f 
C6368 a_3483_46348# VSS 4.80498f 
C6369 a_3147_46376# VSS 0.52775f 
C6370 a_2804_46116# VSS 0.222855f 
C6371 a_2698_46116# VSS 0.215567f 
C6372 a_2521_46116# VSS 0.220999f 
C6373 a_167_45260# VSS 1.32487f 
C6374 a_2202_46116# VSS 0.273578f 
C6375 a_1823_45246# VSS 2.36307f 
C6376 a_1138_42852# VSS 0.456566f 
C6377 a_1176_45822# VSS 0.278365f 
C6378 a_1208_46090# VSS 0.348206f 
C6379 a_805_46414# VSS 0.27506f 
C6380 a_472_46348# VSS 0.32751f 
C6381 a_376_46348# VSS 0.285607f 
C6382 a_n1076_46494# VSS 0.262147f 
C6383 a_n901_46420# VSS 0.762523f 
C6384 a_n1641_46494# VSS 0.256945f 
C6385 a_n1423_46090# VSS 0.176189f 
C6386 a_n1991_46122# VSS 0.305274f 
C6387 a_n1853_46287# VSS 0.341802f 
C6388 a_n2157_46122# VSS 0.525314f 
C6389 a_n2293_46098# VSS 0.690447f 
C6390 a_n2472_46090# VSS 0.290925f 
C6391 a_n2840_46090# VSS 0.340313f 
C6392 a_21076_30879# VSS 2.09664f 
C6393 a_22959_46660# VSS 0.338967f 
C6394 a_12741_44636# VSS 0.979225f 
C6395 a_20820_30879# VSS 1.68221f 
C6396 a_22591_46660# VSS 0.292786f 
C6397 a_11415_45002# VSS 1.63684f 
C6398 a_20202_43084# VSS 1.05073f 
C6399 a_22365_46825# VSS 0.208388f 
C6400 a_18280_46660# VSS 0.29316f 
C6401 a_17639_46660# VSS 0.308795f 
C6402 a_22000_46634# VSS 0.295895f 
C6403 a_21188_46660# VSS 0.261124f 
C6404 a_21363_46634# VSS 0.488515f 
C6405 a_20623_46660# VSS 0.258464f 
C6406 a_20841_46902# VSS 0.180869f 
C6407 a_20273_46660# VSS 0.309206f 
C6408 a_20411_46873# VSS 0.393328f 
C6409 a_20107_46660# VSS 0.575208f 
C6410 a_19123_46287# VSS 0.477642f 
C6411 a_18285_46348# VSS 0.577053f 
C6412 a_765_45546# VSS 0.902406f 
C6413 a_17339_46660# VSS 0.927636f 
C6414 a_16721_46634# VSS 0.305539f 
C6415 a_16388_46812# VSS 1.42609f 
C6416 a_13059_46348# VSS 2.36107f 
C6417 a_14513_46634# VSS 0.29862f 
C6418 a_14180_46812# VSS 0.368158f 
C6419 a_14035_46660# VSS 0.322858f 
C6420 a_13885_46660# VSS 0.297377f 
C6421 a_19692_46634# VSS 1.97188f 
C6422 a_19466_46812# VSS 0.675335f 
C6423 a_19333_46634# VSS 0.289568f 
C6424 a_15227_44166# VSS 2.80559f 
C6425 a_18834_46812# VSS 0.198054f 
C6426 a_17609_46634# VSS 0.205547f 
C6427 a_16292_46812# VSS 0.271203f 
C6428 a_15559_46634# VSS 0.394779f 
C6429 a_15368_46634# VSS 0.278142f 
C6430 a_14976_45028# VSS 0.479565f 
C6431 a_3090_45724# VSS 2.6372f 
C6432 a_15009_46634# VSS 0.270859f 
C6433 a_14084_46812# VSS 0.251005f 
C6434 a_13607_46688# VSS 0.218935f 
C6435 a_12816_46660# VSS 0.260317f 
C6436 a_12991_46634# VSS 0.475827f 
C6437 a_12251_46660# VSS 0.270927f 
C6438 a_12469_46902# VSS 0.193369f 
C6439 a_11901_46660# VSS 0.303844f 
C6440 a_11813_46116# VSS 0.563718f 
C6441 a_11735_46660# VSS 0.520568f 
C6442 a_8270_45546# VSS 0.779033f 
C6443 a_6969_46634# VSS 0.289597f 
C6444 a_6755_46942# VSS 3.33348f 
C6445 a_10249_46116# VSS 0.414443f 
C6446 a_10554_47026# VSS 0.191251f 
C6447 a_10623_46897# VSS 0.283572f 
C6448 a_10467_46802# VSS 0.523954f 
C6449 a_10428_46928# VSS 0.314538f 
C6450 a_10150_46912# VSS 0.276624f 
C6451 a_9863_46634# VSS 0.607398f 
C6452 a_8492_46660# VSS 0.283316f 
C6453 a_8667_46634# VSS 0.596387f 
C6454 a_7927_46660# VSS 0.269867f 
C6455 a_8145_46902# VSS 0.179735f 
C6456 a_7577_46660# VSS 0.314978f 
C6457 a_7715_46873# VSS 0.546182f 
C6458 a_7411_46660# VSS 0.532412f 
C6459 a_5257_43370# VSS 1.42323f 
C6460 a_6540_46812# VSS 0.248814f 
C6461 a_5732_46660# VSS 0.260482f 
C6462 a_5907_46634# VSS 0.473347f 
C6463 a_5167_46660# VSS 0.263586f 
C6464 a_5385_46902# VSS 0.17737f 
C6465 a_4817_46660# VSS 0.296797f 
C6466 a_4955_46873# VSS 0.365781f 
C6467 a_4651_46660# VSS 0.548065f 
C6468 a_4646_46812# VSS 2.12519f 
C6469 a_3877_44458# VSS 2.8543f 
C6470 a_3524_46660# VSS 0.267612f 
C6471 a_3699_46634# VSS 0.499647f 
C6472 a_2959_46660# VSS 0.261026f 
C6473 a_3177_46902# VSS 0.184239f 
C6474 a_2609_46660# VSS 0.302878f 
C6475 a_2443_46660# VSS 0.657702f 
C6476 a_n2661_46098# VSS 2.05975f 
C6477 a_1799_45572# VSS 0.30194f 
C6478 a_1983_46706# VSS 0.205951f 
C6479 a_2107_46812# VSS 1.13475f 
C6480 a_948_46660# VSS 0.263413f 
C6481 a_1123_46634# VSS 0.776627f 
C6482 a_383_46660# VSS 0.269735f 
C6483 a_601_46902# VSS 0.192316f 
C6484 a_33_46660# VSS 0.309712f 
C6485 a_171_46873# VSS 0.579977f 
C6486 a_n133_46660# VSS 0.576523f 
C6487 a_n2438_43548# VSS 2.99787f 
C6488 a_n743_46660# VSS 3.29885f 
C6489 a_n1021_46688# VSS 0.271211f 
C6490 a_n1925_46634# VSS 1.33202f 
C6491 a_n2312_38680# VSS 2.0221f 
C6492 a_n2104_46634# VSS 0.340006f 
C6493 a_n2293_46634# VSS 1.52366f 
C6494 a_n2442_46660# VSS 1.32617f 
C6495 a_n2472_46634# VSS 0.323981f 
C6496 a_n2661_46634# VSS 0.742038f 
C6497 a_n2956_39768# VSS 1.30197f 
C6498 a_n2840_46634# VSS 0.328049f 
C6499 a_22612_30879# VSS 3.44331f 
C6500 a_21588_30879# VSS 2.81097f 
C6501 a_20916_46384# VSS 0.827544f 
C6502 a_20843_47204# VSS 0.121976f 
C6503 a_19594_46812# VSS 0.277274f 
C6504 a_19321_45002# VSS 1.15234f 
C6505 a_13747_46662# VSS 2.11905f 
C6506 a_13661_43548# VSS 2.82749f 
C6507 a_5807_45002# VSS 2.5828f 
C6508 a_768_44030# VSS 3.03052f 
C6509 a_12549_44172# VSS 2.68201f 
C6510 a_12891_46348# VSS 1.22195f 
C6511 a_11309_47204# VSS 0.423399f 
C6512 a_9804_47204# VSS 0.528639f 
C6513 a_8128_46384# VSS 0.573494f 
C6514 a_n881_46662# VSS 4.56296f 
C6515 a_n1613_43370# VSS 4.90074f 
C6516 a_2747_46873# VSS 0.287894f 
C6517 a_n2312_39304# VSS 1.49307f 
C6518 a_n2312_40392# VSS 2.25565f 
C6519 a_22959_47212# VSS 0.322938f 
C6520 a_11453_44696# VSS 0.689179f 
C6521 SMPL_ON_N VSS 2.57201f 
C6522 a_22731_47423# VSS 0.227778f 
C6523 a_22223_47212# VSS 0.332189f 
C6524 a_12465_44636# VSS 5.61685f 
C6525 a_21811_47423# VSS 0.23358f 
C6526 a_4883_46098# VSS 1.54736f 
C6527 a_21496_47436# VSS 0.249536f 
C6528 a_13507_46334# VSS 4.83848f 
C6529 a_21177_47436# VSS 0.223524f 
C6530 a_20990_47178# VSS 0.224581f 
C6531 a_20894_47436# VSS 0.233111f 
C6532 a_19787_47423# VSS 0.258015f 
C6533 a_19386_47436# VSS 0.209882f 
C6534 a_18597_46090# VSS 2.82344f 
C6535 a_18780_47178# VSS 0.319719f 
C6536 a_18479_47436# VSS 1.19826f 
C6537 a_18143_47464# VSS 0.579061f 
C6538 a_10227_46804# VSS 8.12328f 
C6539 a_17591_47464# VSS 0.576556f 
C6540 a_16588_47582# VSS 0.263715f 
C6541 a_16763_47508# VSS 0.587861f 
C6542 a_16023_47582# VSS 0.264352f 
C6543 a_16327_47482# VSS 5.17799f 
C6544 a_16241_47178# VSS 0.18232f 
C6545 a_15673_47210# VSS 0.315684f 
C6546 a_15811_47375# VSS 0.349499f 
C6547 a_15507_47210# VSS 0.556554f 
C6548 a_11599_46634# VSS 2.84967f 
C6549 a_14955_47212# VSS 0.358339f 
C6550 a_14311_47204# VSS 0.248858f 
C6551 a_13487_47204# VSS 0.643275f 
C6552 a_12861_44030# VSS 3.64545f 
C6553 a_13717_47436# VSS 1.02478f 
C6554 a_n1435_47204# VSS 9.72476f 
C6555 a_13381_47204# VSS 0.225132f 
C6556 a_11459_47204# VSS 0.553679f 
C6557 a_9313_45822# VSS 1.04727f 
C6558 a_11031_47542# VSS 0.247302f 
C6559 a_9863_47436# VSS 0.265619f 
C6560 a_9067_47204# VSS 0.606182f 
C6561 a_6575_47204# VSS 0.798434f 
C6562 a_7903_47542# VSS 0.258657f 
C6563 a_7227_47204# VSS 0.610401f 
C6564 a_6851_47204# VSS 0.346433f 
C6565 a_6491_46660# VSS 0.343406f 
C6566 a_6545_47178# VSS 0.597936f 
C6567 a_6151_47436# VSS 2.12954f 
C6568 a_5815_47464# VSS 0.594449f 
C6569 a_5129_47502# VSS 0.361487f 
C6570 a_4915_47217# VSS 2.79467f 
C6571 a_n443_46116# VSS 4.167f 
C6572 a_4791_45118# VSS 2.65418f 
C6573 a_4700_47436# VSS 0.271201f 
C6574 a_4007_47204# VSS 0.628996f 
C6575 a_3815_47204# VSS 0.440491f 
C6576 a_3785_47178# VSS 0.541893f 
C6577 a_3381_47502# VSS 0.320926f 
C6578 a_n1151_42308# VSS 3.78206f 
C6579 a_3160_47472# VSS 0.607125f 
C6580 a_2905_45572# VSS 0.47073f 
C6581 a_2952_47436# VSS 0.275026f 
C6582 a_2553_47502# VSS 0.294118f 
C6583 a_2063_45854# VSS 1.92678f 
C6584 a_584_46384# VSS 2.10508f 
C6585 a_2124_47436# VSS 0.276508f 
C6586 a_1431_47204# VSS 0.595895f 
C6587 a_1239_47204# VSS 0.33333f 
C6588 a_1209_47178# VSS 0.474725f 
C6589 a_327_47204# VSS 0.581187f 
C6590 a_n785_47204# VSS 0.361759f 
C6591 a_n23_47502# VSS 0.278861f 
C6592 a_n237_47217# VSS 3.05697f 
C6593 a_n746_45260# VSS 0.993718f 
C6594 a_n971_45724# VSS 4.81311f 
C6595 a_n452_47436# VSS 0.28781f 
C6596 a_n815_47178# VSS 0.513835f 
C6597 a_n1605_47204# VSS 0.250546f 
C6598 SMPL_ON_P VSS 4.92073f 
C6599 a_n1741_47186# VSS 1.81488f 
C6600 a_n1920_47178# VSS 0.310881f 
C6601 a_n2109_47186# VSS 0.936844f 
C6602 a_n2288_47178# VSS 0.346995f 
C6603 a_n2497_47436# VSS 2.31207f 
C6604 a_n2833_47464# VSS 0.602779f 
C6605 w_11334_34010# VSS 50.9426f 
C6606 w_1575_34946# VSS 51.2247f 
.ends
