magic
tech sky130A
magscale 1 2
timestamp 1711813427
<< error_p >>
rect -29 272 29 278
rect 163 272 221 278
rect -29 238 -17 272
rect 163 238 175 272
rect -29 232 29 238
rect 163 232 221 238
<< pwell >>
rect 77 222 245 299
<< nmos >>
rect -111 -200 -81 200
rect -15 -200 15 200
rect 81 -200 111 200
<< ndiff >>
rect -173 188 -111 200
rect -173 -188 -161 188
rect -127 -188 -111 188
rect -173 -200 -111 -188
rect -81 188 -15 200
rect -81 -188 -65 188
rect -31 -188 -15 188
rect -81 -200 -15 -188
rect 15 188 81 200
rect 15 -188 31 188
rect 65 -188 81 188
rect 15 -200 81 -188
rect 111 188 173 200
rect 111 -188 127 188
rect 161 -188 173 188
rect 111 -200 173 -188
<< ndiffc >>
rect -161 -188 -127 188
rect -65 -188 -31 188
rect 31 -188 65 188
rect 127 -188 161 188
<< poly >>
rect -33 279 33 288
rect 159 279 225 288
rect -111 272 33 279
rect -111 238 -17 272
rect 17 238 33 272
rect -111 226 33 238
rect -111 200 -81 226
rect -33 222 33 226
rect 81 272 225 279
rect 81 238 175 272
rect 209 238 225 272
rect 81 226 225 238
rect -15 200 15 222
rect 81 200 111 226
rect 159 222 225 226
rect -111 -226 -81 -200
rect -15 -226 15 -200
rect 81 -226 111 -200
<< polycont >>
rect -17 238 17 272
rect 175 238 209 272
<< locali >>
rect -33 238 -17 272
rect 17 238 33 272
rect 159 238 175 272
rect 209 238 225 272
rect -161 188 -127 204
rect -161 -204 -127 -188
rect -65 188 -31 204
rect -65 -204 -31 -188
rect 31 188 65 204
rect 31 -204 65 -188
rect 127 188 161 204
rect 127 -204 161 -188
<< viali >>
rect -17 238 17 272
rect 175 238 209 272
rect -161 -188 -127 188
rect -65 -188 -31 188
rect 31 -188 65 188
rect 127 -188 161 188
<< metal1 >>
rect -29 272 29 278
rect -29 238 -17 272
rect 17 238 29 272
rect -29 232 29 238
rect 163 272 221 278
rect 163 238 175 272
rect 209 238 221 272
rect 163 232 221 238
rect -167 188 -121 200
rect -167 -188 -161 188
rect -127 -188 -121 188
rect -167 -200 -121 -188
rect -71 188 -25 200
rect -71 -188 -65 188
rect -31 -188 -25 188
rect -71 -200 -25 -188
rect 25 188 71 200
rect 25 -188 31 188
rect 65 -188 71 188
rect 25 -200 71 -188
rect 121 188 167 200
rect 121 -188 127 188
rect 161 -188 167 188
rect 121 -200 167 -188
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.150 m 1 nf 3 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
