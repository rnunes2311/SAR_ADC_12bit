* SPICE3 file created from SAR_ADC_12bit_flat.ext - technology: sky130A

.subckt SAR_ADC_12bit VDD VCM VSS VREF VIN_P VIN_N RST_Z CLK_DATA DATA[5] DATA[4] DATA[3] DATA[2] DATA[1] DATA[0] START EN_OFFSET_CAL CLK VREF_GND
+ SINGLE_ENDED
X0 a_13076_44458# a_13259_45724# a_13296_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2 VSS a_12427_45724# a_10490_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VDD a_2324_44458# a_949_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=361.2627 ps=3.22652k w=0.87 l=2.89
X5 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X6 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X7 VDD a_2903_42308# a_3080_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X8 VDD a_12861_44030# a_17829_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VSS a_1209_43370# a_n1557_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_16237_45028# a_16147_45260# a_16019_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X11 a_2075_43172# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VDD a_n755_45592# a_1176_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X13 a_6756_44260# a_5937_45572# a_6453_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X14 a_15868_43402# a_15681_43442# a_15781_43660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X15 a_n1533_42852# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X16 a_8103_44636# a_8375_44464# a_8333_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 VSS a_16327_47482# a_16377_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X18 a_2437_43646# a_n443_46116# a_2437_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_5088_37509# VSS VDAC_Ni VDD sky130_fd_pr__pfet_01v8_hvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X20 a_n2810_45028# a_n2840_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X21 a_2113_38308# VDAC_Ni a_2112_39137# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X22 VDD a_3626_43646# a_19647_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X23 VSS a_10334_44484# a_10440_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X24 a_1576_42282# a_1755_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X25 a_10933_46660# a_10554_47026# a_10861_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X26 a_14021_43940# a_13483_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X27 a_16867_43762# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X28 VREF a_21076_30879# C8_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X29 VSS a_n2946_37690# a_n3565_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 a_n913_45002# a_1307_43914# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 a_n2840_43370# a_n2661_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X32 a_3457_43396# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X33 a_14180_46482# a_14035_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X34 VSS a_18989_43940# a_19006_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X35 VSS a_9672_43914# a_2107_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X36 a_n1059_45260# a_17499_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X37 a_n1696_34930# a_n1794_35082# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X38 VSS a_10695_43548# a_10057_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X39 a_n2104_42282# a_n1925_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X40 a_20749_43396# a_12549_44172# a_743_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X41 VDD a_3877_44458# a_2382_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X42 a_n1699_44726# a_n1917_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X43 VSS a_n4334_39616# a_n4064_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X44 a_9241_45822# a_5066_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X45 VDD a_12883_44458# a_n2293_43922# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X46 a_11909_44484# a_3232_43370# a_11827_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X47 a_835_46155# a_584_46384# a_376_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X48 VSS a_1666_39043# a_1169_39043# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X49 a_5210_46155# a_5164_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X50 VDD a_n3690_39392# a_n3420_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X51 VDD a_167_45260# a_1609_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X52 VSS a_526_44458# a_3363_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X53 a_19268_43646# a_19319_43548# a_19095_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X54 VSS a_22959_44484# a_19237_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X55 a_n2216_39072# a_n2312_39304# a_n2302_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X56 a_19987_42826# a_10193_42453# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X57 a_6151_47436# a_14311_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X58 a_8145_46902# a_7927_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X59 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X60 a_14275_46494# a_13925_46122# a_14180_46482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X61 a_20512_43084# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X62 a_14539_43914# a_17701_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X63 a_6298_44484# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X64 a_644_44056# a_626_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X65 a_10949_43914# a_12429_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.28 ps=2.56 w=1 l=0.15
X66 VSS a_n2302_39866# a_n4209_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X67 VSS a_21811_47423# a_20916_46384# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X68 VDD a_3699_46634# a_3686_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X69 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X70 a_8035_47026# a_7411_46660# a_7927_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X71 a_5691_45260# a_5111_44636# a_5837_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X72 VDD a_1307_43914# a_1241_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X73 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X74 a_18249_42858# a_18083_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X75 VDD a_104_43370# a_n971_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X76 VDD a_n2833_47464# CLK_DATA VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X77 a_3363_44484# a_1823_45246# a_3232_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X78 a_n1331_43914# a_n1549_44318# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X79 VCM a_4958_30871# C9_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X80 VSS a_n3565_39590# a_n3607_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X81 VSS a_12281_43396# a_12563_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X82 VSS a_18780_47178# a_13661_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X83 a_n4318_39768# a_n2840_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X84 DATA[5] a_11459_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X85 a_7230_45938# a_6472_45840# a_6667_45809# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X86 VDD a_8049_45260# a_22959_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X87 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X88 a_8746_45002# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X89 a_15004_44636# a_11691_44458# a_15146_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X90 a_16223_45938# a_15599_45572# a_16115_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X91 a_n984_44318# a_n1899_43946# a_n1331_43914# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X92 a_n809_44244# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X93 a_n4064_39616# a_n4334_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X94 a_17124_42282# a_17303_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X95 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X96 VSS a_3065_45002# a_2680_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X97 a_5193_42852# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X98 VDD a_6969_46634# a_6999_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X99 VDD a_10623_46897# a_10554_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X100 a_16137_43396# a_15781_43660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X101 VDD a_n2472_46634# a_n2442_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X102 VDD a_4185_45028# a_22959_45036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X103 a_15225_45822# a_15037_45618# a_15143_45578# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X104 VSS a_3537_45260# a_4640_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X105 a_n2012_43396# a_n2129_43609# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X106 VDD a_n13_43084# a_n1853_43023# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X107 a_5068_46348# a_n1151_42308# a_5210_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X108 a_873_42968# a_685_42968# a_791_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X109 a_17730_32519# a_22591_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X110 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X111 VDD a_22485_44484# a_20974_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X112 a_n1021_46688# a_n1151_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X113 VSS a_11599_46634# a_11735_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X114 a_13163_45724# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.14075 ps=1.325 w=0.42 l=0.15
X115 C9_P_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X116 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X117 a_n2012_44484# a_n2129_44697# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X118 VIN_N EN_VIN_BSTR_N a_10890_34112# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X119 a_13940_44484# a_13556_45296# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X120 VSS a_1414_42308# a_1525_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X121 a_8487_44056# a_4223_44672# a_8415_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X122 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X123 a_16434_46660# a_16388_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X124 a_22613_38993# a_22527_39145# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X125 a_3315_47570# a_n1151_42308# a_2952_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X126 a_2680_45002# a_1823_45246# a_2903_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X127 a_1307_43914# a_2779_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X128 a_22731_47423# SMPL_ON_N VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X129 VDD a_1307_43914# a_3681_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X130 a_n863_45724# a_1667_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X131 VDD a_11459_47204# DATA[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X132 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X133 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X134 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=218.18214 ps=2.11206k w=0.55 l=0.59
X135 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X136 a_n4209_38216# a_n2302_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X137 a_10467_46802# a_11599_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X138 VDD a_13747_46662# a_19862_44208# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X139 a_n2946_39866# a_n2956_39768# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X140 a_n1013_45572# a_n1079_45724# a_n1099_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.182 ps=1.86 w=0.65 l=0.15
X141 VSS a_15279_43071# a_14579_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X142 DATA[3] a_7227_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X143 VSS a_8049_45260# a_22959_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X144 a_7584_44260# a_7542_44172# a_7281_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X145 a_n97_42460# a_19700_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X146 VDD a_19647_42308# a_13258_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X147 a_3754_39466# a_7754_39300# VSS sky130_fd_pr__res_high_po_0p35 l=18
X148 VSS a_2952_47436# a_2747_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X149 VDD a_16751_45260# a_6171_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X150 a_18326_43940# a_18079_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X151 a_9248_44260# a_8270_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X152 a_3503_45724# a_3775_45552# a_3733_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X153 a_n2017_45002# a_19987_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X154 a_288_46660# a_171_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X155 a_10037_46155# a_9804_47204# a_9823_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X156 a_20075_46420# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X157 VDD a_196_42282# a_n3674_37592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X158 VSS a_14513_46634# a_14447_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X159 a_n4064_39072# a_n4334_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X160 a_1149_42558# a_961_42354# a_1067_42314# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X161 a_13569_47204# a_13381_47204# a_13487_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X162 VDD a_14840_46494# a_15015_46420# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X163 C6_P_btm a_n3565_39304# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=0.35
X164 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X165 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X166 a_14537_43396# a_14358_43442# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X167 VDD a_14955_47212# a_10227_46804# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X168 VDD a_7754_40130# a_11206_38545# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X169 a_n3565_39590# a_n2946_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X170 a_n901_43156# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X171 a_17668_45572# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X172 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X173 a_15493_43396# a_14955_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X174 a_7309_43172# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X175 VDD a_1138_42852# a_1337_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X176 a_1427_43646# a_1568_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X177 a_18184_42460# a_15743_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X178 VDD a_13351_46090# a_10903_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X179 a_8379_46155# a_8128_46384# a_7920_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X180 VSS a_3483_46348# a_17325_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X181 VDD a_9290_44172# a_10949_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X182 VSS a_11823_42460# a_14358_43442# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X183 a_18310_42308# a_10193_42453# a_18220_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X184 VDD a_n2288_47178# a_n2312_40392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X185 a_17719_45144# a_16375_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X186 VDD a_5891_43370# a_5147_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X187 a_7287_43370# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X188 a_11173_44260# a_2063_45854# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X189 a_11897_42308# a_11823_42460# a_11551_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X190 VDD a_12861_44030# a_13759_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X191 a_19466_46812# a_19778_44110# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X192 a_9049_44484# a_8701_44490# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X193 a_n3565_38502# a_n2946_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X194 VDD a_16588_47582# a_16763_47508# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X195 a_9396_43370# a_4883_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X196 C0_P_btm a_n784_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X197 a_n1736_42282# a_n1557_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X198 VDD a_14113_42308# a_16522_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X199 a_10651_43940# a_3090_45724# a_10555_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.165 ps=1.33 w=1 l=0.15
X200 VDD a_8667_46634# a_n237_47217# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X201 a_6123_31319# a_7227_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X202 a_7499_43078# a_10083_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X203 VSS a_n755_45592# a_1145_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X204 C7_P_btm a_5534_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X205 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X206 VSS a_n4064_37984# a_n2302_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X207 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X208 a_3581_42558# a_3539_42460# a_3497_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X209 a_n3674_38680# a_n2840_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X210 VSS a_5907_45546# a_5937_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X211 VDD a_22589_40055# a_22527_39145# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X212 a_18783_43370# a_15743_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X213 VSS a_1799_45572# a_1983_46706# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X214 VDD a_22959_46660# a_21076_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X215 a_13467_32519# a_21487_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X216 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X217 a_2864_46660# a_2747_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X218 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X219 a_8199_44636# a_10355_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X220 a_14403_45348# a_13259_45724# a_14309_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X221 a_556_44484# a_742_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X222 VSS a_15433_44458# a_15367_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X223 a_n1794_35082# a_564_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X224 a_n2840_43370# a_n2661_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X225 w_1575_34786# a_n1696_34930# EN_VIN_BSTR_P w_1575_34786# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X226 VSS a_13747_46662# a_13693_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X227 a_18245_44484# a_17767_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X228 a_19741_43940# a_19862_44208# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X229 a_16855_43396# a_16409_43396# a_16759_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X230 a_13113_42826# a_12895_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X231 VSS a_22365_46825# a_20202_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X232 a_n1079_45724# a_n755_45592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X233 a_19386_47436# a_19321_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X234 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X235 VSS a_526_44458# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X236 a_n89_47570# a_n237_47217# a_n452_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X237 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X238 a_1176_45822# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X239 a_10341_43396# a_9803_43646# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X240 VDD a_n4209_38502# a_n4334_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X241 a_5111_42852# a_4905_42826# a_5193_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X242 a_13887_32519# a_22223_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X243 a_5437_45600# a_n881_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X244 a_18953_45572# a_18909_45814# a_18787_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X245 VDD a_4791_45118# a_6165_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X246 VDD a_3429_45260# a_3316_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.28 ps=2.56 w=1 l=0.15
X247 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X248 a_n3607_39616# a_n3674_39768# a_n3690_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X249 a_4842_47570# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X250 a_1337_46116# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X251 a_11136_45572# a_11322_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X252 a_n2661_42834# a_10809_44734# a_12189_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X253 VSS a_10249_46116# a_11186_47026# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X254 a_16655_46660# a_n743_46660# a_16292_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X255 a_n1991_46122# a_n2157_46122# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X256 VREF_GND a_n3420_39072# C6_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X257 a_n3565_37414# a_n2946_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X258 VDD a_1576_42282# a_1606_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X259 a_5159_47243# a_n443_46116# a_4700_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X260 VSS a_5891_43370# a_8375_44464# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X261 a_2075_43172# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X262 VDD a_13076_44458# a_12883_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X263 VSS a_14539_43914# a_14485_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X264 C0_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X265 a_15297_45822# a_11823_42460# a_15225_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X266 VSS a_18194_34908# a_10890_34112# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X267 VDD a_1169_39043# comp_n VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X268 a_18479_47436# a_20075_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X269 a_1423_45028# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X270 a_2382_45260# a_3877_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X271 a_8103_44636# a_8199_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X272 a_n1899_43946# a_n2065_43946# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X273 a_6765_43638# a_6547_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X274 VSS a_22400_42852# a_22848_40945# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X275 a_n2293_43922# a_12741_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X276 a_n3565_38216# a_n2946_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X277 VDD a_n3690_39392# a_n3420_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X278 a_945_42968# a_n1059_45260# a_873_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X279 VDD a_3785_47178# a_3815_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X280 VDD a_14084_46812# a_14035_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X281 a_765_45546# a_12549_44172# a_17829_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X282 VDD a_20974_43370# a_20556_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X283 a_14275_46494# a_13759_46122# a_14180_46482# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X284 VSS a_15051_42282# a_11823_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X285 a_1609_45822# a_n443_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X286 a_17517_44484# a_16979_44734# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X287 VDD a_4915_47217# a_12891_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X288 a_20679_44626# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X289 VSS a_1423_45028# a_9838_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X290 a_13921_42308# a_13259_45724# a_13575_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X291 VCM a_n784_42308# C0_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X292 VSS a_11599_46634# a_13759_46122# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X293 a_14127_45572# a_11823_42460# a_14033_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X294 VSS a_19998_34978# a_21753_35474# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X295 a_13569_43230# a_12379_42858# a_13460_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X296 a_5072_46660# a_4955_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X297 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X298 a_8037_42858# a_7871_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X299 VSS a_22591_46660# a_20820_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X300 VDD a_n2833_47464# CLK_DATA VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X301 a_3686_47026# a_2609_46660# a_3524_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X302 a_9672_43914# a_10057_43914# a_9801_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X303 VDD a_18429_43548# a_16823_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X304 a_17339_46660# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X305 VSS a_1606_42308# a_2351_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X306 a_16409_43396# a_16243_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X307 VSS a_9625_46129# a_10044_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X308 VDD a_n4209_37414# a_n4334_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X309 a_13468_44734# a_768_44030# a_13213_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X310 VSS a_n2302_39072# a_n4209_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X311 a_2124_47436# a_584_46384# a_2266_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X312 VDD a_n971_45724# a_2809_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X313 a_10809_44734# a_2063_45854# a_10809_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X314 a_7577_46660# a_7411_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X315 a_4921_42308# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X316 a_16023_47582# a_15507_47210# a_15928_47570# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X317 a_12791_45546# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X318 a_10193_42453# a_20712_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X319 VSS a_n881_46662# a_n659_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X320 a_6481_42558# a_n913_45002# a_1755_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X321 a_n2956_38680# a_n2472_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X322 a_14955_43940# a_14537_43396# a_15037_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X323 VREF_GND a_14097_32519# C4_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X324 VDD a_21188_45572# a_21363_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X325 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X326 a_15682_43940# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X327 a_18907_42674# a_18727_42674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X328 a_12545_42858# a_12379_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X329 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X330 C9_P_btm a_n4064_39616# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X331 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X332 a_13720_44458# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X333 a_15125_43396# a_15095_43370# a_15037_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X334 VREF a_20692_30879# C6_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=0.35
X335 a_2998_44172# a_584_46384# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X336 a_20974_43370# a_22485_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X337 a_18548_42308# a_18494_42460# a_18057_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X338 a_n875_44318# a_n2065_43946# a_n984_44318# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X339 a_n2293_42834# a_8049_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X340 VSS a_4743_44484# a_4791_45118# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X341 a_3626_43646# a_3232_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X342 VSS a_n2438_43548# a_n2433_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X343 a_n1076_43230# a_n2157_42858# a_n1423_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X344 VDD a_17973_43940# a_18079_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X345 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X346 VREF_GND a_17538_32519# C8_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X347 VDD a_22223_46124# a_20205_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X348 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X349 a_4704_46090# a_4883_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X350 a_5815_47464# a_6151_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X351 a_17478_45572# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X352 DATA[3] a_7227_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X353 VDD a_n1794_35082# a_18194_34908# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X354 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X355 a_17034_45572# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X356 VSS a_n3420_39616# a_n2946_39866# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X357 a_133_42852# a_n97_42460# a_n13_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X358 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X359 a_n1925_46634# a_8162_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X360 a_21350_47026# a_20273_46660# a_21188_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X361 VDD a_2713_42308# a_2903_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X362 a_n3674_39304# a_n2840_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X363 a_13565_43940# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X364 a_n4315_30879# a_n2302_40160# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X365 VDD a_1823_45246# a_2202_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X366 VSS a_n3690_38304# a_n3420_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X367 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X368 a_2211_45572# a_2063_45854# a_1848_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X369 VSS a_16112_44458# a_14673_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X370 VSS a_3316_45546# a_3260_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X371 VDD a_n443_46116# a_2896_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X372 a_n310_47570# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X373 a_21177_47436# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X374 VSS a_9290_44172# a_13943_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X375 a_n3674_37592# a_196_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X376 a_18780_47178# a_18597_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X377 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X378 VSS a_8791_42308# a_5934_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X379 a_421_43172# a_n97_42460# a_n13_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X380 VDD a_17339_46660# a_18051_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X381 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X382 VSS a_n2840_46090# a_n2956_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X383 a_n2661_43370# a_10907_45822# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X384 a_9396_43370# a_4883_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X385 VDD a_19333_46634# a_19123_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X386 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X387 a_5755_42852# a_n97_42460# a_5837_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X388 a_n4251_39392# a_n4318_39304# a_n4334_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X389 a_805_46414# a_472_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X390 VDD a_n1076_43230# a_n901_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X391 a_21845_43940# a_12549_44172# a_19692_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X392 VDD a_4520_42826# a_4093_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X393 a_12469_46902# a_12251_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X394 a_15415_45028# a_15227_44166# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X395 a_19479_31679# a_22223_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X396 a_7542_44172# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X397 a_3080_42308# a_2903_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X398 VSS a_22165_42308# a_22223_42860# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X399 VDD a_10249_46116# a_11186_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X400 a_3905_42558# a_2382_45260# a_3823_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X401 a_12347_46660# a_11901_46660# a_12251_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X402 VSS a_16137_43396# a_16414_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.089375 ps=0.925 w=0.65 l=0.15
X403 a_5066_45546# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X404 a_14581_44484# a_13249_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X405 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X406 a_2113_38308# a_1273_38525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X407 a_n473_42460# a_n755_45592# a_n327_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X408 VDD a_n1699_43638# a_n1809_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X409 a_13759_47204# a_13717_47436# a_13675_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X410 a_n3420_39616# a_n3690_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X411 C4_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X412 a_n967_46494# a_n2157_46122# a_n1076_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X413 a_2779_44458# a_1423_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X414 VDD a_19319_43548# a_19268_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.195 ps=1.39 w=1 l=0.15
X415 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X416 VDD a_9127_43156# a_5891_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X417 a_1123_46634# a_948_46660# a_1302_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X418 a_n755_45592# a_n809_44244# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X419 a_2952_47436# a_3160_47472# a_3094_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X420 a_5807_45002# a_16763_47508# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X421 a_3726_37500# a_3754_38470# VDAC_Ni VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X422 a_6293_42852# a_5755_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X423 a_8120_45572# a_8034_45724# a_n1925_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X424 a_11541_44484# a_11691_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X425 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X426 VSS a_10083_42826# a_7499_43078# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X427 a_5257_43370# a_5907_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X428 a_4880_45572# a_5066_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X429 VIN_P EN_VIN_BSTR_P C0_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X430 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X431 a_3497_42558# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X432 VSS a_1123_46634# a_584_46384# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X433 a_16223_45938# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X434 a_4883_46098# a_21363_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X435 a_2711_45572# a_768_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X436 VSS a_2553_47502# a_2487_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X437 VDD a_12469_46902# a_12359_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X438 a_6453_43914# a_6109_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X439 a_7765_42852# a_7227_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X440 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X441 a_17786_45822# a_15861_45028# a_17478_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X442 a_18450_45144# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X443 a_6765_43638# a_6547_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X444 a_n914_46116# a_n1991_46122# a_n1076_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X445 VSS a_n4334_40480# a_n4064_40160# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X446 a_12089_42308# a_11551_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X447 a_16547_43609# a_16414_43172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X448 a_3221_46660# a_3177_46902# a_3055_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X449 a_6667_45809# a_6472_45840# a_6977_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X450 a_n1190_43762# a_n2267_43396# a_n1352_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X451 a_6643_43396# a_6197_43396# a_6547_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X452 a_5837_45348# a_5807_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X453 a_5565_43396# a_4905_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X454 a_7418_45067# a_7229_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X455 a_1307_43914# a_2779_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X456 a_1793_42852# a_742_44458# a_1709_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X457 VDD a_10227_46804# a_10083_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X458 a_11301_43218# a_10922_42852# a_11229_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X459 VSS a_13291_42460# a_13249_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X460 a_18341_45572# a_18175_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X461 w_1575_34786# a_n1057_35014# w_1575_34786# w_1575_34786# sky130_fd_pr__pfet_01v8 ad=0.986 pd=7.38 as=10.006 ps=72.76 w=3.4 l=16.6
X462 a_19113_45348# a_19321_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X463 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X464 a_8696_44636# a_16855_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X465 a_12189_44484# a_8975_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X466 a_n1736_46482# a_n1853_46287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X467 a_1239_47204# a_1209_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X468 VSS a_n1696_34930# a_n217_35014# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X469 VDD VDAC_Ni a_6886_37412# VSS sky130_fd_pr__nfet_03v3_nvt ad=0.0725 pd=0.79 as=0.145 ps=1.58 w=0.5 l=0.5
X470 a_n4064_37984# a_n4334_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X471 a_1606_42308# a_1576_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X472 VDD a_n443_42852# a_6481_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X473 VDD a_12005_46116# a_n1741_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X474 a_18315_45260# a_18587_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X475 VSS a_768_44030# a_3600_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X476 VDD a_4958_30871# a_17531_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X477 a_16795_42852# a_n97_42460# a_16877_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X478 a_18900_46660# a_18834_46812# a_18285_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X479 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X480 a_17973_43940# a_17737_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X481 a_6419_46155# a_5257_43370# a_6347_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X482 a_18597_46090# a_19431_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X483 a_3737_43940# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X484 comp_n a_1169_39043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X485 VDD a_1823_45246# a_4419_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X486 a_22848_40945# COMP_P a_22589_40599# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X487 VDD a_4007_47204# DATA[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X488 VSS a_21496_47436# a_13507_46334# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X489 VDD a_n2002_35448# SMPL_ON_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X490 VSS a_10723_42308# a_5742_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X491 a_22737_36887# a_22527_39145# a_22629_37990# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X492 a_11823_42460# a_15051_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X493 VSS a_n4209_38216# a_n4251_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X494 a_12891_46348# a_4915_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X495 VSS a_20679_44626# a_20640_44752# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X496 a_21115_43940# a_20935_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X497 a_n1821_43396# a_n2267_43396# a_n1917_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X498 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X499 VDD a_10951_45334# a_10775_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X500 a_20850_46155# a_19692_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X501 VDD a_13661_43548# a_18587_45118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X502 a_11649_44734# a_3232_43370# a_n2661_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.174 ps=1.39 w=1 l=0.15
X503 a_20820_30879# a_22591_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X504 VSS a_21359_45002# a_21101_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X505 EN_VIN_BSTR_N a_18194_34908# w_10694_33990# w_10694_33990# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X506 a_17364_32525# a_22959_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X507 a_18989_43940# a_18451_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X508 a_6197_43396# a_6031_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X509 VDD a_12891_46348# a_13213_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X510 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X511 VREF_GND a_13467_32519# C1_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X512 VDD a_584_46384# a_3540_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.175 ps=1.35 w=1 l=0.15
X513 a_8873_43396# a_5891_43370# a_8791_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X514 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X515 VSS a_n4334_39392# a_n4064_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X516 C9_P_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X517 a_10809_44484# a_10057_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X518 C6_N_btm a_5742_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X519 a_6545_47178# a_6419_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X520 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X521 a_6109_44484# a_5518_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X522 a_n4318_38216# a_n2472_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X523 VDD a_n901_46420# a_n443_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X524 a_13258_32519# a_19647_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X525 VDD a_11599_46634# a_18819_46122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X526 a_18194_34908# a_n1794_35082# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X527 a_n1435_47204# a_n1605_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X528 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X529 a_15682_43940# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X530 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X531 a_14113_42308# a_13575_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X532 VSS a_4646_46812# a_4651_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X533 a_13381_47204# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X534 VSS a_n2472_46090# a_n2956_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X535 a_4958_30871# a_17124_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X536 VSS a_22223_42860# a_22400_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X537 C0_P_btm a_n3565_37414# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X538 VDD a_1208_46090# a_472_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X539 VSS a_18479_47436# a_19452_47524# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X540 VSS a_n2302_39072# a_n4209_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X541 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X542 a_n443_46116# a_n901_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X543 a_20623_45572# a_20107_45572# a_20528_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X544 a_12281_43396# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X545 VSS a_n1794_35082# a_18194_34908# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X546 C1_P_btm a_n4209_37414# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X547 VSS a_n3565_39304# a_n3607_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X548 a_15486_42560# a_15764_42576# a_15720_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X549 VSS a_n1613_43370# a_8649_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X550 a_15765_45572# a_15599_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X551 VSS a_n2946_39866# a_n3565_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X552 a_n1613_43370# a_5815_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X553 VSS a_14495_45572# a_n881_46662# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X554 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X555 a_10617_44484# a_10440_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X556 VDD a_5111_44636# a_8487_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X557 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X558 VCM a_5932_42308# C3_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X559 a_20708_46348# a_15227_44166# a_20850_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X560 a_n2267_44484# a_n2433_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X561 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X562 a_1115_44172# a_453_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X563 VSS COMP_P a_n1329_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X564 VSS a_1847_42826# a_2905_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X565 VSS a_15861_45028# a_17023_45118# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X566 a_16292_46812# a_5807_45002# a_16434_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X567 a_17325_44484# a_15227_44166# a_16979_44734# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X568 a_n4064_39072# a_n4334_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X569 a_15803_42450# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X570 a_5534_30871# a_12563_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X571 VSS a_3381_47502# a_3315_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X572 VDD a_9863_46634# a_2063_45854# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X573 VDD a_n2840_43370# a_n4318_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X574 VSS a_584_46384# a_3457_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X575 VIN_N EN_VIN_BSTR_N C3_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X576 a_3863_42891# a_3681_42891# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X577 VDD a_9049_44484# a_9313_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X578 VDD a_376_46348# a_171_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X579 a_11541_44484# a_11453_44696# a_n2661_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X580 VDD a_1431_47204# DATA[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X581 a_19553_46090# a_19335_46494# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X582 a_n1613_43370# a_5815_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X583 a_18727_42674# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X584 a_n1925_42282# a_4185_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X585 VDD a_n2302_37984# a_n4209_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X586 VSS a_17591_47464# a_16327_47482# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X587 VSS a_n3690_38304# a_n3420_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X588 VDD a_19164_43230# a_19339_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X589 a_2479_44172# a_2905_42968# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X590 VSS a_4361_42308# a_21855_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X591 a_n1741_47186# a_12891_46348# a_12839_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X592 VDD a_8103_44636# a_7640_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X593 a_8192_45572# a_8162_45546# a_8120_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X594 a_5009_45028# a_3090_45724# a_4927_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X595 a_12549_44172# a_20567_45036# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X596 VSS a_n2840_42282# a_n3674_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X597 a_5129_47502# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X598 a_14840_46494# a_13759_46122# a_14493_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X599 VSS a_2324_44458# a_949_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X600 VDD EN_VIN_BSTR_N w_10694_33990# w_10694_33990# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X601 VSS a_n913_45002# a_2713_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X602 VDD a_n863_45724# a_1221_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X603 a_8601_46660# a_7411_46660# a_8492_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X604 a_2307_45899# a_n237_47217# a_1848_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X605 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X606 VDD a_n4209_39304# a_n4334_39392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X607 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X608 a_n2946_39072# a_n2956_39304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X609 a_15861_45028# a_15595_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X610 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X611 VSS a_n1613_43370# a_3221_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X612 a_1756_43548# a_768_44030# a_1987_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X613 a_3754_39134# a_7754_39300# VSS sky130_fd_pr__res_high_po_0p35 l=18
X614 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X615 a_n4318_40392# a_n2840_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X616 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X617 VSS a_18143_47464# a_12861_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X618 a_19332_42282# a_19511_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X619 VSS a_17583_46090# a_13259_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X620 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X621 a_20623_43914# a_19321_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X622 VSS a_17499_43370# a_n1059_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X623 VSS a_7754_38470# a_6886_37412# VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X624 a_n3420_39616# a_n3690_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X625 a_4185_45348# a_3065_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X626 a_n2661_46634# a_13017_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X627 VDD a_19321_45002# a_20567_45036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X628 VDD a_6545_47178# a_6575_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X629 VDD a_18285_46348# a_18051_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.16 ps=1.32 w=1 l=0.15
X630 a_2864_46660# a_2747_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X631 VSS a_n809_44244# a_n755_45592# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X632 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X633 VDD a_1307_43914# a_2253_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X634 a_n2002_35448# a_n1550_35448# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X635 a_13351_46090# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X636 a_18374_44850# a_18248_44752# a_17970_44736# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X637 a_n913_45002# a_1307_43914# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X638 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X639 a_13657_42308# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X640 a_375_42282# a_413_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X641 a_3090_45724# a_19321_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=1.67 w=1 l=0.15
X642 a_n1696_34930# a_n1794_35082# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X643 a_10334_44484# a_10157_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X644 VSS a_10903_43370# a_10057_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X645 a_5700_37509# VSS VDAC_Pi VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X646 a_2113_38308# a_2113_38308# a_2113_38308# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=3.02 ps=24.88 w=1 l=0.15
X647 VSS a_n2438_43548# a_n133_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X648 a_584_46384# a_1123_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X649 VSS a_22959_46124# a_20692_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X650 a_n3674_39768# a_n2472_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X651 VREF a_n4209_39304# C7_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X652 VSS a_20107_42308# a_7174_31319# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X653 a_n4209_39590# a_n2302_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X654 a_526_44458# a_3147_46376# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X655 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X656 a_20301_43646# a_19692_46634# a_20556_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X657 VDD a_n901_46420# a_n914_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X658 a_n971_45724# a_104_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X659 a_20447_31679# a_22959_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X660 VSS a_13348_45260# a_13159_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X661 a_n4334_38304# a_n4318_38216# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X662 VSS a_n881_46662# a_6517_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X663 a_8685_42308# a_8515_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X664 VSS a_6491_46660# a_6851_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X665 a_768_44030# a_13487_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X666 VDD a_14493_46090# a_14383_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X667 a_n327_42308# a_n357_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X668 a_22485_44484# a_22315_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X669 a_15673_47210# a_15507_47210# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X670 a_8605_42826# a_8387_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X671 a_1709_42852# a_n863_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X672 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X673 VDD a_n1736_42282# a_n4318_37592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X674 VREF a_19721_31679# C2_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X675 VSS a_895_43940# a_2537_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X676 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X677 a_17609_46634# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X678 VDD a_11599_46634# a_18175_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X679 a_8945_43396# a_3537_45260# a_8873_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X680 a_13249_42308# a_10903_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X681 a_601_46902# a_383_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X682 a_4640_45348# a_4574_45260# a_4558_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X683 a_n467_45028# a_n745_45366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X684 a_1208_46090# a_765_45546# a_1337_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X685 a_3820_44260# a_2382_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X686 VSS a_n863_45724# a_2905_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X687 VSS a_16721_46634# a_16655_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X688 C5_P_btm a_n4064_38528# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X689 a_21588_30879# a_22223_47212# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X690 a_16877_42852# a_16823_43084# a_16795_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X691 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X692 VSS a_17715_44484# a_17737_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X693 a_16241_47178# a_16023_47582# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X694 a_12359_47026# a_11735_46660# a_12251_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X695 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X696 a_5883_43914# a_8333_44056# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X697 a_16759_43396# a_16409_43396# a_16664_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X698 VDD a_n3565_39590# a_n3690_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X699 a_17665_42852# a_17595_43084# a_14539_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X700 VSS a_n2438_43548# a_n2157_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X701 VDD a_4007_47204# DATA[2] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X702 a_1990_45572# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X703 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X704 a_5072_46660# a_4955_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X705 a_22889_38993# a_22400_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X706 VDD a_3357_43084# a_22591_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X707 VSS a_3815_47204# a_4007_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X708 a_1666_39587# a_1666_39043# a_2112_39137# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X709 a_15803_42450# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X710 a_20528_46660# a_20411_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X711 a_n3607_39392# a_n3674_39304# a_n3690_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X712 VDD a_n4064_39616# a_n2216_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X713 a_21421_42336# a_16327_47482# a_21335_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X714 a_6655_43762# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X715 a_14371_46494# a_13925_46122# a_14275_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X716 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X717 VDD a_3503_45724# a_3218_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X718 VDD a_n2840_43914# a_n4318_39768# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X719 a_15037_43940# a_13556_45296# a_14955_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X720 VSS a_n901_43156# a_n443_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X721 VDD a_10467_46802# a_10428_46928# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X722 a_15060_45348# a_13661_43548# a_14976_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X723 a_9895_44260# a_9290_44172# a_9801_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X724 VDD a_6171_42473# a_5379_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X725 a_5009_45028# a_5147_45002# a_5093_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X726 a_13904_45546# a_10903_43370# a_14127_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X727 a_3537_45260# a_7287_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X728 SMPL_ON_N a_21753_35474# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X729 a_19900_46494# a_18985_46122# a_19553_46090# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X730 VDD a_8696_44636# a_17478_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X731 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X732 a_3935_42891# a_3905_42865# a_3863_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X733 DATA[0] a_327_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X734 VSS a_n881_46662# a_11117_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X735 C3_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X736 VSS a_n4334_39616# a_n4064_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X737 DATA[2] a_4007_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X738 a_15682_46116# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X739 a_1057_46660# a_n133_46660# a_948_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X740 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X741 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X742 VSS a_2982_43646# a_21487_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X743 a_21363_45546# a_21188_45572# a_21542_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X744 VSS a_11823_42460# a_11322_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X745 a_18204_44850# a_17767_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X746 a_n447_43370# a_n2497_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X747 a_17324_43396# a_16409_43396# a_16977_43638# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X748 VSS a_n4064_38528# a_n2302_38778# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X749 a_n443_42852# a_n901_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X750 a_15095_43370# a_15567_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X751 a_10150_46912# a_10428_46928# a_10384_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X752 VSS a_n2472_42282# a_n4318_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X753 VDD a_21753_35474# SMPL_ON_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X754 a_8492_46660# a_7577_46660# a_8145_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X755 a_5649_42852# a_5111_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X756 VDD a_18287_44626# a_18248_44752# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X757 a_20894_47436# a_20990_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X758 a_19636_46660# a_19594_46812# a_19333_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X759 a_10249_46116# a_9823_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X760 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X761 a_10227_46804# a_14955_47212# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X762 a_739_46482# a_n743_46660# a_376_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X763 VSS a_10775_45002# a_10180_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X764 a_2896_43646# a_2479_44172# a_2982_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X765 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X766 a_12791_45546# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X767 VSS a_5807_45002# a_11691_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X768 VSS a_3357_43084# a_22591_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X769 VSS a_2382_45260# a_2304_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X770 a_n4315_30879# a_n2302_40160# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X771 VDD a_n901_46420# a_n443_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X772 a_6298_44484# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X773 a_949_44458# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X774 VDD a_2277_45546# a_2307_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X775 a_10053_45546# a_8746_45002# a_10306_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X776 a_18194_34908# a_n1794_35082# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X777 a_n2956_39768# a_n2840_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X778 VDD a_4361_42308# a_21855_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X779 VDD a_17591_47464# a_16327_47482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X780 VSS a_6945_45028# a_22223_46124# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X781 VDD a_5257_43370# a_5263_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X782 a_n3565_39590# a_n2946_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X783 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X784 VDAC_Ni VSS a_5088_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X785 a_18494_42460# a_18907_42674# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X786 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X787 a_n1151_42308# a_n1329_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X788 a_16763_47508# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X789 a_21259_43561# a_4190_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X790 a_8349_46414# a_8016_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X791 VDD a_1431_47204# DATA[1] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X792 a_17970_44736# a_18287_44626# a_18245_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X793 a_1123_46634# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X794 a_n237_47217# a_8667_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3012 ps=2.66 w=1 l=0.15
X795 a_5837_42852# a_3537_45260# a_5755_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X796 VSS a_19692_46634# a_19636_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X797 a_8697_45572# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X798 a_1145_45348# a_n863_45724# a_626_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X799 VSS a_5934_30871# a_8515_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X800 VSS a_1239_47204# a_1431_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X801 VSS a_17591_47464# a_16327_47482# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X802 a_11173_44260# a_10729_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X803 VDD a_n4334_38304# a_n4064_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X804 a_22165_42308# a_21887_42336# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X805 a_5244_44056# a_5147_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X806 VSS a_n4064_37440# a_n2302_37690# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X807 VDD a_8952_43230# a_9127_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X808 a_n2956_37592# a_n2472_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X809 VSS a_2127_44172# a_n2661_45010# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X810 VSS a_15493_43940# a_22959_43948# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X811 a_n3565_38502# a_n2946_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X812 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X813 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X814 a_19339_43156# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X815 VDD a_n1920_47178# a_n2312_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X816 VDD a_n1177_44458# a_n1190_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X817 VDD a_16292_46812# a_15811_47375# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X818 a_5164_46348# a_4927_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X819 a_9482_43914# a_9838_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X820 a_20835_44721# a_20679_44626# a_20980_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X821 VSS a_5937_45572# a_8781_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X822 a_5837_42852# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X823 a_10037_47542# a_n881_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X824 a_7221_43396# a_6031_43396# a_7112_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X825 VSS a_5937_45572# a_8560_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X826 C7_N_btm a_20820_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X827 VSS a_15559_46634# a_13059_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X828 a_5385_46902# a_5167_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X829 VDD a_10334_44484# a_10440_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X830 a_19597_46482# a_19553_46090# a_19431_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X831 VDD a_n2302_37984# a_n4209_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X832 a_18051_46116# a_18189_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.165 ps=1.33 w=1 l=0.15
X833 a_15493_43940# a_14955_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X834 a_19250_34978# VDD EN_VIN_BSTR_N VSS sky130_fd_pr__nfet_05v0_nvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.9
X835 a_16414_43172# a_n1059_45260# a_16328_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X836 a_21297_46660# a_20107_46660# a_21188_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X837 a_11813_46116# a_11387_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X838 VSS a_1666_39587# a_1169_39587# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X839 VSS SMPL_ON_P a_n1605_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X840 DATA[4] a_9067_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X841 a_5894_47026# a_4817_46660# a_5732_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X842 VDD a_4699_43561# a_3539_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X843 VSS a_n3420_39072# a_n2946_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X844 VDD a_n97_42460# a_16245_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X845 VDD a_13163_45724# a_11962_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X846 a_15433_44458# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X847 VDD a_16327_47482# a_20980_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X848 a_18114_32519# a_22223_45036# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X849 a_n452_44636# a_n1151_42308# a_n310_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X850 VDD a_22959_43396# a_17364_32525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X851 a_n4064_37984# a_n4334_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X852 VDD a_1307_43914# a_4149_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X853 VSS a_n357_42282# a_7573_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X854 VDD a_9863_47436# a_9804_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X855 a_3754_39134# a_7754_38968# VSS sky130_fd_pr__res_high_po_0p35 l=18
X856 a_4649_43172# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X857 a_526_44458# a_3147_46376# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X858 VSS a_1848_45724# a_1799_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X859 a_22485_38105# a_22775_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X860 a_20885_45572# a_20841_45814# a_20719_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X861 a_10554_47026# a_10428_46928# a_10150_46912# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X862 a_n746_45260# a_n1177_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X863 a_7_44811# a_n1151_42308# a_n452_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X864 VDD a_2324_44458# a_15682_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X865 VDD a_10355_46116# a_8199_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X866 a_4181_43396# a_4093_43548# a_n2661_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X867 VDD a_2437_43646# a_22223_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X868 a_21005_45260# a_21101_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X869 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X870 a_n3565_37414# a_n2946_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X871 a_3754_38802# a_7754_38968# VSS sky130_fd_pr__res_high_po_0p35 l=18
X872 a_2075_43172# a_1307_43914# a_n913_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X873 VSS a_17499_43370# a_n1059_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X874 VSS a_12861_44030# a_17339_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X875 VDD a_n2840_45002# a_n2810_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X876 a_10057_43914# a_10807_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X877 a_5343_44458# a_7963_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X878 a_n1423_42826# a_n1641_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X879 a_526_44458# a_3147_46376# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X880 VDD a_11827_44484# a_22223_45036# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X881 VDD a_n2472_43914# a_n3674_39768# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X882 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X883 a_6945_45028# a_5937_45572# a_6945_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X884 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X885 a_20301_43646# a_13661_43548# a_743_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X886 VDD a_n3690_39616# a_n3420_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X887 a_n2216_39866# a_n2442_46660# a_n2302_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X888 VDD a_22000_46634# a_15227_44166# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X889 VSS a_2889_44172# a_413_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X890 VSS a_n97_42460# a_n144_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X891 a_n3674_38216# a_n2104_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X892 a_16321_45348# a_1307_43914# a_16019_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.183625 ps=1.215 w=0.65 l=0.15
X893 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X894 VDD a_9290_44172# a_13070_42354# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X895 a_133_42852# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X896 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X897 a_n3420_39072# a_n3690_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X898 a_n2860_38778# a_n2956_38680# a_n2946_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X899 a_22485_38105# a_22775_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X900 a_6517_45366# a_5937_45572# a_6431_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X901 a_10555_44260# a_10729_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X902 VDD a_5111_44636# a_5837_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X903 a_14401_32519# a_22223_43948# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X904 VSS a_9290_44172# a_13070_42354# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X905 VSS a_5068_46348# a_4955_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X906 VDD a_9290_44172# a_10586_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X907 a_16751_45260# a_8696_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X908 a_1666_39587# a_1666_39043# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X909 a_n913_45002# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X910 VSS a_11599_46634# a_15507_47210# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X911 VSS a_768_44030# a_644_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X912 a_12465_44636# a_5807_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X913 VDD a_n357_42282# a_16877_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X914 a_5193_43172# a_3905_42865# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X915 VSS a_18783_43370# a_18525_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X916 a_3540_43646# a_1414_42308# a_3626_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.14 ps=1.28 w=1 l=0.15
X917 a_21363_45546# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X918 VSS a_n3690_38528# a_n3420_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X919 a_5421_42558# a_5379_42460# a_5337_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X920 VDD a_12861_44030# a_17609_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X921 a_n2956_38216# a_n2472_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X922 a_13885_46660# a_13607_46688# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X923 VCM a_4958_30871# C9_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X924 a_2232_45348# a_1609_45822# a_n2293_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X925 a_5691_45260# a_6171_45002# a_5837_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X926 a_9801_44260# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X927 VCM a_3080_42308# C2_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X928 a_327_44734# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X929 VSS a_7499_43078# a_8746_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X930 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X931 a_15743_43084# a_19339_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X932 VSS a_22591_43396# a_14209_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X933 VSS a_2437_43646# a_22223_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X934 a_6547_43396# a_6197_43396# a_6452_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X935 a_20556_43646# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X936 a_1987_43646# a_742_44458# a_1891_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X937 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X938 a_648_43396# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X939 VDD a_n23_47502# a_7_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X940 a_17609_46634# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X941 a_3602_45348# a_3537_45260# a_3495_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X942 VDD CLK a_8953_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X943 VDD a_2982_43646# a_21487_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X944 a_13661_43548# a_18780_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X945 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X946 a_9313_44734# a_3232_43370# a_9159_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X947 C6_P_btm a_5742_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X948 a_11323_42473# a_5742_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X949 a_14383_46116# a_13759_46122# a_14275_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X950 a_2813_43396# a_2479_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X951 a_16721_46634# a_16388_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X952 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X953 VDD a_526_44458# a_9885_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X954 VSS a_22537_40625# a_22737_36887# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X955 VREF a_20820_30879# C7_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X956 VDD a_15681_43442# a_15781_43660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X957 a_6125_45348# a_3232_43370# a_5691_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X958 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X959 a_10907_45822# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X960 a_14955_43396# a_9145_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X961 a_8128_46384# a_7903_47542# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X962 a_3429_45260# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X963 VDD a_15227_44166# a_17969_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06405 ps=0.725 w=0.42 l=0.15
X964 DATA[0] a_327_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X965 a_n2860_37690# a_n2956_37592# a_n2946_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X966 a_15682_46116# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X967 VSS a_7287_43370# a_3537_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X968 C4_P_btm a_n3420_38528# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X969 a_18599_43230# a_18083_42858# a_18504_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X970 DATA[2] a_4007_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X971 a_18057_42282# a_18494_42460# a_18214_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X972 a_11117_47542# a_4915_47217# a_11031_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X973 w_10694_33990# a_18194_34908# EN_VIN_BSTR_N w_10694_33990# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X974 a_7112_43396# a_6197_43396# a_6765_43638# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X975 a_584_46384# a_1123_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X976 VSS a_n3690_37440# a_n3420_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X977 VSS a_n901_43156# a_n443_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X978 a_19240_46482# a_19123_46287# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X979 VCM a_5742_30871# C6_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X980 VSS a_10193_42453# a_10149_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X981 VDD a_10193_42453# a_10210_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X982 VSS a_2324_44458# a_15682_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X983 EN_VIN_BSTR_N VDD a_19250_34978# VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.9
X984 VSS a_n967_45348# a_n961_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X985 a_564_42282# a_743_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X986 a_21195_42852# a_20922_43172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X987 VDD a_6575_47204# a_9067_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X988 a_22612_30879# a_22959_47212# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X989 a_21188_46660# a_20273_46660# a_20841_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X990 a_13749_43396# a_13661_43548# a_13667_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X991 VSS a_n2840_45546# a_n2810_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X992 a_13490_45394# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X993 a_n2840_43914# a_n2661_43922# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X994 a_n822_43940# a_n1899_43946# a_n984_44318# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X995 a_21613_42308# a_21335_42336# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X996 a_7112_43396# a_6031_43396# a_6765_43638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X997 a_14537_43396# a_13059_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X998 VDAC_Pi a_3754_38470# a_4338_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X999 a_n4064_39616# a_n4334_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1000 a_n23_47502# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X1001 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1002 a_14543_43071# a_5534_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1003 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1004 VDD a_19900_46494# a_20075_46420# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1005 VDD a_7227_45028# a_7230_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1006 VSS a_16327_47482# a_19597_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1007 a_9823_46155# a_n743_46660# a_9751_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1008 VDD a_22959_43948# a_17538_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1009 a_18214_42558# a_16137_43396# a_18057_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1010 a_n3690_38304# a_n3674_38216# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1011 a_15009_46634# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1012 a_17591_47464# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X1013 VSS a_10227_46804# a_15521_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1014 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1015 a_22485_44484# a_22315_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1016 a_n1644_44306# a_n1761_44111# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1017 VDD RST_Z a_8530_39574# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1018 VDD a_n1329_42308# a_n1151_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1019 VSS a_13507_46334# a_18184_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1020 a_n630_44306# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1021 a_18783_43370# a_15743_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1022 a_n4064_38528# a_n4334_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1023 a_8325_42308# a_n913_45002# a_8337_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1024 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X1025 a_21973_42336# a_20202_43084# a_21887_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1026 VSS a_n1613_43370# a_645_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1027 a_10341_42308# a_9803_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1028 a_n1920_47178# a_n1741_47186# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1029 VSS a_16327_47482# a_20885_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1030 VSS a_10807_43548# a_11173_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1031 VSS a_5257_43370# a_3905_42865# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1032 a_9127_43156# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1033 VDD a_n2472_45002# a_n2956_37592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1034 VSS a_n2946_39072# a_n3565_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1035 a_13259_45724# a_17583_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1036 VSS a_10586_45546# a_10544_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X1037 a_16751_45260# a_17023_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1038 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1039 VSS a_n4209_38502# a_n4251_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X1040 VSS a_7227_42308# a_6123_31319# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1041 VSS a_10083_42826# a_7499_43078# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1042 a_n2840_42826# a_n2661_42834# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1043 a_1302_46660# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1044 a_5907_45546# a_6194_45824# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1045 a_13059_46348# a_15559_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1046 a_n2302_37984# a_n2810_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1047 VREF_GND a_14209_32519# C5_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1048 a_3065_45002# a_3318_42354# a_3581_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X1049 a_16023_47582# a_15673_47210# a_15928_47570# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1050 VSS a_n881_46662# a_n935_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1051 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1052 C6_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1053 VDD a_21487_43396# a_13467_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1054 a_2553_47502# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X1055 VDD a_n443_42852# a_997_45618# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X1056 a_8568_45546# a_8199_44636# a_8791_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1057 a_4338_37500# a_3754_38470# VDAC_Pi VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1058 a_13635_43156# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1059 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1060 VDD a_564_42282# a_n1794_35082# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1061 a_n473_42460# a_n971_45724# a_n327_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X1062 a_16335_44484# a_13661_43548# a_16241_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X1063 VDD a_15861_45028# a_17023_45118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1064 a_5205_44734# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1065 a_7499_43078# a_10083_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=2.61 w=1 l=0.15
X1066 VSS a_1123_46634# a_1057_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1067 a_5700_37509# VSS VDAC_Pi VDD sky130_fd_pr__pfet_01v8_hvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1068 a_n4064_37440# a_n4334_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1069 VSS a_13259_45724# a_18315_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1070 a_22737_37285# a_22527_39145# a_22629_38406# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1071 a_n1453_44318# a_n1899_43946# a_n1549_44318# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1072 VSS a_22400_42852# a_22848_40081# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1073 VSS a_22223_43396# a_13887_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1074 a_11682_45822# a_11322_45546# a_11525_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1075 VDD a_22591_45572# a_19963_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1076 a_5934_30871# a_8791_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1077 a_18429_43548# a_18525_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X1078 a_509_45822# a_n1099_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X1079 a_20980_44850# a_20766_44850# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1080 a_4190_30871# a_19332_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1081 a_3381_47502# a_2905_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1082 VDD a_3537_45260# a_4649_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1083 a_6682_46660# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X1084 a_20273_45572# a_20107_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1085 VDD a_11963_45334# a_11787_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X1086 VDD a_1423_45028# a_9838_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1087 a_19256_45572# a_18175_45572# a_18909_45814# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1088 a_n755_45592# a_n809_44244# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1089 VSS a_3699_46634# a_3633_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1090 VSS a_5937_45572# a_9159_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1091 a_14226_46987# a_14180_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X1092 VSS a_n2438_43548# a_n2157_46122# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1093 VSS a_8953_45546# a_9241_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1094 a_n2840_45002# a_n2661_45010# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1095 a_n722_43218# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1096 a_12005_46436# a_2063_45854# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1097 a_9885_43396# a_8270_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1098 VSS a_n4209_37414# a_n4251_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X1099 VDD a_n3690_39616# a_n3420_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X1100 a_18817_42826# a_18599_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1101 VDD a_167_45260# a_1423_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1102 VDAC_Pi VSS a_5700_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1103 VSS a_4704_46090# a_1823_45246# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1104 a_16886_45144# a_8696_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X1105 a_11688_45572# a_11652_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X1106 a_8953_45002# CLK VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1107 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1108 a_4520_42826# a_1823_45246# a_4743_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1109 a_949_44458# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1110 a_n3420_39072# a_n3690_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1111 VSS a_22889_38993# a_22944_39857# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1112 VIN_P EN_VIN_BSTR_P a_n1057_35014# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1113 VDD a_n2104_42282# a_n3674_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1114 VDD RST_Z a_14311_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1115 a_19721_31679# a_22959_45036# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1116 a_458_43396# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X1117 a_19339_43156# a_19164_43230# a_19518_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1118 a_11453_44696# a_17719_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1119 VDD a_n3420_37984# a_n2860_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X1120 a_13711_45394# a_12891_46348# a_13348_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X1121 a_16664_43396# a_16547_43609# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1122 a_1138_42852# a_791_42968# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X1123 a_21259_43561# a_4190_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1124 a_10586_45546# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1125 VSS a_11599_46634# a_15599_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1126 VSS a_n3690_38528# a_n3420_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1127 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1128 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X1129 a_196_42282# a_375_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1130 VSS a_n881_46662# a_7989_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1131 a_7832_46660# a_7715_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1132 VDD a_n2109_45247# en_comp VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1133 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1134 a_15928_47570# a_15811_47375# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1135 a_3633_46660# a_2443_46660# a_3524_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1136 VSS a_n2472_45546# a_n2956_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1137 a_2127_44172# a_2675_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X1138 a_9885_43646# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X1139 a_n2472_43914# a_n2293_43922# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1140 VDD a_12991_46634# a_12978_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1141 VDD a_1667_45002# a_n863_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1142 a_n4209_39304# a_n2302_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1143 a_14084_46812# a_n1151_42308# a_14226_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X1144 a_5837_45028# a_3232_43370# a_5691_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X1145 a_21753_35474# a_19998_34978# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1146 VDD a_21195_42852# a_21671_42860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1147 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1148 a_12427_45724# a_12791_45546# a_12749_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1149 VSS a_n913_45002# a_4921_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1150 a_14209_32519# a_22591_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1151 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1152 a_12553_44484# a_12465_44636# a_n2661_43922# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1153 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1154 a_5829_43940# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X1155 a_16237_45028# a_n743_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X1156 VDD a_22959_45036# a_19721_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1157 a_14761_44260# a_14673_44172# a_n2293_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1158 VSS a_n1613_43370# a_5429_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1159 CAL_P a_22485_38105# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X1160 VSS a_21363_46634# a_21297_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1161 VDD a_n452_45724# a_n1853_46287# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1162 VDD a_584_46384# a_2998_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1163 VSS a_4699_43561# a_3539_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1164 VDD a_15959_42545# a_15890_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1165 VSS a_10227_46804# a_13157_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1166 a_n4209_38502# a_n2302_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X1167 VSS a_n2946_39866# a_n3565_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1168 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1169 a_17538_32519# a_22959_43948# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1170 a_n144_43396# a_n971_45724# a_n447_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X1171 a_16680_45572# a_15599_45572# a_16333_45814# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1172 VSS a_5937_45572# a_6101_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X1173 a_9672_43914# a_8199_44636# a_9895_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1174 a_15231_43396# a_9145_43396# a_15125_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1175 a_8387_43230# a_7871_42858# a_8292_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1176 VDD a_22731_47423# a_13717_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1177 VDD a_9290_44172# a_13667_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X1178 a_n3420_37984# a_n3690_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X1179 VDD a_10903_43370# a_13163_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.06615 ps=0.735 w=0.42 l=0.15
X1180 VDD a_17767_44458# a_17715_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X1181 VDD a_7845_44172# a_7542_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.28 ps=2.56 w=1 l=0.15
X1182 a_n2840_44458# a_n2661_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1183 a_22400_42852# a_22223_42860# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1184 VDD a_n863_45724# a_945_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X1185 VSS a_9482_43914# a_10157_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1186 VDD a_12549_44172# a_10949_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.195 ps=1.39 w=1 l=0.15
X1187 a_4933_42558# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1188 a_19333_46634# a_19466_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1189 a_13565_44260# a_12891_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1190 VSS a_n3690_37440# a_n3420_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1191 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1192 a_n2293_46098# a_5663_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X1193 EN_VIN_BSTR_P VDD a_n217_35014# VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.9
X1194 VSS a_11453_44696# a_22959_47212# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1195 VSS a_12563_42308# a_5534_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1196 a_n2472_42826# a_n2293_42834# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1197 a_7920_46348# a_8128_46384# a_8062_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1198 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1199 a_n13_43084# a_n443_42852# a_133_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1200 a_2698_46116# a_2521_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1201 a_15785_43172# a_15743_43084# a_15095_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X1202 a_8654_47026# a_7577_46660# a_8492_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1203 VDD a_21363_46634# a_21350_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1204 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1205 VDD a_n809_44244# a_n822_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1206 a_766_43646# a_626_44172# a_458_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X1207 a_n784_42308# a_n961_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1208 a_12895_43230# a_12379_42858# a_12800_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1209 VSS a_805_46414# a_739_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1210 VSS a_8191_45002# a_8137_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1211 a_15959_42545# a_15803_42450# a_16104_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1212 a_5210_46482# a_5164_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X1213 a_11341_43940# a_3232_43370# a_11173_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.19825 ps=1.26 w=0.65 l=0.15
X1214 VDD a_7705_45326# a_7735_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1215 a_13720_44458# a_13661_43548# a_13940_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1216 a_2162_46660# a_2107_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X1217 VSS a_n4334_39392# a_n4064_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1218 a_n1423_42826# a_n1641_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1219 a_n2956_39304# a_n2840_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1220 VDD a_11415_45002# a_n2661_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1221 a_15037_43940# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X1222 VDD a_1606_42308# a_2351_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1223 a_2277_45546# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1224 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1225 a_6903_46660# a_6755_46942# a_6540_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X1226 VDD a_14180_45002# a_13017_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1227 a_3232_43370# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1228 VDD a_n2302_40160# a_n4315_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1229 VDD a_8199_44636# a_8191_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X1230 a_n4209_37414# a_n2302_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X1231 a_1576_42282# a_1755_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1232 a_7573_43172# a_7499_43078# a_7227_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1233 VSS a_21855_43396# a_13678_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1234 VDD a_18989_43940# a_19006_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1235 VSS a_6540_46812# a_6491_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1236 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1237 VDD a_22223_45572# a_19479_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1238 VIN_N EN_VIN_BSTR_N C0_dummy_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1239 VSS a_2903_42308# a_3080_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1240 VSS a_n863_45724# a_n906_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X1241 a_n2840_44458# a_n2661_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1242 a_22629_37990# a_22581_37893# CAL_P VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1243 a_3823_42558# a_3065_45002# a_3905_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1244 VSS a_2779_44458# a_1307_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X1245 VSS a_5263_45724# a_5204_45822# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1246 VDD a_2124_47436# a_1209_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1247 a_12925_46660# a_11735_46660# a_12816_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1248 VSS a_2957_45546# a_2905_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1249 a_376_46348# a_n743_46660# a_518_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X1250 a_11415_45002# a_4915_47217# a_14581_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1251 VDD a_7754_40130# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.5
X1252 a_n2104_42282# a_n1925_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1253 a_n2472_45002# a_n2293_45010# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1254 a_21398_44850# a_20679_44626# a_20835_44721# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1255 VDD a_16333_45814# a_16223_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1256 a_16241_44484# a_2711_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1257 a_3905_42865# a_5257_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1258 VSS a_8685_43396# a_15231_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1259 VSS a_10623_46897# a_10554_47026# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1260 a_13485_45572# a_12549_44172# a_13385_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X1261 C3_P_btm a_n4209_38216# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1262 VSS a_22959_45572# a_20447_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1263 a_22848_39857# a_22485_38105# a_22581_37893# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1264 VDD a_19987_42826# a_n2017_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.135 ps=1.27 w=1 l=0.15
X1265 a_9028_43914# a_9482_43914# a_9420_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X1266 VSS a_17973_43940# a_18079_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X1267 a_n2860_39072# a_n2956_39304# a_n2946_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X1268 a_9290_44172# a_13635_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1269 a_3059_42968# a_742_44458# a_2987_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1270 a_n452_44636# a_n467_45028# a_n310_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X1271 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1272 VDD a_768_44030# a_2711_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1273 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1274 VDD a_12281_43396# a_12563_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1275 VDD a_12741_44636# a_22959_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1276 a_8333_44734# a_3537_45260# a_8238_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X1277 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1278 a_17124_42282# a_17303_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1279 a_12156_46660# a_11813_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1280 VDD a_10809_44734# a_22959_46124# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1281 VSS a_1115_44172# a_n2293_45010# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.169 ps=1.82 w=0.65 l=0.15
X1282 a_5013_44260# a_1307_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1283 VDD a_n447_43370# a_n2129_43609# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1284 a_3357_43084# a_5257_43370# a_5565_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1285 a_1568_43370# a_1847_42826# a_1793_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1286 a_n967_43230# a_n2157_42858# a_n1076_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1287 a_11682_45822# a_10586_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X1288 a_18315_45260# a_15227_44166# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X1289 a_n2012_44484# a_n2129_44697# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1290 a_14543_43071# a_5534_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1291 a_16147_45260# a_17478_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1292 a_22848_40081# en_comp a_22589_40055# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1293 a_19963_31679# a_22591_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1294 a_n967_45348# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1295 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1296 VDD a_11599_46634# a_20107_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1297 VSS a_7276_45260# a_7227_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1298 a_1241_44260# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.102375 ps=0.965 w=0.65 l=0.15
X1299 VDD a_n809_44244# a_n755_45592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1300 VSS a_n815_47178# a_n785_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1301 a_n4334_40480# a_n4318_40392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1302 a_3175_45822# a_3090_45724# a_2957_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X1303 a_14621_43646# a_14579_43548# a_14537_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1304 VDD a_n2946_37984# a_n3565_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1305 VREF a_20205_31679# C4_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1306 VSS a_15227_44166# a_18900_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X1307 a_n310_44811# a_n356_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X1308 VDD a_16977_43638# a_16867_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1309 VDD a_15227_44166# a_17749_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X1310 a_3147_46376# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X1311 a_12638_46436# a_12594_46348# a_12379_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1312 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1313 VSS a_2324_44458# a_6298_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1314 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1315 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1316 a_21071_46482# a_15227_44166# a_20708_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X1317 a_n1059_45260# a_17499_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1318 VDD a_1273_38525# a_2684_37794# VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1319 a_961_42354# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1320 a_9127_43156# a_8952_43230# a_9306_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1321 VSS a_12741_44636# a_22959_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1322 VSS a_8349_46414# a_8283_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1323 VSS a_11787_45002# a_11652_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X1324 a_4223_44672# a_3537_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1325 a_509_45822# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1326 a_16119_47582# a_15673_47210# a_16023_47582# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1327 a_6452_43396# a_6293_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1328 VSS CLK a_8953_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1329 a_6194_45824# a_6472_45840# a_6428_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1330 a_3754_38802# a_7754_38636# VSS sky130_fd_pr__res_high_po_0p35 l=18
X1331 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1332 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1333 VDD a_n881_46662# a_11031_47542# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1334 VSS a_1209_47178# a_1239_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1335 a_15559_46634# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X1336 a_12429_44172# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1337 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1338 a_11229_43218# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1339 a_16020_45572# a_15903_45785# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1340 C3_P_btm a_5932_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1341 a_10149_42308# a_9290_44172# a_9803_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1342 VSS a_20708_46348# a_20411_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X1343 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1344 C9_N_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1345 a_10793_43218# a_10083_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1346 a_n863_45724# a_1667_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1347 a_13635_43156# a_13460_43230# a_13814_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1348 a_12379_46436# a_12594_46348# a_12638_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X1349 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1350 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1351 a_1209_43370# a_1049_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1352 a_2982_43646# a_3232_43370# a_2813_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1353 a_n443_46116# a_n901_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1354 a_21542_45572# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1355 VSS a_19647_42308# a_13258_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1356 a_18985_46122# a_18819_46122# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1357 VSS a_n1794_35082# a_18194_34908# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1358 a_12839_46116# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1359 VDD a_n2438_43548# a_2443_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1360 VDD a_9028_43914# a_8975_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1361 VDD a_17124_42282# a_4958_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1362 VSS a_10053_45546# a_9625_46129# VSS sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X1363 a_17639_46660# a_17609_46634# a_765_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1364 VSS a_380_45546# a_n356_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X1365 VSS a_20193_45348# a_21973_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1366 VSS a_196_42282# a_n3674_37592# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1367 VDD a_5257_43370# a_5826_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X1368 a_9803_42558# a_n97_42460# a_9885_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1369 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1370 VSS a_10227_46804# a_10553_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1371 VSS a_18597_46090# a_16375_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1372 VSS a_n913_45002# a_12281_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1373 a_12816_46660# a_11901_46660# a_12469_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1374 a_n3565_39590# a_n2946_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1375 a_20205_45028# a_18184_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1376 a_n3420_37984# a_n3690_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1377 VDD a_13259_45724# a_13667_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1378 a_n1736_42282# a_n1557_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1379 a_13747_46662# a_19386_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1380 VSS a_4791_45118# a_6165_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X1381 a_261_44278# a_n863_45724# a_175_44278# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1382 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1383 a_8325_42308# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1384 a_10623_46897# a_10467_46802# a_10768_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1385 a_17957_46116# a_765_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.208 ps=1.94 w=0.65 l=0.15
X1386 a_2675_43914# a_2998_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1387 a_18695_43230# a_18249_42858# a_18599_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1388 a_17613_45144# a_8696_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1389 a_n4318_39304# a_n2840_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1390 a_18799_45938# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1391 VSS a_19862_44208# a_20922_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.089375 ps=0.925 w=0.65 l=0.15
X1392 a_6151_47436# a_14311_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1393 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1394 VSS a_5129_47502# a_5063_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1395 VSS a_167_45260# a_2521_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1396 a_3733_45822# a_n755_45592# a_3638_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X1397 a_16333_45814# a_16115_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1398 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1399 a_1337_46116# a_1176_45822# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X1400 a_13163_45724# a_13527_45546# a_13485_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1401 a_8605_42826# a_8387_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1402 VDD a_4419_46090# a_n1925_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1403 a_n4209_38216# a_n2302_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1404 a_20712_42282# a_n357_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1405 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1406 a_1241_43940# a_1467_44172# a_1443_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1407 a_9145_43396# a_8791_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1408 VDD a_n961_42308# a_n784_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1409 a_7227_42852# a_n97_42460# a_7309_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1410 a_14976_45348# a_13059_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X1411 a_9863_47436# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X1412 a_743_42282# a_19692_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1413 a_4915_47217# a_12991_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1414 VSS a_12891_46348# a_12638_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1415 a_n3674_38680# a_n2840_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1416 VCM a_4958_30871# C9_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1417 VSS a_3539_42460# a_3065_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1418 a_17801_45144# a_17613_45144# a_17719_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X1419 VDD a_n4209_39590# a_n4334_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X1420 a_18787_45572# a_18341_45572# a_18691_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1421 a_10922_42852# a_10796_42968# a_10518_42984# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1422 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1423 a_3754_39964# a_7754_40130# VSS sky130_fd_pr__res_high_po_0p35 l=18
X1424 VDD a_n4334_40480# a_n4064_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1425 VDD a_526_44458# a_3232_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1426 a_n1794_35082# a_564_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1427 a_167_45260# a_2202_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1428 VDD a_11967_42832# a_20512_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1429 VDD a_16019_45002# a_15903_45785# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1430 a_2896_43646# a_n443_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1431 VSS a_9067_47204# DATA[4] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1432 a_n2312_38680# a_n2104_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1433 a_12005_46116# a_10903_43370# a_12005_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1434 a_n2288_47178# a_n2109_47186# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1435 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1436 a_14097_32519# a_22959_42860# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1437 a_6999_46987# a_3877_44458# a_6540_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1438 a_8199_44636# a_10355_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X1439 a_3429_45260# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1440 C8_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1441 a_4338_37500# VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.589 ps=4.42 w=1.9 l=0.15
X1442 a_9293_42558# a_9223_42460# a_8953_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X1443 VDD a_n452_47436# a_n815_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1444 VDD a_n2302_40160# a_n4315_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1445 a_14309_45348# a_2711_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1446 a_13807_45067# a_13556_45296# a_13348_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1447 a_2981_46116# a_2804_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1448 a_1176_45822# a_997_45618# a_1260_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X1449 a_4185_45028# a_3877_44458# a_4185_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1450 VDD a_13159_45002# a_n2661_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1451 VSS a_20269_44172# a_19319_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1452 a_n1655_43396# a_n1699_43638# a_n1821_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1453 a_16104_42674# a_15890_42674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1454 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1455 a_22731_47423# SMPL_ON_N VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1456 a_n722_46482# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1457 VSS a_n443_42852# a_997_45618# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1458 a_6945_45348# a_5205_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1459 a_21513_45002# a_21363_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1460 a_4791_45118# a_4743_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X1461 VSS a_1576_42282# a_1606_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1462 a_n1533_46116# a_n2157_46122# a_n1641_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1463 a_15227_44166# a_22000_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1464 a_n743_46660# a_n1021_46688# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1465 a_n4064_40160# a_n4334_40480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X1466 a_2075_43172# a_1307_43914# a_n913_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1467 VSS a_5205_44484# a_6756_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1468 VDD a_327_44734# a_375_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1469 VDD a_19321_45002# a_3090_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X1470 VSS a_3483_46348# a_13829_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X1471 VDD a_7754_40130# a_11206_38545# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X1472 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1473 VDD a_5937_45572# a_6671_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1474 VDD a_n863_45724# a_458_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X1475 VDD a_n4334_38304# a_n4064_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X1476 VDD a_526_44458# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1477 VDD a_1756_43548# a_1467_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.28 ps=2.56 w=1 l=0.15
X1478 VDD a_4791_45118# a_5066_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1479 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1480 a_20269_44172# a_20365_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X1481 VDD a_14976_45028# a_15227_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1482 VSS a_13904_45546# a_12594_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X1483 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1484 VSS a_8953_45546# a_8568_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X1485 VDAC_Pi a_3754_38470# a_4338_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1486 a_16112_44458# a_15227_44166# a_16335_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1487 VSS a_16327_47482# a_17021_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1488 a_n913_45002# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1489 VSS a_20974_43370# a_20749_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1490 a_16388_46812# a_17957_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1725 ps=1.345 w=1 l=0.15
X1491 VSS a_20159_44458# a_19321_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X1492 VDD a_9672_43914# a_2107_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1493 VSS a_22589_40599# a_22737_37285# VSS sky130_fd_pr__nfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X1494 a_n4318_37592# a_n1736_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1495 VSS a_6151_47436# a_8189_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1496 VDD a_12549_44172# a_17609_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1497 a_6229_45572# a_6194_45824# a_5907_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1498 VDD a_19700_43370# a_n97_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1499 a_6851_47204# a_6491_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1500 VDD a_19615_44636# a_18579_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X1501 a_8423_43396# a_n443_42852# a_8317_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1502 VDD a_7499_43078# a_8697_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1503 a_18799_45938# a_18175_45572# a_18691_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1504 a_1755_42282# a_n913_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1505 a_n1741_47186# a_12005_46116# a_12379_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X1506 VSS a_2324_44458# a_6298_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1507 VDD a_6765_43638# a_6655_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1508 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1509 a_n4209_39304# a_n2302_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X1510 VDD a_22223_47212# a_21588_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1511 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1512 a_685_42968# a_n443_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1513 a_10467_46802# a_11599_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1514 VDD a_n443_42852# a_15781_43660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X1515 a_17749_42852# a_17701_42308# a_17665_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1516 a_18599_43230# a_18249_42858# a_18504_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1517 CLK_DATA a_n2833_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X1518 VDD a_7920_46348# a_7715_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1519 a_3537_45260# a_7287_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1520 a_2809_45028# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X1521 a_7832_46660# a_7715_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1522 a_3873_46454# a_n881_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X1523 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1524 VSS a_4905_42826# a_4520_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X1525 a_6709_45028# a_6431_45366# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1526 VSS a_20202_43084# a_21421_42336# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1527 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1528 a_20623_43914# a_19321_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1529 a_20193_45348# a_18494_42460# a_20205_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1530 VSS a_9313_45822# a_11459_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X1531 a_n4318_39768# a_n2840_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1532 a_n443_42852# a_n901_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1533 a_6428_45938# a_5907_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1534 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1535 a_1273_38525# a_1107_38525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1536 a_n2104_46634# a_n1925_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1537 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1538 VSS a_7287_43370# a_3537_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1539 a_2987_42968# a_1847_42826# a_2905_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1540 a_11031_47542# a_4915_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1541 VSS a_12991_46634# a_12925_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1542 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1543 VDAC_Ni a_7754_38636# VSS sky130_fd_pr__res_high_po_0p35 l=18
X1544 VSS a_20894_47436# a_20843_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1545 a_13076_44458# a_9482_43914# a_13468_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X1546 a_10752_42852# a_10083_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1547 a_n1809_43762# a_n2433_43396# a_n1917_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1548 a_17970_44736# a_18248_44752# a_18204_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1549 a_5663_43940# a_5883_43914# a_5841_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X1550 a_n2302_38778# a_n2312_38680# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1551 a_16588_47582# a_15507_47210# a_16241_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1552 VSS a_4099_45572# a_3483_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1553 VSS a_14539_43914# a_16112_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X1554 a_16867_43762# a_16243_43396# a_16759_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1555 VDD a_1107_38525# a_1273_38525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1556 a_n745_45366# a_n746_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1557 a_10518_42984# a_10835_43094# a_10793_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1558 C2_P_btm a_n3420_37984# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1559 VIN_P EN_VIN_BSTR_P C5_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1560 a_n37_45144# a_n443_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1561 a_18287_44626# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1562 a_20159_44458# a_20362_44736# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1563 VSS a_11341_43940# a_22223_43948# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1564 VSS a_8530_39574# a_3754_38470# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1565 DATA[5] a_11459_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1566 a_6969_46634# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1567 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1568 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1569 a_18861_43218# a_18817_42826# a_18695_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1570 a_11322_45546# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1571 a_n3674_37592# a_196_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1572 a_n1809_43762# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1573 a_4419_46090# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X1574 VDD a_11189_46129# a_11133_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X1575 VDD a_7227_47204# DATA[3] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1576 a_n1076_46494# a_n1991_46122# a_n1423_46090# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1577 VSS a_7640_43914# a_7584_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1578 VSS a_21753_35474# SMPL_ON_N VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1579 a_15959_42545# a_15764_42576# a_16269_42308# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1580 a_16375_45002# a_18597_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1581 VDD a_n1699_44726# a_n1809_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1582 a_4235_43370# a_3935_42891# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X1583 a_21177_47436# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X1584 a_7418_45394# a_7229_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X1585 a_22000_46634# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1586 VDD a_7542_44172# a_7499_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1587 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1588 a_11309_47204# a_11031_47542# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1589 VDD a_1307_43914# a_3353_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1590 a_3905_42308# a_2382_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X1591 a_8483_43230# a_8037_42858# a_8387_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1592 a_n2104_46634# a_n1925_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1593 a_453_43940# a_175_44278# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1594 a_7281_43914# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X1595 a_9028_43914# a_9290_44172# a_9248_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1596 EN_VIN_BSTR_P VDD a_n1550_35448# VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.9
X1597 VDD a_n2302_38778# a_n4209_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1598 VDD a_4700_47436# a_3785_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1599 a_18909_45814# a_18691_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1600 a_15521_42308# a_15486_42560# a_15051_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1601 a_11551_42558# a_n97_42460# a_11633_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1602 VSS a_11459_47204# DATA[5] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1603 VDD a_15227_44166# a_15415_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X1604 VSS a_16327_47482# a_20397_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1605 a_n809_44244# a_n984_44318# a_n630_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1606 VDD a_8270_45546# a_9165_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1607 VDD a_948_46660# a_1123_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1608 VDD a_15009_46634# a_14180_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1609 a_20766_44850# a_20679_44626# a_20362_44736# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1610 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1611 a_13385_45572# a_10903_43370# a_13297_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X1612 VDD a_13777_45326# a_13807_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1613 VSS a_n755_45592# a_n39_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1614 a_14976_45028# a_14797_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X1615 VSS a_22589_40599# a_22537_40625# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1616 a_6886_37412# VDAC_Pi VDD VSS sky130_fd_pr__nfet_03v3_nvt ad=0.145 pd=1.58 as=0.0725 ps=0.79 w=0.5 l=0.5
X1617 a_6419_46482# a_6165_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X1618 VSS a_768_44030# a_5244_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1619 a_n2302_37690# a_n2810_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1620 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1621 VSS a_n2946_39072# a_n3565_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1622 VDD a_8199_44636# a_8336_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X1623 a_20623_45572# a_20273_45572# a_20528_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1624 VSS a_9396_43370# a_5111_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1625 a_n2312_39304# a_n1920_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1626 a_20009_46494# a_18819_46122# a_19900_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1627 a_n1190_44850# a_n2267_44484# a_n1352_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1628 a_7309_42852# a_5891_43370# a_7227_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1629 a_743_42282# a_13661_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1630 VSS a_n4064_40160# a_n2302_40160# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X1631 a_22397_42558# a_n913_45002# a_17303_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1632 a_12991_43230# a_12545_42858# a_12895_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1633 VSS a_3905_42865# a_5013_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1634 a_22765_42852# a_15743_43084# a_18184_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1635 a_7705_45326# a_7229_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1636 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1637 VSS a_10405_44172# a_8016_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1638 a_3065_45002# a_1823_45246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X1639 a_742_44458# a_n443_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1640 a_310_45028# a_n37_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1641 VDD a_3232_43370# a_2982_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1642 VDD a_526_44458# a_3905_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X1643 VSS a_18184_42460# a_20256_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.11375 ps=1 w=0.65 l=0.15
X1644 VDD a_16241_47178# a_16131_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1645 a_19466_46812# a_13747_46662# a_19929_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1646 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1647 a_20850_46482# a_19692_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X1648 VSS a_768_44030# a_9028_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X1649 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1650 a_12089_42308# a_11551_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1651 a_11173_43940# a_2063_45854# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1652 a_3457_43396# a_1414_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1653 VDD a_5907_46634# a_5894_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1654 a_8034_45724# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1655 a_5841_46660# a_4651_46660# a_5732_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1656 a_22000_46634# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1657 VSS a_3699_46348# a_3160_47472# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X1658 VSS a_22223_45036# a_18114_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1659 a_2437_43396# a_1568_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1660 VDD a_n2104_46634# a_n2312_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1661 a_2448_45028# a_2382_45260# a_n2293_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X1662 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1663 a_21167_46155# a_20916_46384# a_20708_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1664 a_22725_37990# a_22589_40055# a_22629_37990# VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X1665 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1666 a_5205_44484# a_5343_44458# a_5289_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1667 a_7499_43078# a_10083_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1668 a_948_46660# a_33_46660# a_601_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1669 VSS a_21005_45260# a_19778_44110# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1670 VDD a_n2302_37690# a_n4209_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1671 VSS a_13487_47204# a_768_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X1672 a_9241_46436# a_n237_47217# a_8049_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1673 a_15015_46420# a_14840_46494# a_15194_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1674 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1675 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1676 VDD a_20567_45036# a_12549_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1677 a_21398_44850# a_20640_44752# a_20835_44721# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1678 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1679 a_1823_45246# a_4704_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1680 a_5527_46155# a_5204_45822# a_5068_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1681 a_1606_42308# a_1576_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1682 VSS a_4235_43370# a_4181_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1683 VDD a_18783_43370# a_18525_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X1684 w_1575_34786# a_n1696_34930# EN_VIN_BSTR_P w_1575_34786# sky130_fd_pr__pfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1685 a_n881_46662# a_14495_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X1686 a_21188_45572# a_20107_45572# a_20841_45814# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1687 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1688 a_n1821_44484# a_n2267_44484# a_n1917_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1689 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1690 a_22944_39857# a_22613_38993# a_22848_39857# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1691 VCM a_5534_30871# C7_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X1692 VSS a_8270_45546# a_8192_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X1693 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1694 a_5891_43370# a_9127_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1695 VDD a_n863_45724# a_3059_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1696 VDD a_17609_46634# a_765_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1697 VSS a_n755_45592# a_3503_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1698 a_19237_31679# a_22959_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1699 a_12156_46660# a_11813_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1700 a_n4334_38528# a_n4318_38680# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1701 a_n901_43156# a_n1076_43230# a_n722_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1702 a_n2810_45028# a_n2840_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1703 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1704 a_16333_45814# a_16115_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1705 a_16795_42852# a_n97_42460# a_16877_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X1706 a_n913_45002# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1707 VDD a_21188_46660# a_21363_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1708 a_6905_45572# a_6151_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1709 a_14180_45002# a_13059_46348# a_14403_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X1710 a_16405_45348# a_16375_45002# a_16321_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1711 VDD a_5934_30871# a_8515_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1712 VREF a_19963_31679# C3_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1713 VDD a_3422_30871# a_22315_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1714 a_2123_42473# a_n784_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1715 VSS a_n1613_43370# a_n1287_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1716 VSS a_22223_43948# a_14401_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1717 EN_VIN_BSTR_P a_n1696_34930# w_1575_34786# w_1575_34786# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X1718 a_19518_43218# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1719 w_1575_34786# a_n1057_35014# w_1575_34786# w_1575_34786# sky130_fd_pr__pfet_01v8 ad=0.986 pd=7.38 as=0 ps=0 w=3.4 l=16.6
X1720 VSS a_20075_46420# a_20009_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1721 VSS a_16922_45042# a_16751_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1722 VDD a_3232_43370# a_11341_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.3925 ps=1.785 w=1 l=0.15
X1723 a_1049_43396# a_458_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1724 VDD a_1169_39587# COMP_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1725 VDD a_526_44458# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1726 VDD a_n237_47217# a_8270_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1727 a_1848_45724# a_n237_47217# a_1990_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1728 VDD a_14539_43914# a_12465_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1729 VDD a_n881_46662# a_7903_47542# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1730 VDD a_1666_39043# a_1169_39043# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1731 VSS a_n1696_34930# a_n1057_35014# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X1732 VDD a_n1423_46090# a_n1533_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1733 VDD a_5111_44636# a_5421_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X1734 a_20623_46660# a_20107_46660# a_20528_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1735 a_11778_45572# a_10193_42453# a_11688_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X1736 a_6347_46155# a_6165_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1737 a_4700_47436# a_n443_46116# a_4842_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X1738 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1739 VDD a_21359_45002# a_21101_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X1740 C4_P_btm a_n3565_38502# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1741 a_14113_42308# a_13575_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1742 VDD a_5755_42308# a_5932_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1743 a_10695_43548# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1744 a_4958_30871# a_17124_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1745 a_17333_42852# a_16795_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1746 VSS a_19339_43156# a_19273_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1747 a_8387_43230# a_8037_42858# a_8292_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1748 VDD a_n2840_44458# a_n4318_40392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1749 VDD a_15004_44636# a_14815_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1750 VSS a_16327_47482# a_18861_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1751 VSS a_1823_45246# a_3602_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X1752 VDD a_18780_47178# a_13661_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1753 a_n4334_37440# a_n4318_37592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1754 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1755 a_2455_43940# a_895_43940# a_2253_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1756 a_2680_45002# a_3065_45002# a_2809_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1757 a_13667_43396# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X1758 a_21381_43940# a_21115_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1759 a_380_45546# a_765_45546# a_509_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X1760 a_15781_43660# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X1761 a_16019_45002# a_16147_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.183625 pd=1.215 as=0.160875 ps=1.145 w=0.65 l=0.15
X1762 VDD a_3537_45260# a_4558_45348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X1763 a_12741_44636# a_6755_46942# a_16789_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1764 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1765 a_5534_30871# a_12563_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1766 VSS a_2324_44458# a_15682_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1767 VDD en_comp a_1107_38525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1768 VDD a_n473_42460# a_n1761_44111# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X1769 VSS a_7754_38470# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0 ps=0 w=2 l=0.15
X1770 a_20836_43172# a_20193_45348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1771 a_12895_43230# a_12545_42858# a_12800_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1772 VSS a_n2833_47464# CLK_DATA VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1773 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X1774 VDD a_1123_46634# a_584_46384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1775 a_726_44056# a_626_44172# a_644_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1776 a_6655_43762# a_6031_43396# a_6547_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1777 DATA[5] a_11459_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X1778 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X1779 a_2889_44172# a_1414_42308# a_3052_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1780 VDD a_3232_43370# a_3626_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1781 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X1782 a_5343_44458# a_7963_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1783 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1784 a_3483_46348# a_4099_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1785 a_9313_44734# a_5883_43914# a_9241_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X1786 a_2809_45028# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X1787 VDD a_6171_45002# a_11827_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1788 w_10694_33990# a_10890_34112# w_10694_33990# w_10694_33990# sky130_fd_pr__pfet_01v8 ad=0.493 pd=3.69 as=10.006 ps=72.76 w=3.4 l=16.6
X1789 VDD a_9625_46129# a_9569_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1176 ps=1.4 w=0.42 l=0.15
X1790 a_15567_42826# a_15227_44166# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1791 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X1792 a_2113_38308# a_2113_38308# a_2113_38308# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X1793 a_7_45899# a_n443_46116# a_n452_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X1794 a_n2810_45572# a_n2840_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1795 a_5732_46660# a_4817_46660# a_5385_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1796 a_5708_44484# a_3483_46348# a_5608_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X1797 VDD a_13259_45724# a_22397_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1798 a_11823_42460# a_15051_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.305 ps=2.61 w=1 l=0.15
X1799 VDD a_13507_46334# a_22765_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1800 a_13678_32519# a_21855_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X1801 a_5365_45348# a_5111_44636# a_4927_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1802 a_17021_43396# a_16977_43638# a_16855_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1803 VDD a_7227_47204# DATA[3] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1804 VREF_GND a_n4064_39616# C9_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1805 a_7989_47542# a_n237_47217# a_7903_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1806 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1807 a_19332_42282# a_19511_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1808 VSS a_6851_47204# a_7227_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X1809 a_13607_46688# a_6755_46942# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1810 a_4880_45572# a_526_44458# a_4808_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X1811 a_20922_43172# a_10193_42453# a_20836_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.091 ps=0.93 w=0.65 l=0.15
X1812 a_12978_47026# a_11901_46660# a_12816_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1813 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1814 VDD a_13720_44458# a_12607_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1815 VDD a_2952_47436# a_2747_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X1816 a_5147_45002# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1817 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1818 VDD a_14513_46634# a_14543_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1819 VDD a_21259_43561# a_16922_45042# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1820 VDD a_n4334_38528# a_n4064_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1821 VSS a_11459_47204# DATA[5] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1822 VDD a_21137_46414# a_21167_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1823 C9_N_btm a_17730_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1824 a_3905_42558# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X1825 VSS a_22959_47212# a_22612_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1826 a_383_46660# a_33_46660# a_288_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1827 VSS a_6755_46942# a_13556_45296# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1828 a_n4209_38216# a_n2302_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X1829 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1830 a_17061_44734# a_11691_44458# a_16979_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1831 a_4149_42891# a_2382_45260# a_3935_42891# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X1832 DATA[3] a_7227_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1833 VDD a_n755_45592# a_3318_42354# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X1834 VDD a_n443_46116# a_1427_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1835 VDD a_5497_46414# a_5527_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1836 a_5937_45572# a_5907_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1837 a_11323_42473# a_5742_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1838 VSS a_4921_42308# a_5755_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1839 a_21076_30879# a_22959_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1840 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X1841 VDD a_n2302_38778# a_n4209_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1842 a_n3565_39304# a_n2946_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1843 a_3699_46634# a_3524_46660# a_3878_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1844 VDD a_17583_46090# a_13259_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1845 VSS a_3600_43914# a_3499_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X1846 VSS a_n755_45592# a_3318_42354# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X1847 a_5111_44636# a_9396_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1848 a_17595_43084# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1849 a_13829_44260# a_13059_46348# a_13483_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X1850 a_18341_45572# a_18175_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1851 a_9290_44172# a_13635_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1852 a_12991_46634# a_12816_46660# a_13170_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1853 VSS a_2277_45546# a_2211_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1854 a_18429_43548# a_18525_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.5
X1855 VSS a_6453_43914# a_n2661_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1856 a_6773_42558# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1857 a_2253_44260# a_n443_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.102375 ps=0.965 w=0.65 l=0.15
X1858 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1859 a_9885_42558# a_7499_43078# a_9803_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1860 a_16414_43172# a_16137_43396# a_16245_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X1861 a_21811_47423# SINGLE_ENDED VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1862 a_2304_45348# a_n863_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X1863 a_3726_37500# a_6886_37412# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=0.15
X1864 a_13351_46090# a_13507_46334# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X1865 a_n4064_38528# a_n4334_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X1866 a_n1435_47204# a_n1605_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1867 a_n935_46688# a_n1151_42308# a_n1021_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1868 VSS a_12549_44172# a_17639_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.099125 ps=0.955 w=0.65 l=0.15
X1869 a_6977_45572# a_6598_45938# a_6905_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1870 VSS a_n23_44458# a_n89_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X1871 VSS a_n1177_43370# a_n1243_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1872 VDD a_13460_43230# a_13635_43156# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1873 VSS a_n913_45002# a_n967_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1874 VDD a_11525_45546# a_11189_46129# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X1875 VDD a_n755_45592# a_626_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1876 a_n1287_44306# a_n1331_43914# a_n1453_44318# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1877 VDD a_10227_46804# a_10768_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1878 a_n755_45592# a_n809_44244# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1879 a_895_43940# a_644_44056# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X1880 a_n699_43396# a_n1177_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1881 a_11136_42852# a_10922_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1882 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1883 VDD a_8568_45546# a_8162_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1884 VDD a_n4334_37440# a_n4064_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1885 a_11551_42558# a_n97_42460# a_11633_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1886 a_6293_42852# a_5755_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1887 a_n2840_42826# a_n2661_42834# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1888 a_16131_47204# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1889 a_14033_45572# a_3483_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X1890 a_5289_44734# a_4223_44672# a_5205_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1891 VSS a_n1736_42282# a_n4318_37592# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1892 VDD a_10083_42826# a_7499_43078# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1893 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1894 a_768_44030# a_13487_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1895 VDD a_11415_45002# a_22591_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X1896 VSS a_5147_45002# a_5708_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X1897 VIN_N EN_VIN_BSTR_N C8_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X1898 VDD a_13259_45724# a_14309_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X1899 VSS a_6886_37412# a_4338_37500# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=0.15
X1900 a_10053_45546# a_10490_45724# a_10210_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X1901 a_n4064_40160# a_n4334_40480# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1902 VDD a_19332_42282# a_4190_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1903 a_n998_43396# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1904 a_3090_45724# a_18911_45144# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1468 ps=1.34 w=1 l=0.15
X1905 VSS a_18287_44626# a_18248_44752# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1906 a_6671_43940# a_6109_44484# a_6453_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X1907 a_n1352_43396# a_n2433_43396# a_n1699_43638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1908 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1909 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1910 VDD a_n2302_37690# a_n4209_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1911 VDD a_n2946_37984# a_n3565_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1912 a_16131_47204# a_15507_47210# a_16023_47582# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1913 a_n23_44458# a_n356_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X1914 VSS a_2779_44458# a_1307_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1915 a_11750_44172# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1916 a_7845_44172# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1917 VIN_N EN_VIN_BSTR_N C1_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X1918 VSS a_6123_31319# a_7963_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1919 a_5907_46634# a_5732_46660# a_6086_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1920 a_8560_45348# a_8746_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X1921 a_19095_43396# a_13661_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X1922 a_21363_46634# a_21188_46660# a_21542_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1923 VSS a_n4315_30879# a_n4251_40480# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X1924 VSS a_n4064_39616# a_n2302_39866# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X1925 a_14180_46482# a_14035_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1926 a_n4064_37440# a_n4334_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X1927 a_18315_45260# a_18587_45118# a_18545_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1928 a_8349_46414# a_8016_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X1929 a_2537_44260# a_2479_44172# a_2127_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X1930 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1931 VSS a_3499_42826# a_3445_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1932 VDD a_3815_47204# a_4007_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1933 a_9306_43218# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1934 VDD a_6667_45809# a_6598_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1935 a_7230_45938# a_6511_45714# a_6667_45809# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1936 VDD a_2779_44458# a_1307_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X1937 a_8685_43396# a_8147_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X1938 VDD a_22400_42852# a_22589_40599# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1939 VDD a_1273_38525# a_1666_39043# VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1940 VSS VSS a_3726_37500# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.589 pd=4.42 as=0.3135 ps=2.23 w=1.9 l=0.15
X1941 COMP_P a_1169_39587# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1942 a_8270_45546# a_n237_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1943 a_15765_45572# a_15599_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1944 a_3992_43940# a_768_44030# a_3737_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X1945 a_3815_47204# a_3785_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1946 a_2063_45854# a_9863_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1947 VSS a_11415_45002# a_22591_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1948 a_6755_46942# a_15015_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1949 VDD a_19431_45546# a_19418_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1950 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1951 VSS a_14021_43940# a_22959_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1952 a_19328_44172# a_19478_44306# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1386 ps=1.08 w=0.42 l=0.15
X1953 VSS a_10227_46804# a_14537_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1954 a_21073_44484# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1955 VDD a_768_44030# a_726_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X1956 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1957 VDD a_13059_46348# a_15297_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X1958 VSS a_12465_44636# a_22223_47212# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1959 VDD a_n1352_43396# a_n1177_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1960 VDD a_19998_34978# a_21753_35474# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1961 VSS a_n863_45724# a_1067_42314# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1962 a_19164_43230# a_18083_42858# a_18817_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1963 a_383_46660# a_n133_46660# a_288_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1964 a_3524_46660# a_2443_46660# a_3177_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1965 a_13814_43218# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1966 VSS a_9127_43156# a_9061_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1967 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1968 a_n217_35014# a_n1696_34930# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X1969 VDD a_9482_43914# a_10157_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X1970 VSS a_12607_44458# a_12553_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1971 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X1972 VSS a_10903_43370# a_11963_45334# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1973 VSS a_17499_43370# a_17433_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1974 C1_P_btm a_1606_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X1975 VDD a_12427_45724# a_10490_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X1976 a_13213_44734# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1977 VSS a_14815_43914# a_14761_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1978 a_12513_46660# a_12469_46902# a_12347_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1979 VDD a_n2302_39072# a_n4209_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1980 VSS a_11323_42473# a_10807_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1981 a_18989_43940# a_18451_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X1982 VDD a_1209_43370# a_n1557_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1983 VSS a_8667_46634# a_8601_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1984 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1985 a_2889_44172# a_2998_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X1986 VSS a_7281_43914# a_7229_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X1987 VSS a_21195_42852# a_21671_42860# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1988 a_n2956_38680# a_n2472_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1989 VSS a_n699_43396# a_4743_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X1990 VDD a_n443_46116# a_2437_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1991 a_n3565_39590# a_n2946_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X1992 a_10553_43218# a_10518_42984# a_10083_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1993 a_16789_44484# a_14537_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1994 VSS a_13635_43156# a_13569_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1995 a_18834_46812# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X1996 a_10405_44172# a_7499_43078# a_10555_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.13325 pd=1.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X1997 a_n1151_42308# a_n1329_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X1998 VSS a_n2833_47464# CLK_DATA VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X1999 VSS a_18315_45260# a_18189_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X2000 a_n1917_43396# a_n2433_43396# a_n2012_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2001 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2002 a_n1441_43940# a_n2065_43946# a_n1549_44318# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2003 VDD a_17499_43370# a_17486_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2004 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2005 VDD a_22223_42860# a_22400_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2006 VDD a_3524_46660# a_3699_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2007 a_n1059_45260# a_17499_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2008 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2009 VSS a_12861_44030# a_17639_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2010 a_10765_43646# a_10695_43548# a_10057_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X2011 VDD a_12549_44172# a_20556_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2012 a_15890_42674# a_15803_42450# a_15486_42560# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X2013 VDD a_5815_47464# a_n1613_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2014 a_17433_43396# a_16243_43396# a_17324_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2015 VCM a_4958_30871# C9_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2016 a_11827_44484# a_3232_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2017 a_1847_42826# a_2351_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2018 VSS a_6151_47436# a_14955_47212# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2019 a_20205_31679# a_22223_46124# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2020 VSS a_15227_44166# a_15785_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2021 VDD a_1239_47204# a_1431_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2022 VDD a_8667_46634# a_8654_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2023 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2024 a_n452_45724# a_n443_46116# a_n310_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2025 a_700_44734# a_n746_45260# a_327_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X2026 a_19862_44208# a_13747_46662# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2027 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2028 a_10775_45002# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X2029 a_3232_43370# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2030 VDD a_22959_44484# a_19237_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2031 a_1115_44172# a_453_43940# a_1443_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2032 a_484_44484# a_n863_45724# a_327_44734# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X2033 a_n3690_38528# a_n3674_38680# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2034 VDD a_14543_43071# a_13291_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2035 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2036 a_20512_43084# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2037 VSS a_12549_44172# a_21205_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2038 a_20256_43172# a_20202_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.203125 ps=1.275 w=0.65 l=0.15
X2039 a_6761_42308# a_n913_45002# a_6773_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2040 a_6298_44484# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2041 a_n2840_42282# a_n2661_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2042 a_n2661_46098# a_1983_46706# a_2162_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2043 a_5429_46660# a_5385_46902# a_5263_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2044 VSS a_15368_46634# a_15312_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2045 VDD a_8685_43396# a_14955_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X2046 VDD a_16855_45546# a_16842_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2047 VSS a_5815_47464# a_n1613_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2048 a_11315_46155# a_11133_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2049 a_16522_42674# a_15803_42450# a_15959_42545# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X2050 a_1221_42558# a_1184_42692# a_1149_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X2051 a_20885_46660# a_20841_46902# a_20719_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2052 a_20719_45572# a_20273_45572# a_20623_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2053 a_1756_43548# a_1307_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X2054 a_14456_42282# a_14635_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2055 a_n2472_42826# a_n2293_42834# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2056 a_7276_45260# a_6709_45028# a_7418_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2057 VDD a_1823_45246# a_3232_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2058 a_n4315_30879# a_n2302_40160# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2059 a_3260_45572# a_3218_45724# a_2957_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X2060 a_n2497_47436# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2061 VSS a_3422_30871# a_22315_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2062 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2063 VDD a_10341_42308# a_11554_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2064 a_11280_45822# a_2063_45854# a_10907_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X2065 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2066 a_603_45572# a_310_45028# a_509_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X2067 a_15002_46116# a_13925_46122# a_14840_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2068 a_8746_45002# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2069 a_n906_45572# a_n971_45724# a_n1013_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X2070 a_11064_45572# a_10903_43370# a_10907_45822# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X2071 a_21205_44306# a_20935_43940# a_21115_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X2072 a_2479_44172# a_2905_42968# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X2073 a_12861_44030# a_18143_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2074 DATA[3] a_7227_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X2075 VDD a_n2840_46090# a_n2956_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2076 VDD a_6945_45028# a_22223_46124# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2077 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2078 a_13556_45296# a_6755_46942# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2079 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2080 VCM a_7174_31319# C0_dummy_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2081 VDD a_8199_44636# a_9377_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X2082 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X2083 a_n4334_39392# a_n4318_39304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2084 a_12710_44260# a_10903_43370# a_12603_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X2085 a_13777_45326# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2086 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2087 a_16522_42674# a_15764_42576# a_15959_42545# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X2088 a_14205_43396# a_13667_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196275 ps=1.33 w=0.65 l=0.15
X2089 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2090 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2091 VDD a_5732_46660# a_5907_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2092 a_6419_46155# a_5807_45002# a_6419_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2093 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X2094 a_n2860_39866# a_n2956_39768# a_n2946_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X2095 VDD a_13556_45296# a_13857_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2096 a_18533_44260# a_18326_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2097 a_n901_46420# a_n1076_46494# a_n722_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2098 a_5066_45546# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2099 a_12861_44030# a_18143_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2100 VSS a_11599_46634# a_18175_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2101 VSS a_13635_43156# a_9290_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2102 VSS a_11599_46634# a_18819_46122# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2103 a_n3690_37440# a_n3674_37592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2104 VSS a_n3690_39616# a_n3420_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2105 a_n2442_46660# a_n2472_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2106 VSS a_n1435_47204# a_13487_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X2107 VDD a_3147_46376# a_526_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X2108 a_8317_43396# a_n755_45592# a_8229_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2109 a_n3674_38216# a_n2104_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2110 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2111 a_n2312_40392# a_n2288_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2112 VDD a_n1079_45724# a_n1099_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.28 ps=2.56 w=1 l=0.15
X2113 VSS a_22591_44484# a_17730_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2114 a_n914_42852# a_n1991_42858# a_n1076_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2115 a_n97_42460# a_19700_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2116 VDD a_n809_44244# a_n755_45592# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2117 a_3877_44458# a_3699_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2118 VDD a_22537_40625# a_22725_37990# VDD sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X2119 a_n913_45002# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2120 a_15368_46634# a_15143_45578# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X2121 a_11206_38545# CAL_N a_4338_37500# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X2122 a_4905_42826# a_5379_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2123 VSS a_10467_46802# a_10428_46928# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2124 VSS a_3147_46376# a_526_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X2125 a_9313_45822# a_9049_44484# a_9159_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2126 a_21145_44484# a_20766_44850# a_21073_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X2127 VDD a_n4334_40480# a_n4064_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2128 VSS a_2680_45002# a_2274_45254# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X2129 VDD a_2324_44458# a_15682_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2130 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2131 a_22613_38993# a_22527_39145# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2132 a_10768_47026# a_10554_47026# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X2133 VSS a_21671_42860# a_3422_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2134 a_n785_47204# a_n815_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2135 a_5837_45028# a_5807_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X2136 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2137 C0_dummy_P_btm a_7174_31319# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2138 a_14537_43396# a_14358_43442# a_14621_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X2139 a_n3565_38216# a_n2946_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2140 a_n1736_43218# a_n1853_43023# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2141 a_6640_46482# a_5257_43370# a_6419_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X2142 VDD a_3090_45724# a_17786_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X2143 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2144 a_15493_43396# a_14955_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X2145 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2146 a_16877_42852# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X2147 a_9823_46482# a_9569_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X2148 VDD a_14021_43940# a_22959_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2149 VDD a_n3420_38528# a_n2860_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X2150 VSS a_10227_46804# a_12513_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2151 VDD a_3483_46348# a_17061_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2152 VSS a_17339_46660# a_19095_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2153 a_3699_46348# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X2154 VSS a_10533_42308# a_10723_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2155 VSS a_3537_45260# a_4223_44672# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2156 a_18214_42558# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X2157 VSS a_14537_43396# a_14180_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X2158 a_16501_45348# a_10193_42453# a_16405_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2159 VSS a_15743_43084# a_15567_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2160 VSS a_21259_43561# a_16922_45042# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2161 VSS a_n2840_46634# a_n2956_39768# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2162 a_9049_44484# a_8701_44490# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X2163 VDD a_2382_45260# a_3737_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2164 VDD a_n967_45348# a_n961_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2165 a_19615_44636# a_12861_44030# a_19789_44512# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2166 a_22589_40599# COMP_P VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2167 a_1273_38525# a_1107_38525# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2168 VSS a_1169_39043# comp_n VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2169 a_9863_46634# a_10150_46912# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X2170 VDD a_n881_46662# a_n745_45366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2171 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2172 VDD a_21496_47436# a_13507_46334# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X2173 a_n2109_45247# a_n2017_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2174 VSS a_n143_45144# a_n37_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2175 SMPL_ON_P a_n2002_35448# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2176 a_19418_45938# a_18341_45572# a_19256_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2177 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2178 VDD a_n2438_43548# a_n2433_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2179 VDD a_5907_45546# a_5937_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.135 ps=1.27 w=1 l=0.15
X2180 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2181 C5_P_btm a_n4209_38502# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2182 VSS a_n452_44636# a_n2129_44697# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X2183 a_n2472_42282# a_n2293_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2184 a_n4318_38680# a_n2472_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2185 a_5608_44484# a_5111_44636# a_5518_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X2186 VDD a_742_44458# a_700_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X2187 VDD a_n901_43156# a_n443_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2188 VSS a_768_44030# a_13720_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X2189 VSS a_7287_43370# a_7221_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2190 VDD a_327_47204# DATA[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2191 a_2609_46660# a_2443_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2192 a_n89_44484# a_n467_45028# a_n452_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X2193 VDD a_9290_44172# a_9801_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X2194 VSS a_n1613_43370# a_6809_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2195 a_n4064_39616# a_n4334_39616# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2196 a_556_44484# a_526_44458# a_484_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X2197 VDD a_n4334_39392# a_n4064_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2198 VSS a_4007_47204# DATA[2] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2199 VDD a_2324_44458# a_15682_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2200 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2201 a_2112_39137# a_1273_38525# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2202 VSS a_19328_44172# a_19279_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.1201 pd=1.085 as=0.169 ps=1.82 w=0.65 l=0.15
X2203 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X2204 VDD a_n3420_37440# a_n2860_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X2205 a_n3420_38528# a_n3690_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X2206 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2207 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2208 a_10554_47026# a_10467_46802# a_10150_46912# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X2209 a_11387_46155# a_n1151_42308# a_11315_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X2210 a_10341_43396# a_9803_43646# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2211 a_13887_32519# a_22223_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2212 VSS a_10227_46804# a_20885_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2213 C0_P_btm a_n3420_37440# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2214 VIN_P EN_VIN_BSTR_P C2_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2215 VSS a_16137_43396# a_18548_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X2216 a_n452_45724# a_n743_46660# a_n310_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2217 a_11682_45822# a_11652_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X2218 a_n443_42852# a_n901_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2219 VDD a_n2472_46090# a_n2956_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2220 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X2221 VDD a_11322_45546# a_11280_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X2222 VSS a_13747_46662# a_14495_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X2223 VDD a_10809_44734# a_n2661_42834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2224 C0_dummy_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2225 VSS a_n4209_39590# a_n4251_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X2226 VSS a_n1329_42308# a_n1151_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2227 a_3381_47502# a_2905_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2228 VDD a_18479_47436# a_13747_46662# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X2229 VSS a_n746_45260# a_261_44278# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2230 VDD a_n2302_39072# a_n4209_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2231 a_5649_42852# a_5111_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2232 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2233 a_11136_45572# a_3483_46348# a_11064_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X2234 VSS a_13249_42308# a_13904_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X2235 a_17486_43762# a_16409_43396# a_17324_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2236 VSS a_n913_45002# a_8325_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2237 VSS a_1307_43914# a_2675_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2238 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2239 a_3699_46634# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2240 VSS a_13259_45724# a_14797_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X2241 VSS a_2324_44458# a_949_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2242 a_20841_45814# a_20623_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2243 VIN_N EN_VIN_BSTR_N C9_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X2244 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2245 a_17639_46660# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2246 a_10341_42308# a_9803_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X2247 a_16327_47482# a_17591_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2248 a_19998_34978# VDD EN_VIN_BSTR_N VSS sky130_fd_pr__nfet_05v0_nvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.9
X2249 VSS a_2324_44458# a_15682_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2250 a_1260_45572# a_n755_45592# a_1176_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X2251 a_20397_44484# a_20362_44736# a_20159_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X2252 a_12991_46634# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2253 a_518_46155# a_472_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2254 a_n4064_39072# a_n4334_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X2255 VDD a_20841_45814# a_20731_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2256 a_9751_46155# a_9569_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X2257 a_1443_43940# a_1414_42308# a_1241_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2258 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=0.35
X2259 DATA[1] a_1431_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2260 VDD a_11823_42460# a_14033_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X2261 VSS a_n2840_42826# a_n3674_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2262 VSS a_3537_45260# a_5365_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.102375 pd=0.965 as=0.10725 ps=0.98 w=0.65 l=0.15
X2263 a_3065_45002# a_3318_42354# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X2264 a_n310_45899# a_n356_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2265 C8_P_btm a_n3420_39616# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2266 a_16327_47482# a_17591_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2267 VDD a_22591_46660# a_20820_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2268 a_n3420_37440# a_n3690_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X2269 a_8337_42558# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2270 VDD a_4646_46812# a_7411_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2271 a_11186_47026# a_10428_46928# a_10623_46897# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X2272 a_20273_46660# a_20107_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2273 VSS a_3877_44458# a_2382_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2274 VDD a_n1331_43914# a_n1441_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2275 VDD a_10835_43094# a_10796_42968# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2276 VSS a_5066_45546# a_9159_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2277 VSS a_12883_44458# a_12829_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2278 a_11341_43940# a_10729_43914# a_11257_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3925 pd=1.785 as=0.135 ps=1.27 w=1 l=0.15
X2279 VREF a_n4209_39590# C9_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2280 VSS a_564_42282# a_n1794_35082# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2281 a_12549_44172# a_20567_45036# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2282 VDD a_14456_42282# a_5342_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2283 a_645_46660# a_601_46902# a_479_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2284 VDD a_2063_45854# a_10809_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2285 VDD a_2127_44172# a_n2661_45010# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.26 ps=2.52 w=1 l=0.15
X2286 VDD a_10227_46804# a_16104_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X2287 a_12861_44030# a_18143_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2288 a_14513_46634# a_14180_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2289 a_n2840_46090# a_n2661_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2290 a_5088_37509# VSS VDAC_Ni VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2291 a_21137_46414# a_19692_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2292 a_1609_45822# a_167_45260# a_1609_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2293 VREF_GND a_17730_32519# C9_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2294 a_14635_42282# a_n913_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2295 a_10544_45572# a_10490_45724# a_10053_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X2296 a_10555_44260# a_10949_43914# a_10405_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.1885 pd=1.88 as=0.13325 ps=1.06 w=0.65 l=0.15
X2297 C2_P_btm a_n3565_38216# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2298 VSS a_1431_47204# DATA[1] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2299 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2300 a_8952_43230# a_7871_42858# a_8605_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2301 a_3067_47026# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2302 a_9377_42558# a_8685_42308# a_9293_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2303 a_4190_30871# a_19332_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2304 VDD a_9067_47204# DATA[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2305 a_15861_45028# a_15595_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2306 a_15194_46482# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2307 a_6469_45572# a_5907_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X2308 a_13720_44458# a_9482_43914# a_14112_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X2309 a_15493_43940# a_14955_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2310 a_n1352_43396# a_n2267_43396# a_n1699_43638# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2311 a_16245_42852# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X2312 VSS a_n357_42282# a_6101_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2313 a_20692_30879# a_22959_46124# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2314 VSS a_n2302_37984# a_n4209_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2315 a_3177_46902# a_2959_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2316 a_5907_46634# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2317 a_5497_46414# a_5164_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2318 VSS a_104_43370# a_n971_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2319 VREF_GND a_13258_32519# C0_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2320 VDD a_4743_44484# a_4791_45118# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2321 a_19700_43370# a_18579_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2322 a_12861_44030# a_18143_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X2323 a_21363_46634# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2324 VSS a_n443_42852# a_15940_43402# VSS sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X2325 a_12427_45724# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.14075 ps=1.325 w=0.42 l=0.15
X2326 VSS a_n3690_39616# a_n3420_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X2327 a_5891_43370# a_9127_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2328 a_n1920_47178# a_n1741_47186# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2329 a_10903_43370# a_13351_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2330 a_n955_45028# a_n1059_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2331 SMPL_ON_P a_n2002_35448# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2332 VDD a_n357_42282# a_7309_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2333 VDD a_3147_46376# a_526_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2334 a_18596_45572# a_18479_45785# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2335 a_4185_45028# a_3065_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2336 a_6575_47204# a_6545_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2337 a_16137_43396# a_15781_43660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X2338 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2339 VSS a_22775_42308# a_22485_38105# VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2340 VSS a_n2472_46634# a_n2442_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2341 a_4649_42852# a_526_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2342 VSS a_2711_45572# a_20107_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2343 VSS a_n2104_42282# a_n3674_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2344 VSS a_15015_46420# a_14949_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2345 VSS a_5691_45260# a_n2109_47186# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2346 a_17583_46090# a_17715_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X2347 a_17730_32519# a_22591_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2348 a_3600_43914# a_1307_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X2349 VSS a_n1550_35448# a_n2002_35448# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2350 a_13925_46122# a_13759_46122# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2351 VDD a_n901_43156# a_n914_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2352 a_8191_45002# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X2353 VDD a_22959_46124# a_20692_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2354 a_n310_44484# a_n356_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X2355 a_21125_42558# a_18597_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2356 VDD a_1169_39587# COMP_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2357 a_5932_42308# a_5755_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2358 VSS a_14543_43071# a_13291_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2359 VDD a_1307_43914# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2360 VSS a_3147_46376# a_526_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2361 VDD a_n2946_38778# a_n3565_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2362 VDD a_16112_44458# a_14673_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X2363 a_n1641_46494# a_n1991_46122# a_n1736_46482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2364 a_3175_45822# a_3316_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2365 VSS a_16763_47508# a_5807_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2366 VREF a_20447_31679# C5_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2367 a_14226_46660# a_14180_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X2368 VDD a_13348_45260# a_13159_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X2369 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2370 VDD a_6491_46660# a_6851_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2371 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X2372 a_n4209_39590# a_n2302_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X2373 a_6511_45714# a_4646_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2374 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2375 VDD a_22775_42308# a_22485_38105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X2376 a_3422_30871# a_21671_42860# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2377 VSS a_16763_47508# a_16697_47582# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2378 VDD a_2889_44172# a_413_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.34 ps=2.68 w=1 l=0.15
X2379 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2380 VSS a_n443_42852# a_1755_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2381 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2382 a_10405_44172# a_10729_43914# a_10651_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X2383 a_n2840_45546# a_n2661_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2384 a_14401_32519# a_22223_43948# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2385 VREF a_21076_30879# C8_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2386 a_4558_45348# a_4574_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2387 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2388 a_5193_42852# a_3905_42865# a_5111_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2389 a_18143_47464# a_18479_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X2390 a_10533_42308# a_n913_45002# a_10545_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2391 VDD a_16721_46634# a_16751_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2392 a_18909_45814# a_18691_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2393 a_n2840_45002# a_n2661_45010# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2394 a_948_46660# a_n133_46660# a_601_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2395 a_3699_46348# a_3877_44458# a_3873_46454# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2396 a_117_45144# a_n443_42852# a_45_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X2397 a_11415_45002# a_13249_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2398 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2399 a_15681_43442# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2400 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2401 a_n4209_38502# a_n2302_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X2402 VREF_GND a_18114_32519# C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2403 VDD CAL_N VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=10
X2404 VDD a_n1059_45260# a_18727_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X2405 VSS a_5013_44260# a_5663_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2406 a_9801_43940# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2407 VSS a_10193_42453# a_18797_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2408 a_n4251_38304# a_n4318_38216# a_n4334_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X2409 a_2779_44458# a_1423_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2410 a_19789_44512# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X2411 VDD a_1107_38525# a_1273_38525# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2412 comp_n a_1169_39043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2413 VDD a_18057_42282# a_n356_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X2414 a_13113_42826# a_12895_43230# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2415 a_16197_42308# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X2416 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2417 VDD a_8034_45724# a_n1925_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X2418 VDD a_11691_44458# a_11649_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2419 VSS a_22581_37893# a_22537_39537# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2420 VSS a_n2002_35448# SMPL_ON_P VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2421 a_n3690_39392# a_n3674_39304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2422 a_15761_42308# a_15051_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X2423 a_16680_45572# a_15765_45572# a_16333_45814# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2424 VSS a_1568_43370# a_1512_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2425 VDD a_n1794_35082# a_n1696_34930# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2426 VDD a_5066_45546# a_5024_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X2427 VSS a_n809_44244# a_n875_44318# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2428 VDD a_n2946_37690# a_n3565_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2429 a_n2267_43396# a_n2433_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2430 a_10518_42984# a_10796_42968# a_10752_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X2431 VDD a_1123_46634# a_584_46384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2432 a_8189_46660# a_8145_46902# a_8023_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2433 VDD a_13661_43548# a_14976_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X2434 a_11691_44458# a_5807_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2435 VSS a_n4064_39072# a_n2302_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X2436 a_20062_46116# a_18985_46122# a_19900_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2437 a_20269_44172# a_20365_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X2438 VSS a_5891_43370# a_5837_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2439 VSS a_n2472_42826# a_n4318_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2440 VSS a_7754_38470# a_7754_38470# VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2441 a_18707_42852# a_18083_42858# a_18599_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2442 VDD a_327_47204# DATA[0] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2443 a_12638_46436# a_13059_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2444 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X2445 a_n784_42308# a_n961_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2446 a_13157_43218# a_13113_42826# a_12991_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2447 VSS a_4007_47204# DATA[2] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2448 VDD a_15015_46420# a_15002_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2449 VDD a_16327_47482# a_20159_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2450 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2451 VSS a_n785_47204# a_327_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X2452 a_18834_46812# a_13661_43548# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X2453 a_n2840_45546# a_n2661_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2454 VSS a_21177_47436# a_20990_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2455 VSS a_7499_43078# a_11816_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X2456 a_n3420_38528# a_n3690_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2457 a_6761_42308# a_3537_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2458 a_10623_46897# a_10428_46928# a_10933_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X2459 a_5263_45724# a_n881_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X2460 VDD a_11823_42460# a_11322_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2461 VSS a_5111_44636# a_8018_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X2462 a_7903_47542# a_n237_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2463 VSS a_8667_46634# a_n237_47217# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2464 a_3357_43084# a_4905_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2465 a_n2472_46090# a_n2293_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2466 VREF a_19237_31679# C0_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2467 SMPL_ON_N a_21753_35474# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2468 VCM a_5742_30871# C6_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2469 VSS a_22589_40055# a_22527_39145# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2470 VDD a_n901_43156# a_n443_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2471 VSS a_22959_46660# a_21076_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2472 a_10249_46116# a_9823_46155# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X2473 VDD a_10775_45002# a_10180_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X2474 CAL_N a_22485_38105# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X2475 a_2684_37794# VDAC_Pi a_2113_38308# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2476 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2477 a_8696_44636# a_16855_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X2478 a_n4209_37414# a_n2302_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X2479 a_13467_32519# a_21487_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2480 a_6633_46155# a_5807_45002# a_6419_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X2481 a_n2661_42834# a_8975_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2482 a_n1243_43396# a_n2433_43396# a_n1352_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2483 a_7274_43762# a_6197_43396# a_7112_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2484 a_10922_42852# a_10835_43094# a_10518_42984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X2485 DATA[0] a_327_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2486 VDD a_5807_45002# a_11691_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2487 a_n1917_43396# a_n2267_43396# a_n2012_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2488 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2489 a_n4209_38502# a_n2302_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2490 VSS RST_Z a_14311_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2491 a_16327_47482# a_17591_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.3 ps=2.6 w=1 l=0.15
X2492 a_18285_46348# a_18834_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2493 EN_VIN_BSTR_N a_18194_34908# w_10694_33990# w_10694_33990# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=0.66 ps=4.33 w=4 l=0.15
X2494 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2495 a_18597_46090# a_19431_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X2496 VSS a_18443_44721# a_18374_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X2497 VSS a_8199_44636# a_10951_45334# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2498 a_1176_45572# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X2499 a_7735_45067# a_6709_45028# a_7276_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X2500 C8_P_btm a_5342_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2501 DATA[4] a_9067_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2502 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=0.35
X2503 a_n3565_39304# a_n2946_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X2504 VSS a_n2109_45247# en_comp VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2505 a_n1076_43230# a_n1991_42858# a_n1423_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2506 DATA[1] a_1431_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X2507 a_13348_45260# a_13556_45296# a_13490_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2508 C10_P_btm a_n4064_40160# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2509 a_n2302_40160# a_n2312_40392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2510 VSS a_21356_42826# a_n357_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2511 VDD a_11453_44696# a_22959_47212# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2512 VSS a_15037_45618# a_15143_45578# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2513 VSS a_8696_44636# a_8701_44490# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2514 a_3878_46660# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2515 a_2277_45546# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2516 a_626_44172# a_n863_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2517 a_18479_45785# a_19268_43646# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.3275 ps=1.655 w=1 l=0.15
X2518 a_16327_47482# a_17591_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X2519 a_20273_45572# a_20107_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2520 a_10555_44260# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X2521 a_n3420_37440# a_n3690_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2522 VSS a_n443_42852# a_742_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2523 VSS a_n901_43156# a_n967_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2524 a_20820_30879# a_22591_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2525 VSS a_13076_44458# a_12883_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X2526 a_685_42968# a_n443_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2527 a_17364_32525# a_22959_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2528 a_13170_46660# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2529 a_11633_42558# a_9290_44172# a_11551_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2530 VDD a_4791_45118# a_6633_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X2531 a_20731_45938# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2532 a_19700_43370# a_18579_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2533 VDD a_11599_46634# a_20107_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2534 a_16751_45260# a_17023_45118# a_16981_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2535 a_2382_45260# a_3877_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2536 C9_N_btm a_21588_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2537 VSS a_13487_47204# a_768_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2538 a_12829_44484# a_12741_44636# a_n2293_43922# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2539 a_11257_43940# a_10807_43548# a_11173_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2540 VCM a_6123_31319# C4_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2541 VSS a_14084_46812# a_14035_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X2542 VDD a_5937_45572# a_8034_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2543 a_5342_30871# a_14456_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2544 a_17639_46660# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.099125 pd=0.955 as=0.169 ps=1.82 w=0.65 l=0.15
X2545 a_10809_44734# a_10057_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2546 VCM a_3422_30871# VDAC_P VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2547 VDD a_11823_42460# a_14853_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2548 a_20749_43396# a_20974_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2549 VDD a_11967_42832# a_16243_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2550 a_19511_42282# a_n913_45002# a_21125_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2551 VSS a_1431_47204# DATA[1] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2552 a_1609_45572# a_n443_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2553 a_17517_44484# a_16979_44734# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X2554 a_20075_46420# a_19900_46494# a_20254_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2555 a_n4209_37414# a_n2302_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2556 VDD a_10083_42826# a_7499_43078# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2557 a_16020_45572# a_15903_45785# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2558 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2559 a_20731_45938# a_20107_45572# a_20623_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2560 a_22629_38406# a_22581_37893# CAL_N VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X2561 VDD a_n3420_39072# a_n2860_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X2562 VSS a_22731_47423# a_13717_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2563 a_16855_45546# a_16680_45572# a_17034_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2564 a_18114_32519# a_22223_45036# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2565 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2566 a_17339_46660# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2567 a_n2472_45546# a_n2293_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2568 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2569 VSS a_18429_43548# a_16823_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2570 VSS a_n4334_38304# a_n4064_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2571 VSS a_8325_42308# a_8791_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2572 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2573 VDD a_n4334_38528# a_n4064_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2574 VSS a_768_44030# a_13076_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X2575 VSS a_12861_44030# a_19692_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2576 VDD a_14495_45572# a_n881_46662# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2577 a_18596_45572# a_18479_45785# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2578 a_n2472_45002# a_n2293_45010# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2579 VDD a_n881_46662# a_6431_45366# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2580 a_5326_44056# a_5147_45002# a_5244_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2581 VSS a_22959_42860# a_14097_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2582 a_3445_43172# a_3357_43084# a_n2293_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2583 a_13003_42852# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2584 VSS a_9127_43156# a_5891_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2585 a_3503_45724# a_3775_45552# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2586 C6_N_btm a_14401_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2587 a_19929_45028# a_19778_44110# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2588 a_3540_43646# a_584_46384# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2589 VSS a_n2302_37984# a_n4209_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2590 DATA[4] a_9067_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2591 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2592 VDD a_167_45260# a_117_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X2593 a_6086_46660# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2594 a_3147_46376# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X2595 a_n1533_46116# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2596 VSS a_n3565_38216# a_n3607_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X2597 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2598 a_5337_42558# a_5267_42460# a_4905_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X2599 a_21542_46660# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2600 a_10216_45572# a_10180_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X2601 a_4699_43561# a_3080_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2602 a_3626_43646# a_3232_43370# a_3457_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2603 a_n4064_37984# a_n4334_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X2604 VDD a_21613_42308# a_22775_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2605 a_16269_42308# a_15890_42674# a_16197_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X2606 a_1067_42314# a_1184_42692# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2607 VDD a_5937_45572# a_6945_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2608 COMP_P a_1169_39587# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2609 a_21356_42826# a_21381_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2610 VDD CLK a_8953_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2611 VDD a_2324_44458# a_949_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2612 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2613 VDD a_1307_43914# a_16237_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2614 a_n1549_44318# a_n2065_43946# a_n1644_44306# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2615 VSS a_19862_44208# a_19808_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2616 VDD a_5891_43370# a_8791_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2617 VSS a_n3690_39392# a_n3420_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2618 a_20256_43172# a_18494_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X2619 a_7927_46660# a_7411_46660# a_7832_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2620 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2621 VREF_GND a_13887_32519# C3_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2622 a_n3420_39072# a_n3690_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X2623 a_n2472_45546# a_n2293_45546# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2624 a_17668_45572# a_n881_46662# a_17568_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X2625 C9_P_btm a_n4064_39616# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2626 a_4649_42852# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2627 a_6540_46812# a_3877_44458# a_6682_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2628 VDD a_6511_45714# a_6472_45840# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2629 VSS a_15493_43396# a_19478_44306# VSS sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.08 as=0.0567 ps=0.69 w=0.42 l=0.15
X2630 a_16664_43396# a_16547_43609# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2631 VDD a_5068_46348# a_4955_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X2632 a_9159_44484# a_5883_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X2633 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2634 VSS a_10341_43396# a_22591_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2635 VDD a_n4334_37440# a_n4064_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2636 VSS a_17124_42282# a_4958_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2637 a_n1545_46494# a_n1991_46122# a_n1641_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2638 C8_P_btm a_n3565_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2639 a_5267_42460# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X2640 a_1138_42852# a_791_42968# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X2641 a_n4318_40392# a_n2840_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2642 a_n1644_44306# a_n1761_44111# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2643 VDD a_7754_40130# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=0 ps=0 w=8 l=0.5
X2644 VDD a_1609_45822# a_n2293_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X2645 a_5267_42460# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X2646 VREF_GND a_17364_32525# C7_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X2647 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2648 a_2127_44172# a_2675_43914# a_2455_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2649 a_11787_45002# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X2650 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2651 VDD a_17499_43370# a_n1059_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2652 a_n1057_35014# EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X2653 VSS a_19333_46634# a_19123_46287# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X2654 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2655 a_n2946_37984# a_n2956_38216# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2656 a_3316_45546# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X2657 VSS a_13777_45326# a_13711_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2658 a_20712_42282# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2659 a_19479_31679# a_22223_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2660 a_20573_43172# a_20512_43084# a_20256_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.118625 ps=1.015 w=0.65 l=0.15
X2661 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2662 a_n2293_46634# a_14673_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2663 a_n1177_43370# a_n1352_43396# a_n998_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2664 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2665 VSS a_526_44458# a_5457_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2666 a_33_46660# a_n133_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2667 a_584_46384# a_1123_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2668 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2669 VDD a_10903_43370# a_10849_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X2670 VDD a_7754_40130# a_7754_40130# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X2671 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X2672 a_8495_42852# a_7871_42858# a_8387_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2673 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2674 a_5495_43940# a_5244_44056# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X2675 a_16842_45938# a_15765_45572# a_16680_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2676 VDD a_167_45260# a_2521_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X2677 VDD a_2779_44458# a_1307_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2678 VSS a_n961_42308# a_n784_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2679 VSS a_13259_45724# a_17303_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2680 VDD a_5937_45572# a_5829_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X2681 a_17538_32519# a_22959_43948# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2682 a_21496_47436# a_4883_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2683 a_11816_44260# a_11750_44172# a_10729_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2684 a_9801_43940# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2685 a_5742_30871# a_10723_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2686 VDD a_15051_42282# a_11823_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2687 a_2123_42473# a_n784_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2688 a_13565_43940# a_12891_46348# a_13483_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2689 a_7227_42852# a_n97_42460# a_7309_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2690 a_5257_43370# a_5907_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2691 VDD a_13747_46662# a_13607_46688# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X2692 a_1667_45002# a_1823_45246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X2693 a_n1655_44484# a_n1699_44726# a_n1821_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2694 a_n2293_46098# a_5663_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1575 ps=1.315 w=1 l=0.15
X2695 a_13003_42852# a_12379_42858# a_12895_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2696 a_2711_45572# a_768_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2697 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X2698 DATA[0] a_327_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X2699 a_16763_47508# a_16588_47582# a_16942_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2700 a_4883_46098# a_21363_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2701 VSS a_16751_45260# a_6171_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X2702 VDD a_20835_44721# a_20766_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X2703 a_11750_44172# a_10903_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X2704 VSS a_15861_45028# a_17668_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X2705 a_7845_44172# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X2706 a_15597_42852# a_15743_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2707 a_n4064_39072# a_n4334_39392# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2708 VSS a_9223_42460# a_8953_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X2709 VDD a_11967_42832# a_18083_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2710 a_13487_47204# a_13381_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.16535 ps=1.82 w=0.65 l=0.15
X2711 a_13297_45572# a_13259_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1034 ps=1 w=0.42 l=0.15
X2712 C10_P_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2713 C2_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2714 w_10694_33990# a_10890_34112# w_10694_33990# w_10694_33990# sky130_fd_pr__pfet_01v8 ad=0.986 pd=7.38 as=0 ps=0 w=3.4 l=16.6
X2715 C10_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2716 VDD a_n3565_38216# a_n3690_38304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X2717 a_6101_43172# a_5891_43370# a_5755_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2718 a_11901_46660# a_11735_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2719 a_16979_44734# a_14539_43914# a_17061_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2720 VSS a_14955_47212# a_10227_46804# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2721 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2722 a_18443_44721# a_18248_44752# a_18753_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X2723 VDD a_18909_45814# a_18799_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2724 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2725 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2726 a_1431_46436# a_1138_42852# a_1337_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X2727 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2728 VDD a_n4064_37984# a_n2216_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X2729 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2730 a_18443_44721# a_18287_44626# a_18588_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X2731 VDD a_768_44030# a_5326_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X2732 VSS a_n4209_39304# a_n4251_39392# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X2733 a_n357_42282# a_21356_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2734 VSS a_n2288_47178# a_n2312_40392# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2735 a_491_47026# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2736 a_n901_46420# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2737 VSS a_3483_46348# a_15301_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2738 VCM a_1606_42308# C1_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2739 VDD a_20712_42282# a_10193_42453# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2740 VSS a_13635_43156# a_9290_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2741 a_5068_46348# a_5204_45822# a_5210_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2742 a_14033_45822# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X2743 VSS a_11599_46634# a_20107_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2744 a_3537_45260# a_7287_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2745 VSS a_6761_42308# a_7227_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2746 VDD a_13661_43548# a_15595_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2747 a_9803_42558# a_n97_42460# a_9885_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2748 VDD a_10227_46804# a_11136_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X2749 a_n1177_43370# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2750 VREF_GND a_n3420_39616# C8_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2751 VDD a_n2946_39072# a_n3565_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2752 a_601_46902# a_383_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2753 a_5024_45822# a_n443_46116# a_4419_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X2754 VDAC_Ni a_3754_38470# a_3726_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X2755 a_17701_42308# a_17531_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2756 VSS a_12861_44030# a_13487_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X2757 a_4808_45572# a_1823_45246# a_4419_46090# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X2758 a_6598_45938# a_6472_45840# a_6194_45824# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X2759 a_n229_43646# a_n2497_47436# a_n447_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X2760 a_n3607_38304# a_n3674_38216# a_n3690_38304# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X2761 VSS a_6969_46634# a_6903_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2762 a_18214_42558# a_18184_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X2763 a_491_47026# a_n133_46660# a_383_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2764 VSS a_4883_46098# a_10355_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X2765 VDD a_16327_47482# a_18588_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X2766 VDD a_4646_46812# a_6031_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2767 VSS a_n1613_43370# a_n1655_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2768 a_6812_45938# a_6598_45938# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X2769 a_8147_43396# a_n443_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X2770 VDAC_Ni VSS a_5088_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2771 a_12427_45724# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.1281 ps=1.03 w=0.42 l=0.15
X2772 C9_N_btm a_17730_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2773 VDD a_19594_46812# a_19551_46910# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X2774 a_n4318_37592# a_n1736_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2775 a_9290_44172# a_13635_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2776 VSS a_2698_46116# a_2804_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2777 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2778 a_1414_42308# a_1067_42314# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X2779 w_1575_34786# a_n1057_35014# w_1575_34786# w_1575_34786# sky130_fd_pr__pfet_01v8 ad=0.493 pd=3.69 as=0 ps=0 w=3.4 l=16.6
X2780 VSS a_5649_42852# a_22223_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2781 VDD a_13259_45724# a_14797_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2782 a_n2288_47178# a_n2109_47186# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X2783 a_4817_46660# a_4651_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2784 a_8062_46155# a_8016_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2785 a_949_44458# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2786 a_13296_44484# a_12891_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X2787 VDD a_20623_43914# a_20365_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X2788 a_11601_46155# a_11309_47204# a_11387_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
X2789 a_10210_45822# a_8746_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X2790 a_18287_44626# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2791 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2792 VSS a_11189_46129# a_11133_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X2793 a_n3565_38216# a_n2946_37984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X2794 a_6431_45366# a_5937_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2795 a_6109_44484# a_5518_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2796 a_14021_43940# a_13483_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X2797 a_17499_43370# a_17324_43396# a_17678_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2798 a_3495_45348# a_3429_45260# a_3316_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.182 ps=1.86 w=0.65 l=0.15
X2799 VDD a_1115_44172# a_n2293_45010# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.26 ps=2.52 w=1 l=0.15
X2800 VDD a_19787_47423# a_19594_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2801 a_18707_42852# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2802 a_19787_47423# START VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2803 a_8667_46634# a_8492_46660# a_8846_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2804 a_1208_46090# a_n881_46662# a_1431_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2805 a_5431_46482# a_n1151_42308# a_5068_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X2806 a_n1809_44850# a_n2433_44484# a_n1917_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2807 a_n2302_39866# a_n2442_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2808 VSS a_n2438_43548# a_2443_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2809 a_18797_44260# a_13661_43548# a_18451_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X2810 a_19551_46910# a_19692_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2811 VDD a_8953_45546# a_8049_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2812 a_8697_45822# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2813 VDD a_10341_43396# a_22591_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2814 a_12005_46116# a_2063_45854# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2815 VSS a_12861_44030# a_18911_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.194 pd=1.95 as=0.1092 ps=1.36 w=0.42 l=0.15
X2816 a_1241_43940# a_584_46384# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1575 ps=1.315 w=1 l=0.15
X2817 VSS a_2123_42473# a_1184_42692# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2818 a_1273_38525# a_1107_38525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2819 a_16285_47570# a_16241_47178# a_16119_47582# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2820 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2821 a_1423_45028# a_167_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2822 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2823 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X2824 a_10617_44484# a_10440_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2825 C7_P_btm a_n4064_39072# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X2826 VSS a_1169_39043# comp_n VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2827 VSS a_961_42354# a_1067_42314# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2828 VDD a_4704_46090# a_1823_45246# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2829 a_18479_47436# a_20075_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2830 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2831 VDD a_9313_45822# a_11459_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X2832 a_n1809_44850# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2833 VSS a_n3690_39392# a_n3420_39072# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X2834 a_19987_42826# a_10193_42453# a_20573_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X2835 VSS a_3785_47178# a_3815_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2836 VDD a_5891_43370# a_8375_44464# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2837 a_n3420_39072# a_n3690_39392# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2838 VSS a_9863_46634# a_2063_45854# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.08775 ps=0.92 w=0.65 l=0.15
X2839 a_7920_46348# a_n1151_42308# a_8062_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2840 VDD a_22889_38993# a_22581_37893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2841 a_19721_31679# a_22959_45036# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2842 a_19808_44306# a_19778_44110# a_19328_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2843 VDD a_10193_42453# a_11633_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2844 VDD a_15559_46634# a_13059_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2845 VDD a_11189_46129# a_11601_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X2846 a_5263_45724# a_5257_43370# a_5437_45600# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2847 a_12495_44260# a_12429_44172# a_10949_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.2275 ps=2 w=0.65 l=0.15
X2848 VSS a_n2840_43370# a_n4318_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2849 a_15037_43396# a_14205_43396# a_14955_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X2850 VSS a_4915_47217# a_12891_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2851 a_14084_46812# a_13885_46660# a_14226_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X2852 a_6452_43396# a_6293_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2853 VSS a_1107_38525# a_1273_38525# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2854 a_7705_45326# a_7229_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2855 a_8953_45002# CLK VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2856 a_16981_45144# a_16922_45042# a_16886_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X2857 a_1115_44172# a_1307_43914# a_1241_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2858 a_19478_44306# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1201 ps=1.085 w=0.42 l=0.15
X2859 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2860 a_4223_44672# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2861 a_7174_31319# a_20107_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2862 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2863 VDD a_n2302_39866# a_n4209_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2864 VDD a_10227_46804# a_15051_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2865 CLK_DATA a_n2833_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2866 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X2867 a_n2833_47464# a_n2497_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X2868 VSS a_8103_44636# a_7640_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X2869 a_15146_44811# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2870 a_n4209_39304# a_n2302_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2871 a_2903_45348# a_n971_45724# a_2809_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X2872 VSS a_3537_45260# a_8103_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2873 VSS a_21137_46414# a_21071_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2874 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2875 VSS a_1414_42308# a_2889_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2876 VDD a_1848_45724# a_1799_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X2877 VSS a_19279_43940# a_21398_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X2878 a_1666_39587# a_1273_38525# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X2879 VSS a_n13_43084# a_n1853_43023# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2880 a_18479_45785# a_19268_43646# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2881 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2882 VSS a_22485_44484# a_20974_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2883 VSS a_n3420_37984# a_n2946_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X2884 a_5275_47026# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2885 a_5841_44260# a_5495_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X2886 C5_N_btm EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2887 a_n2661_45546# a_4093_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2888 VSS a_n2302_38778# a_n4209_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2889 VSS a_5497_46414# a_5431_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X2890 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2891 VDD a_19339_43156# a_19326_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2892 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2893 a_8137_45348# a_8049_45260# a_n2293_42834# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2894 VDD a_17499_43370# a_n1059_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X2895 VDD a_6123_31319# a_7963_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2896 VDD a_12861_44030# a_17339_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2897 a_10849_43646# a_10807_43548# a_10765_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2898 VSS a_13507_46334# a_18997_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X2899 a_8560_45348# a_3483_46348# a_8488_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X2900 VDD a_n3690_38304# a_n3420_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2901 a_13249_42308# a_13070_42354# a_13333_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.135 ps=1.27 w=1 l=0.15
X2902 a_6969_46634# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2903 a_n2216_37984# a_n2810_45572# a_n2302_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X2904 VSS a_22223_46124# a_20205_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X2905 a_6194_45824# a_6511_45714# a_6469_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X2906 a_17613_45144# a_8696_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2907 a_n229_43646# a_n97_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2908 VSS a_n1613_43370# a_n1379_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2909 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2910 VSS a_13747_46662# a_19862_44208# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2911 a_17303_42282# a_n913_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2912 a_8649_43218# a_8605_42826# a_8483_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2913 VSS a_n901_46420# a_n967_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2914 a_15004_44636# a_13556_45296# a_15146_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X2915 a_11186_47026# a_10467_46802# a_10623_46897# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X2916 a_n1076_46494# a_n2157_46122# a_n1423_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2917 VSS a_526_44458# a_4169_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X2918 a_n23_45546# a_n356_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2919 a_3353_43940# a_2998_44172# a_2675_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2920 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2921 a_18326_43940# a_18079_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2922 a_20922_43172# a_19862_44208# a_20753_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1375 ps=1.275 w=1 l=0.15
X2923 a_10334_44484# a_10157_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2924 VSS a_742_44458# a_1756_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2925 C5_P_btm a_5934_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2926 a_n2017_45002# a_19987_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.208 ps=1.94 w=0.65 l=0.15
X2927 a_n2956_38216# a_n2472_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2928 VDD a_10193_42453# a_13657_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X2929 a_13885_46660# a_13607_46688# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2930 VDD a_8191_45002# a_n2293_42834# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2931 VSS RST_Z a_7754_39964# VSS sky130_fd_pr__nfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.15
X2932 VSS a_4223_44672# a_n2497_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2933 a_n217_35014# VDD EN_VIN_BSTR_P VSS sky130_fd_pr__nfet_05v0_nvt ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.9
X2934 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2935 a_4699_43561# a_3080_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2936 a_19511_42282# a_18597_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2937 a_n1991_46122# a_n2157_46122# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2938 a_n3420_37984# a_n3690_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X2939 VSS a_19692_46634# a_743_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2940 VDD a_22591_43396# a_14209_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X2941 VDD a_7499_43078# a_8746_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2942 a_n971_45724# a_104_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2943 a_22889_38993# a_22400_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2944 VDD a_n4334_39392# a_n4064_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X2945 a_20447_31679# a_22959_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X2946 VDD a_15493_43940# a_22959_43948# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2947 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2948 VSS a_n2302_37690# a_n4209_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2949 a_18147_46436# a_17339_46660# a_17957_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2950 a_8336_45822# a_8270_45546# a_n1925_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X2951 VDD a_13527_45546# a_13163_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X2952 a_n4334_39616# a_n4318_39768# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2953 a_n2956_39304# a_n2840_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2954 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2955 VDD a_584_46384# a_766_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1625 ps=1.325 w=1 l=0.15
X2956 w_10694_33990# a_18194_34908# EN_VIN_BSTR_N w_10694_33990# sky130_fd_pr__pfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X2957 a_11361_45348# a_10907_45822# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2958 VDD a_11599_46634# a_11735_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2959 a_19431_45546# a_19256_45572# a_19610_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2960 VSS a_9290_44172# a_12710_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.118125 pd=1.04 as=0.08775 ps=0.92 w=0.65 l=0.15
X2961 VDD a_11323_42473# a_10807_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2962 a_2266_47243# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X2963 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X2964 a_2982_43646# a_2479_44172# a_2896_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2965 a_18280_46660# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2966 VDD a_8492_46660# a_8667_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2967 C1_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X2968 VREF_GND a_n4064_40160# C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2969 VDD a_n1076_46494# a_n901_46420# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2970 a_n4251_38528# a_n4318_38680# a_n4334_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X2971 a_4361_42308# a_3823_42558# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X2972 VDD a_11967_42832# a_12379_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2973 VDD a_21811_47423# a_20916_46384# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2974 VDD a_11599_46634# a_13759_46122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2975 a_18985_46122# a_18819_46122# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2976 VDD a_n971_45724# a_3775_45552# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2977 VDD a_5649_42852# a_22223_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X2978 VSS a_5343_44458# a_8333_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2979 VDD a_7287_43370# a_3537_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2980 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2981 VSS a_3090_45724# a_10555_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.10725 ps=0.98 w=0.65 l=0.15
X2982 a_20528_45572# a_19466_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2983 a_13487_47204# a_13717_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2984 VREF_GND a_13678_32519# C2_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X2985 VDD a_22485_38105# a_22581_37893# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X2986 VDD a_20269_44172# a_19319_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X2987 a_5807_45002# a_16763_47508# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X2988 VSS a_16327_47482# a_16285_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2989 a_n23_44458# a_n356_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X2990 VDD a_n1059_45260# a_8791_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2991 a_1847_42826# a_2351_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2992 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X2993 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2994 VSS a_1169_39587# COMP_P VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2995 a_19553_46090# a_19335_46494# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2996 VDD a_n2840_45546# a_n2810_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2997 VSS a_3503_45724# a_3218_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X2998 a_15037_45618# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2999 a_14537_43646# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X3000 VDD a_1307_43914# a_n913_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3001 a_6671_43940# a_5205_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3002 a_n1699_43638# a_n1917_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3003 C6_P_btm a_n3420_39072# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3004 VDD a_n2946_38778# a_n3565_38502# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3005 VSS a_5111_44636# a_4905_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X3006 VDD a_9313_44734# a_22959_42860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3007 a_2124_47436# a_2063_45854# a_2266_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3008 VSS a_9625_46129# a_9569_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X3009 a_n4064_37984# a_n4334_38304# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3010 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3011 VDD a_19279_43940# a_21398_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X3012 VDD a_3483_46348# a_13565_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3013 a_22725_38406# a_22589_40055# a_22629_38406# VDD sky130_fd_pr__pfet_01v8 ad=0.0693 pd=0.75 as=0.0693 ps=0.75 w=0.42 l=0.15
X3014 a_6171_42473# a_5932_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3015 a_17568_45572# a_8696_44636# a_17478_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X3016 a_18588_44850# a_18374_44850# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X3017 a_18451_43940# a_18579_44172# a_18533_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3018 a_22485_38105# a_22775_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X3019 VSS a_5755_42308# a_5932_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3020 a_2959_46660# a_2609_46660# a_2864_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3021 a_21359_45002# a_21513_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3022 a_7_47243# a_n746_45260# a_n452_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3023 a_15227_46910# a_3090_45724# a_15009_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3024 a_14493_46090# a_14275_46494# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3025 a_19478_44306# a_15493_43396# a_19478_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0441 ps=0.63 w=0.42 l=0.15
X3026 a_7287_43370# a_7112_43396# a_7466_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3027 a_12251_46660# a_11901_46660# a_12156_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3028 a_8495_42852# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3029 a_n4251_37440# a_n4318_37592# a_n4334_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X3030 a_11633_42558# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X3031 VDD a_7276_45260# a_7227_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3032 VSS a_2479_44172# a_2813_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X3033 a_15279_43071# a_5342_30871# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3034 VREF_GND a_14401_32519# C6_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3035 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3036 VDD a_n815_47178# a_n785_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3037 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3038 a_1239_47204# a_1209_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3039 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3040 VDD a_3877_44458# a_3699_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3041 a_9313_45822# a_5937_45572# a_9241_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X3042 a_20841_45814# a_20623_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3043 VDD a_805_46414# a_835_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3044 a_12379_46436# a_12005_46116# a_n1741_47186# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3045 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3046 a_6298_44484# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3047 a_4338_37500# a_3754_38470# VDAC_Pi VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3048 a_961_42354# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3049 a_n2956_39768# a_n2840_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3050 a_n1741_47186# a_12594_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3051 VDD a_5257_43370# a_3905_42865# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3052 VSS en_comp a_1107_38525# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3053 VSS a_n473_42460# a_n1761_44111# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3054 a_13163_45724# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0987 pd=0.89 as=0.1281 ps=1.03 w=0.42 l=0.15
X3055 VDD a_10227_46804# a_9863_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3056 a_10210_45822# a_10586_45546# a_10053_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3057 comp_n a_1169_39043# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3058 VSS a_4185_45028# a_22959_45036# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3059 a_22485_38105# a_22775_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X3060 VDD a_n2438_43548# a_n2065_43946# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3061 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X3062 VSS a_n2002_35448# SMPL_ON_P VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3063 a_5457_43172# a_5111_44636# a_5111_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3064 VDD a_11787_45002# a_11652_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X3065 a_10695_43548# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X3066 VDD a_n1794_35082# a_n1696_34930# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3067 VDD a_n2946_37690# a_n3565_37414# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3068 a_13059_46348# a_15559_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3069 VDD a_n23_44458# a_7_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3070 a_12891_46348# a_4915_47217# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3071 a_8023_46660# a_7577_46660# a_7927_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3072 VSS a_10057_43914# a_9672_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X3073 a_n237_47217# a_8667_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.2087 ps=2.02 w=0.65 l=0.15
X3074 a_n143_45144# a_n755_45592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3075 a_20637_44484# a_20159_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X3076 a_4520_42826# a_4905_42826# a_4649_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3077 VSS a_n971_45724# a_8423_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.196275 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X3078 VSS RST_Z a_8530_39574# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3079 VSS a_n2946_37984# a_n3565_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3080 a_n1379_43218# a_n1423_42826# a_n1545_43230# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3081 a_8697_45822# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3082 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3083 VDD a_n4334_39616# a_n4064_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3084 VSS a_3626_43646# a_19647_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3085 a_n443_42852# a_n901_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3086 VDD a_1209_47178# a_1239_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3087 a_3094_47243# a_2905_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3088 a_15051_42282# a_15486_42560# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X3089 a_n1641_46494# a_n2157_46122# a_n1736_46482# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3090 VDD a_13661_43548# a_16241_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X3091 a_11823_42460# a_15051_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3092 a_5167_46660# a_4817_46660# a_5072_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3093 VSS a_10835_43094# a_10796_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3094 VDD a_20708_46348# a_20411_46873# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3095 VSS a_16327_47482# a_18005_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X3096 VSS a_16292_46812# a_15811_47375# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X3097 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3098 a_9482_43914# a_9838_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3099 a_20623_46660# a_20273_46660# a_20528_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3100 VDD a_12594_46348# a_n1741_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3101 a_18374_44850# a_18287_44626# a_17970_44736# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X3102 a_16750_47204# a_15673_47210# a_16588_47582# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3103 a_6545_47178# a_6419_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X3104 a_8783_44734# a_8696_44636# a_8701_44490# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3105 a_175_44278# a_n863_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3106 VDD a_22400_42852# a_22589_40055# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3107 VDD a_22223_43396# a_13887_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3108 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X3109 VSS a_n901_46420# a_n443_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3110 VDD a_18479_47436# a_20935_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X3111 VSS a_7754_38470# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0 ps=0 w=2 l=0.15
X3112 VSS a_5907_46634# a_5841_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3113 a_5745_43940# a_5883_43914# a_5829_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3114 a_3754_38470# a_7754_38470# VSS sky130_fd_pr__res_high_po_0p35 l=18
X3115 a_1110_47026# a_33_46660# a_948_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3116 a_16434_46987# a_16388_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3117 VSS a_2324_44458# a_15682_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3118 VDD a_n2302_39866# a_n4209_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3119 a_13381_47204# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3120 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3121 a_2998_44172# a_584_46384# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3122 a_20974_43370# a_22485_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3123 VDD a_4921_42308# a_5755_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3124 a_10991_42826# a_10835_43094# a_11136_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X3125 VDD a_6851_47204# a_7227_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3126 a_3052_44056# a_2998_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.14575 ps=1.335 w=0.42 l=0.15
X3127 VSS a_n4334_38528# a_n4064_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3128 a_3177_46902# a_2959_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3129 VSS a_1208_46090# a_472_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X3130 a_9241_44734# a_5937_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3131 a_n1699_43638# a_n1917_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3132 a_22365_46825# EN_OFFSET_CAL VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3133 VSS a_15682_46116# a_11599_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3134 VSS a_13163_45724# a_11962_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.1034 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3135 a_3055_46660# a_2609_46660# a_2959_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3136 a_19326_42852# a_18249_42858# a_19164_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3137 a_n443_46116# a_n901_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3138 a_9885_43646# a_8270_45546# a_9803_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3139 VDD a_18597_46090# a_16375_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3140 a_19431_45546# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3141 VSS a_22959_43396# a_17364_32525# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3142 w_10694_33990# a_10890_34112# w_10694_33990# w_10694_33990# sky130_fd_pr__pfet_01v8 ad=0.493 pd=3.69 as=0 ps=0 w=3.4 l=16.6
X3143 VDD a_n3690_38304# a_n3420_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X3144 a_n4064_39616# a_n4334_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X3145 VSS a_n1177_44458# a_n1243_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3146 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3147 VSS a_n23_45546# a_n89_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X3148 a_n452_47436# a_n746_45260# a_n310_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3149 a_2952_47436# a_n1151_42308# a_3094_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3150 VDD a_12816_46660# a_12991_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3151 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3152 a_7499_43940# a_7640_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3153 VSS a_n2302_38778# a_n4209_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3154 a_4235_43370# a_3935_42891# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15835 ps=1.395 w=1 l=0.15
X3155 a_5105_45348# a_4558_45348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.10725 ps=0.98 w=0.65 l=0.15
X3156 a_18051_46116# a_765_45546# a_17957_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.32 ps=2.64 w=1 l=0.15
X3157 a_n1441_43940# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3158 a_15301_44260# a_15227_44166# a_14955_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3159 a_n746_45260# a_n1177_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X3160 VSS a_n3565_38502# a_n3607_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X3161 a_n2840_43914# a_n2661_43922# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3162 a_6809_43396# a_6765_43638# a_6643_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3163 VSS a_376_46348# a_171_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X3164 a_19443_46116# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3165 VSS a_13059_46348# a_15143_45578# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3166 VSS a_8199_44636# a_8701_44490# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3167 a_7499_43940# a_3090_45724# a_7281_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3168 a_9165_43940# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3169 a_453_43940# a_175_44278# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X3170 a_9885_42308# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3171 a_n3674_39304# a_n2840_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3172 a_2959_46660# a_2443_46660# a_2864_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3173 a_14543_46987# a_13885_46660# a_14084_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3174 VDD a_413_45260# a_22959_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3175 a_17969_45144# a_16375_45002# a_17896_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
X3176 a_n4064_38528# a_n4334_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X3177 a_16292_46812# a_n743_46660# a_16434_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3178 a_21188_46660# a_20107_46660# a_20841_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3179 a_12251_46660# a_11735_46660# a_12156_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3180 a_4365_46436# a_4185_45028# a_n1925_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3181 a_n998_44484# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3182 VDD a_3177_46902# a_3067_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3183 a_7577_46660# a_7411_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3184 VDD a_n2472_45546# a_n2956_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3185 a_14976_45028# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X3186 a_10835_43094# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3187 a_12638_46436# a_12891_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.18525 ps=1.87 w=0.65 l=0.15
X3188 a_n1352_44484# a_n2433_44484# a_n1699_44726# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3189 a_n3420_37984# a_n3690_38304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3190 VSS a_13661_43548# a_743_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3191 a_12839_46116# a_12891_46348# a_n1741_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3192 VSS a_3090_45724# a_4927_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X3193 VSS a_22000_46634# a_15227_44166# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3194 VSS a_n863_45724# a_791_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X3195 a_14209_32519# a_22591_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3196 a_4646_46812# a_6298_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3197 VSS a_n4334_37440# a_n4064_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3198 a_n1613_43370# a_5815_47464# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3199 a_n2661_43922# a_12465_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3200 a_n2012_43396# a_n2129_43609# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3201 VSS a_11823_42460# a_14635_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3202 a_19692_46634# a_12549_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3203 C8_P_btm a_n3565_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3204 VSS a_4520_42826# a_4093_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X3205 a_5013_44260# a_3905_42865# a_5025_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3206 a_8018_44260# a_7499_43078# a_7911_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.125125 ps=1.035 w=0.65 l=0.15
X3207 VDD a_11823_42460# a_14358_43442# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X3208 a_167_45260# a_2202_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3209 a_20254_46482# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3210 VDD a_10405_44172# a_8016_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.335 ps=2.67 w=1 l=0.15
X3211 VIN_N EN_VIN_BSTR_N C10_N_btm VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X3212 a_742_44458# a_n443_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3213 VSS a_19332_42282# a_4190_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3214 a_14840_46494# a_13925_46122# a_14493_46090# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3215 VSS a_1414_42308# a_3457_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.091 ps=0.93 w=0.65 l=0.15
X3216 a_20356_42852# a_18184_42460# a_20256_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.175 ps=1.35 w=1 l=0.15
X3217 a_19006_44850# a_18287_44626# a_18443_44721# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X3218 a_9420_43940# a_768_44030# a_9165_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X3219 VDD a_10903_43370# a_12005_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3220 a_n4209_38216# a_n2302_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3221 VSS a_12861_44030# a_18280_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3222 VSS a_13661_43548# a_15685_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X3223 C4_P_btm a_6123_31319# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X3224 a_13575_42558# a_n97_42460# a_13657_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3225 VSS a_n2302_37690# a_n4209_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3226 a_8667_46634# a_6151_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3227 a_n1613_43370# a_5815_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3228 VDD a_n971_45724# a_n229_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3229 a_n1057_35014# a_n1696_34930# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3230 a_n1533_42852# a_n2157_42858# a_n1641_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3231 a_21335_42336# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3232 VSS a_n3565_37414# a_n3607_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.138125 pd=1.075 as=0.06825 ps=0.86 w=0.65 l=0.15
X3233 a_n2946_38778# a_n2956_38680# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3234 VSS a_9127_43156# a_5891_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X3235 VSS a_13351_46090# a_10903_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X3236 a_14309_45028# a_2711_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X3237 VSS a_413_45260# a_22959_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3238 a_743_42282# a_12549_44172# a_20749_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3239 VDD a_3877_44458# a_4185_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3240 a_13105_45348# a_13017_45260# a_n2661_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3241 VSS a_6545_47178# a_6575_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3242 a_8229_43396# a_7499_43078# a_8147_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X3243 a_19551_46910# a_19466_46812# a_19333_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3244 a_18280_46660# a_12549_44172# a_17609_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X3245 VSS a_18285_46348# a_18243_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.104 ps=0.97 w=0.65 l=0.15
X3246 a_6945_45028# a_5205_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3247 a_3726_37500# a_3754_38470# VDAC_Ni VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3248 a_n4064_37440# a_n4334_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X3249 a_20708_46348# a_20916_46384# a_20850_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3250 a_5167_46660# a_4651_46660# a_5072_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3251 VDD a_n1352_44484# a_n1177_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3252 a_15685_45394# a_15415_45028# a_15595_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3253 VDD a_10193_42453# a_18214_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X3254 a_21350_45938# a_20273_45572# a_21188_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3255 a_n2002_35448# a_n1550_35448# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3256 a_7639_45394# a_n1151_42308# a_7276_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X3257 VSS a_526_44458# a_10149_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3258 a_7765_42852# a_7227_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X3259 a_501_45348# a_413_45260# a_375_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3260 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3261 COMP_P a_1169_39587# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3262 a_16547_43609# a_16414_43172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25675 ps=1.44 w=0.65 l=0.15
X3263 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3264 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3265 a_n3565_38502# a_n2946_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3266 a_5891_43370# a_9127_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3267 a_13857_44734# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3268 a_n2661_46098# a_2107_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X3269 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3270 VSS a_16327_47482# a_18953_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3271 VSS a_742_44458# a_1568_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3272 a_19273_43230# a_18083_42858# a_19164_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3273 a_6123_31319# a_7227_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3274 a_768_44030# a_13487_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X3275 a_584_46384# a_1123_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3276 VDD a_2711_45572# a_4099_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3277 a_12293_43646# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3278 C8_N_btm a_5342_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3279 a_8035_47026# a_6151_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3280 a_10306_45572# a_10193_42453# a_10216_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X3281 a_18545_45144# a_13259_45724# a_18450_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X3282 a_n1917_44484# a_n2433_44484# a_n2012_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3283 a_22629_37990# a_22537_39537# CAL_P VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3284 a_n1423_46090# a_n1641_46494# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3285 a_16977_43638# a_16759_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3286 VDD a_21855_43396# a_13678_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3287 VDD a_6540_46812# a_6491_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X3288 VDD a_22223_43948# a_14401_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3289 VDD a_n863_45724# a_n1099_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3290 C10_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X3291 a_n2946_37690# a_n2956_37592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3292 a_5111_42852# a_4905_42826# a_5193_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3293 VDD a_5263_45724# a_5204_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X3294 a_n467_45028# a_n745_45366# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3295 VSS a_765_45546# a_1208_46090# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X3296 VDD a_15095_43370# a_14955_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X3297 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=0 ps=0 w=10 l=10
X3298 VSS a_n4334_38304# a_n4064_37984# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X3299 VDD a_2957_45546# a_2905_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3300 a_8855_44734# a_4791_45118# a_8783_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3301 a_11963_45334# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X3302 a_n2661_44458# a_11453_44696# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.182 ps=1.92 w=0.7 l=0.15
X3303 VDD a_4915_47217# a_11415_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3304 a_n1741_47186# a_12005_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3305 a_3600_43914# a_3537_45260# a_3820_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3306 a_21588_30879# a_22223_47212# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3307 a_1848_45724# a_2063_45854# a_1990_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3308 a_14537_46482# a_14493_46090# a_14371_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3309 a_10425_46660# a_9863_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X3310 a_16241_44734# a_2711_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X3311 a_3905_42865# a_5257_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3312 a_21811_47423# SINGLE_ENDED VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3313 a_19365_45572# a_18175_45572# a_19256_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3314 VDD a_22959_45572# a_20447_31679# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3315 a_3090_45724# a_18911_45144# a_19113_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3316 DATA[2] a_4007_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3317 a_13777_45326# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X3318 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3319 VCM a_5934_30871# C5_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3320 a_n3690_39616# a_n3674_39768# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3321 a_17333_42852# a_16795_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X3322 a_11525_45546# a_11962_45724# a_11682_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X3323 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3324 a_17595_43084# a_13259_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X3325 a_n13_43084# a_n755_45592# a_133_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11375 ps=1 w=0.65 l=0.15
X3326 a_n1696_34930# a_n1794_35082# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3327 a_19250_34978# a_18194_34908# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3328 a_n3565_37414# a_n2946_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3329 a_n2840_42282# a_n2661_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3330 a_20193_45348# a_18184_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3331 a_20719_46660# a_20273_46660# a_20623_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3332 a_1756_43548# a_768_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3333 VSS a_n1613_43370# a_n1379_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X3334 a_n2472_43914# a_n2293_43922# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3335 a_n2302_39072# a_n2312_39304# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3336 a_14456_42282# a_14635_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3337 VDD a_20075_46420# a_20062_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3338 VSS a_2711_45572# a_4099_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3339 a_4927_45028# a_5147_45002# a_5105_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X3340 a_21381_43940# a_21115_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X3341 SMPL_ON_N a_21753_35474# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3342 VSS a_10227_46804# a_10185_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X3343 a_n3607_38528# a_n3674_38680# a_n3690_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X3344 a_4169_42308# a_1823_45246# a_3823_42558# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3345 CLK_DATA a_n2833_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X3346 VDD a_20894_47436# a_20843_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X3347 a_4704_46090# a_4883_46098# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3348 VSS a_n913_45002# a_6761_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3349 VDD a_12465_44636# a_22223_47212# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3350 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3351 VDD a_15051_42282# a_11823_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3352 VDD a_20193_45348# a_20753_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3353 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3354 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X3355 VDD a_5257_43370# a_3357_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3356 VSS a_14113_42308# a_16522_42674# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X3357 a_22589_40055# en_comp VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3358 a_2324_44458# a_8953_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3359 VSS a_21753_35474# SMPL_ON_N VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3360 a_13460_43230# a_12379_42858# a_13113_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3361 a_19240_46482# a_19123_46287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3362 a_5829_43940# a_5495_43940# a_5745_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3363 a_10227_46804# a_14955_47212# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3364 VSS a_21487_43396# a_13467_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3365 VDD a_7287_43370# a_7274_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3366 VDD a_12861_44030# a_18911_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1468 pd=1.34 as=0.1092 ps=1.36 w=0.42 l=0.15
X3367 a_14955_43940# a_14537_43396# a_15037_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3368 a_15953_42852# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3369 a_9114_42852# a_8037_42858# a_8952_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3370 a_n4315_30879# a_n2302_40160# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X3371 VDD a_21753_35474# SMPL_ON_N VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3372 VSS a_n901_46420# a_n443_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3373 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3374 VSS a_8199_44636# a_8953_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X3375 a_18780_47178# a_18597_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3376 VDD a_15227_44166# a_18285_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3377 a_16375_45002# a_18597_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3378 VDD a_2324_44458# a_6298_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3379 a_15279_43071# a_5342_30871# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3380 a_10193_42453# a_20712_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3381 a_19335_46494# a_18985_46122# a_19240_46482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3382 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3383 a_5205_44484# a_5111_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3384 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3385 a_4842_47243# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3386 VSS a_685_42968# a_791_42968# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3387 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3388 VSS a_22591_45572# a_19963_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3389 C8_N_btm a_21076_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3390 a_509_45572# a_n1099_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X3391 VSS a_11322_45546# a_12016_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X3392 a_n1059_45260# a_17499_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3393 a_20753_42852# a_10193_42453# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X3394 DATA[5] a_11459_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3395 a_16789_45572# a_15599_45572# a_16680_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3396 a_20362_44736# a_20640_44752# a_20596_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X3397 a_13622_42852# a_12545_42858# a_13460_43230# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X3398 a_n1991_42858# a_n2157_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3399 a_15143_45578# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3400 VSS a_n746_45260# a_556_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X3401 a_8701_44490# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3402 a_n3607_37440# a_n3674_37592# a_n3690_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X3403 a_10775_45002# a_10951_45334# a_10903_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X3404 VSS a_7227_47204# DATA[3] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X3405 VDD a_6151_47436# a_14955_47212# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3406 a_15673_47210# a_15507_47210# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3407 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3408 VDD a_22589_40599# a_22537_40625# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3409 a_20679_44626# a_11967_42832# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3410 VDD a_n2946_39072# a_n3565_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3411 VDD a_10991_42826# a_10922_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X3412 a_5815_47464# a_6151_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X3413 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X3414 a_n2956_37592# a_n2472_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3415 a_13667_43396# a_11823_42460# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X3416 VSS a_n1920_47178# a_n2312_39304# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3417 VDD a_n4064_40160# a_n2216_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X3418 a_5164_46348# a_4927_45028# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.102375 ps=0.965 w=0.65 l=0.15
X3419 a_949_44458# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3420 a_15940_43402# a_12549_44172# a_15868_43402# VSS sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X3421 VDD a_4646_46812# a_4651_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3422 a_1427_43646# a_1049_43396# a_1209_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X3423 a_19164_43230# a_18249_42858# a_18817_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3424 VDD a_12861_44030# a_21845_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3425 a_2982_43646# a_3232_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.16 ps=1.32 w=1 l=0.15
X3426 w_1575_34786# EN_VIN_BSTR_P VDD w_1575_34786# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3427 VDD a_3600_43914# a_3499_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X3428 a_648_43396# a_526_44458# a_548_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.11375 ps=1 w=0.65 l=0.15
X3429 a_16409_43396# a_16243_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3430 VSS a_2063_45854# a_11136_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X3431 VSS a_1823_45246# a_2202_46116# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3432 a_10903_45394# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X3433 VDD a_n3420_39616# a_n2860_39866# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X3434 a_18243_46436# a_18189_46348# a_18147_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.10725 ps=0.98 w=0.65 l=0.15
X3435 VSS a_n971_45724# a_3775_45552# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3436 a_9290_44172# a_13635_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3437 a_4700_47436# a_4915_47217# a_4842_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3438 VDD a_6453_43914# a_n2661_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3439 VSS a_n2438_43548# a_n2433_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3440 a_11813_46116# a_11387_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11285 ps=1.045 w=0.65 l=0.15
X3441 VDD a_380_45546# a_n356_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X3442 VDD a_10053_45546# a_9625_46129# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X3443 VDD a_12861_44030# a_19615_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3444 a_2253_43940# a_n443_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1575 ps=1.315 w=1 l=0.15
X3445 VDD a_13113_42826# a_13003_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3446 a_765_45546# a_17609_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X3447 a_3503_45724# a_1823_45246# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X3448 VDD a_3699_46348# a_3160_47472# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X3449 VDD a_9625_46129# a_10037_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.07665 ps=0.785 w=0.42 l=0.15
X3450 VDD a_22223_45036# a_18114_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3451 a_18997_42308# a_18727_42674# a_18907_42674# VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3452 a_5755_42852# a_n97_42460# a_5837_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3453 VDAC_Pi VSS a_5700_37509# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3454 a_12281_43396# a_n913_45002# a_12293_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3455 VDD a_10533_42308# a_10723_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3456 VSS a_9863_47436# a_9804_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X3457 a_8049_45260# a_n237_47217# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3458 a_11387_46482# a_11133_46155# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X3459 VDD a_21005_45260# a_19778_44110# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X3460 VDD a_8791_42308# a_5934_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3461 VDD a_13487_47204# a_768_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3462 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X3463 a_895_43940# a_644_44056# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X3464 VSS a_n3420_38528# a_n2946_38778# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X3465 VDD a_4646_46812# a_7871_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3466 a_3067_47026# a_2443_46660# a_2959_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X3467 a_19256_45572# a_18341_45572# a_18909_45814# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3468 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3469 C3_P_btm a_n4064_37984# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X3470 VSS a_2713_42308# a_2903_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3471 a_9863_47436# a_2063_45854# a_10037_47542# VSS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X3472 a_15037_45618# a_13259_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3473 a_3726_37500# CAL_P a_11206_38545# VDD sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X3474 a_10991_42826# a_10796_42968# a_11301_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X3475 a_2127_44172# a_1307_43914# a_2253_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X3476 a_1823_45246# a_4704_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3477 VDD a_n2438_43548# a_n2433_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3478 a_17678_43396# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3479 a_n452_47436# a_n237_47217# a_n310_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3480 VDD a_10903_43370# a_12427_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.03 as=0.06615 ps=0.735 w=0.42 l=0.15
X3481 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3482 a_3080_42308# a_2903_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3483 a_22581_37893# a_22613_38993# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X3484 a_18057_42282# a_n1059_45260# a_18310_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X3485 VSS a_n452_45724# a_n1853_46287# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X3486 a_n3674_39768# a_n2472_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3487 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3488 a_8846_46660# a_6151_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3489 a_1307_43914# a_2779_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3490 a_22365_46825# EN_OFFSET_CAL VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3491 VDD CAL_P VDD VDD sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=0 ps=0 w=10 l=10
X3492 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3493 a_1273_38525# a_1107_38525# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3494 a_n89_45572# a_n743_46660# a_n452_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X3495 a_n2472_42282# a_n2293_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3496 VSS a_n2840_45002# a_n2810_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3497 a_15928_47570# a_15811_47375# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3498 a_518_46482# a_472_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X3499 a_15463_44811# a_11691_44458# a_15004_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3500 VSS a_17767_44458# a_17715_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X3501 a_20556_43646# a_19692_46634# a_20301_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3502 a_n3420_39616# a_n3690_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1775 ps=1.355 w=1 l=0.15
X3503 a_14309_45028# a_13059_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3504 a_16237_45028# a_16375_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3505 a_8791_43396# a_3537_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X3506 VDD a_22589_40599# a_22725_38406# VDD sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.46 as=0.0693 ps=0.75 w=0.42 l=0.15
X3507 VDD a_n4209_38216# a_n4334_38304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X3508 a_9061_43230# a_7871_42858# a_8952_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3509 a_1568_43370# a_n863_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3510 VDD a_n1423_42826# a_n1533_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3511 a_n1379_46482# a_n1423_46090# a_n1545_46494# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X3512 VSS a_n1794_35082# a_n1696_34930# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3513 a_13575_42558# a_n97_42460# a_13657_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3514 a_6667_45809# a_6511_45714# a_6812_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X3515 a_3754_39964# a_7754_39964# VSS sky130_fd_pr__res_high_po_0p35 l=18
X3516 VSS a_9290_44172# a_10586_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3517 a_16115_45572# a_15765_45572# a_16020_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3518 VDD a_18911_45144# a_3090_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.335 pd=1.67 as=0.165 ps=1.33 w=1 l=0.15
X3519 a_2725_42558# a_n755_45592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3520 a_18504_43218# a_17333_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3521 VDD a_3499_42826# a_n2293_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3522 a_16979_44734# a_14539_43914# a_17061_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3523 a_2253_43940# a_2479_44172# a_2455_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3524 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3525 VSS a_1307_43914# a_3681_42891# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.1092 ps=1.36 w=0.42 l=0.15
X3526 a_n310_47243# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3527 a_5025_43940# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3528 VSS a_626_44172# a_648_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.143 ps=1.09 w=0.65 l=0.15
X3529 VSS a_n3420_37440# a_n2946_37690# VSS sky130_fd_pr__nfet_01v8 ad=0.115375 pd=1.005 as=0.08775 ps=0.92 w=0.65 l=0.15
X3530 a_n3420_38528# a_n3690_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X3531 a_21356_42826# a_21381_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3532 a_16877_43172# a_16823_43084# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3533 a_20841_46902# a_20623_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3534 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X3535 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3536 VSS a_6171_45002# a_6125_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3537 VSS a_17595_43084# a_14539_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X3538 a_21137_46414# a_19692_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X3539 a_5883_43914# a_8333_44056# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X3540 a_20766_44850# a_20640_44752# a_20362_44736# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X3541 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3542 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3543 a_805_46414# a_472_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3544 a_1176_45822# a_997_45618# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.1925 ps=1.385 w=1 l=0.15
X3545 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3546 a_21887_42336# a_20202_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3547 VSS a_11967_42832# a_18083_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3548 DATA[2] a_4007_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X3549 VDD a_1823_45246# a_3316_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X3550 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3551 a_21513_45002# a_21363_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X3552 a_8704_45028# a_5937_45572# a_8191_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.195 ps=1.39 w=1 l=0.15
X3553 a_3232_43370# a_1823_45246# a_3363_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3554 a_13333_42558# a_13291_42460# a_13249_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3555 a_13661_43548# a_18780_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3556 a_5497_46414# a_5164_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X3557 a_12749_45572# a_12549_44172# a_12649_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0735 ps=0.77 w=0.42 l=0.15
X3558 VSS a_n2840_43914# a_n4318_39768# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3559 a_15037_44260# a_13556_45296# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3560 VSS a_22223_45572# a_19479_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3561 VDD a_n2438_43548# a_n133_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3562 VDD a_n984_44318# a_n809_44244# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3563 VDD a_14815_43914# a_n2293_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3564 a_n1545_43230# a_n1991_42858# a_n1641_43230# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3565 a_8128_46384# a_7903_47542# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3566 VDD a_7281_43914# a_7229_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3567 VDD a_13507_46334# a_18907_42674# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3568 CLK_DATA a_n2833_47464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3569 a_479_46660# a_33_46660# a_383_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3570 VSS a_6667_45809# a_6598_45938# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X3571 VDD a_13904_45546# a_12594_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X3572 VDD a_n881_46662# a_n1021_46688# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3573 VDD a_2324_44458# a_15682_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3574 a_8568_45546# a_8953_45546# a_8697_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3575 a_17767_44458# a_17970_44736# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X3576 VREF a_19479_31679# C1_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X3577 VCM a_4190_30871# C10_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3578 VDD a_n755_45592# a_133_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X3579 a_16241_44734# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3580 a_10867_43940# a_7499_43078# a_10405_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=1.41 as=0.195 ps=1.39 w=1 l=0.15
X3581 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3582 VDD a_10723_42308# a_5742_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3583 a_11823_42460# a_15051_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3584 a_20556_43646# a_20974_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3585 a_n3420_37440# a_n3690_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X3586 a_4574_45260# a_4791_45118# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X3587 a_13483_43940# a_13249_42308# a_13565_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3588 VDD a_20159_44458# a_19321_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X3589 a_n1352_44484# a_n2267_44484# a_n1699_44726# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3590 a_2583_47243# a_584_46384# a_2124_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3591 a_22612_30879# a_22959_47212# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3592 VDD a_8349_46414# a_8379_46155# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3593 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3594 VSS a_768_44030# a_2711_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3595 a_n2216_40160# a_n2312_40392# a_n2302_40160# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X3596 VSS a_14456_42282# a_5342_30871# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3597 a_n984_44318# a_n2065_43946# a_n1331_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3598 VREF a_22612_30879# C10_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3599 a_11608_46482# a_n1151_42308# a_11387_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X3600 a_5093_45028# a_5111_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.26 ps=2.52 w=1 l=0.15
X3601 VSS a_8953_45002# a_2324_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3602 a_19862_44208# a_13747_46662# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3603 VDD a_15227_44166# a_15597_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3604 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3605 a_19335_46494# a_18819_46122# a_19240_46482# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3606 VDD a_2324_44458# a_6298_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3607 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X3608 a_8953_45546# a_8685_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3609 a_n4318_38216# a_n2472_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3610 a_18249_42858# a_18083_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3611 a_12816_46660# a_11735_46660# a_12469_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3612 a_19268_43646# a_13661_43548# a_19177_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.1525 ps=1.305 w=1 l=0.15
X3613 a_13258_32519# a_19647_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3614 a_20256_42852# a_20202_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3125 ps=1.625 w=1 l=0.15
X3615 VDD a_16680_45572# a_16855_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X3616 VSS a_n447_43370# a_n2129_43609# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X3617 a_20528_45572# a_19466_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3618 a_11525_45546# a_10586_45546# a_11778_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X3619 VREF a_n3565_39590# C8_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3620 a_3537_45260# a_7287_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3621 VDD a_2711_45572# a_20107_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3622 a_16147_45260# a_17478_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3623 a_n2109_45247# a_n2017_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3624 a_19610_45572# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3625 a_19963_31679# a_22591_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3626 a_5837_43172# a_3537_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3627 a_n143_45144# a_n755_45592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3628 VDD a_18143_47464# a_12861_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X3629 VDD a_22959_47212# a_22612_30879# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3630 a_n310_45572# a_n356_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X3631 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3632 VSS a_7227_47204# DATA[3] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3633 a_15015_46420# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3634 VSS a_7227_45028# a_7230_45938# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X3635 a_20596_44850# a_20159_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X3636 a_2957_45546# a_3090_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X3637 VSS a_14579_43548# a_14537_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3638 VDD a_n2946_39866# a_n3565_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3639 VDD a_11599_46634# a_15507_47210# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3640 VDD a_6151_47436# a_6812_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X3641 VSS a_5111_44636# a_8333_44056# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3642 VDD a_7287_43370# a_3537_45260# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X3643 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3644 VDD a_20679_44626# a_20640_44752# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3645 a_n3565_39304# a_n2946_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3646 VDD COMP_P a_n1329_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X3647 VSS a_19321_45002# a_20567_45036# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3648 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3649 a_14513_46634# a_14180_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X3650 a_10903_43370# a_13351_46090# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3651 VSS a_n2472_45002# a_n2956_37592# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3652 a_10949_43914# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X3653 a_10149_43396# a_5111_44636# a_9803_43646# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X3654 VSS a_19431_45546# a_19365_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3655 VSS a_16922_45042# a_17719_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X3656 a_16112_44458# a_14539_43914# a_16241_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3657 a_13943_43396# a_11823_42460# a_13837_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X3658 C8_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X3659 VDD a_4099_45572# a_3483_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3660 a_6197_43396# a_6031_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3661 VSS a_18143_47464# a_12861_44030# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X3662 a_n2840_46634# a_n2661_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3663 a_380_45546# a_n357_42282# a_603_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X3664 a_18533_43940# a_18326_43940# a_18451_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3665 a_7309_42852# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X3666 VDD a_n863_45724# a_2448_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X3667 VSS a_1169_39587# COMP_P VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3668 a_5932_42308# a_5755_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3669 a_16328_43172# a_n97_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3670 VSS a_n2946_38778# a_n3565_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3671 a_17583_46090# a_17715_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X3672 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3673 VDD a_13635_43156# a_9290_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3674 VDD a_15433_44458# a_15463_44811# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3675 a_n2267_43396# a_n2433_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3676 VDD a_n755_45592# a_8147_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X3677 VSS a_10991_42826# a_10922_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X3678 a_5732_46660# a_4651_46660# a_5385_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3679 a_19615_44636# a_12549_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X3680 a_5088_37509# VDAC_P a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X3681 VDD a_5129_47502# a_5159_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3682 a_n2840_46090# a_n2661_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3683 a_n967_45348# a_n913_45002# a_n955_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3684 a_19006_44850# a_18248_44752# a_18443_44721# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X3685 a_n4209_39590# a_n2302_39866# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X3686 VDD a_18817_42826# a_18707_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3687 a_15559_46634# a_13507_46334# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X3688 a_9803_43646# a_8953_45546# a_9885_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3689 VDD a_3232_43370# a_9313_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X3690 VDD a_n2840_42282# a_n3674_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3691 a_13460_43230# a_12545_42858# a_13113_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3692 a_20362_44736# a_20679_44626# a_20637_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X3693 a_2713_42308# a_n913_45002# a_2725_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3694 a_768_44030# a_13487_47204# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3695 a_16241_47178# a_16023_47582# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X3696 a_14955_43396# a_14205_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X3697 VSS a_n913_45002# a_10533_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3698 a_7466_43396# a_n1613_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3699 a_n4064_40160# a_n4334_40480# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3700 VDD a_6151_47436# a_5907_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3701 a_16697_47582# a_15507_47210# a_16588_47582# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3702 a_n2267_44484# a_n2433_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3703 a_15682_43940# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3704 a_13693_46688# a_6755_46942# a_13607_46688# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X3705 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X3706 VDAC_Ni a_3754_38470# a_3726_37500# VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3707 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X3708 VDD a_19778_44110# a_19741_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3709 a_2609_46660# a_2443_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3710 a_5708_44484# a_5257_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.105625 ps=0.975 w=0.65 l=0.15
X3711 a_18143_47464# a_18479_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X3712 a_5263_46660# a_4817_46660# a_5167_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X3713 VSS a_n2472_43914# a_n3674_39768# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3714 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3715 a_12016_45572# a_11962_45724# a_11525_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X3716 VREF a_21588_30879# C9_N_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3717 VSS a_1107_38525# a_1273_38525# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3718 VSS a_18057_42282# a_n356_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X3719 VDD a_21671_42860# a_3422_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3720 VDD a_8746_45002# a_8704_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.105 ps=1.21 w=1 l=0.15
X3721 C9_N_btm a_4958_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3722 a_3411_47243# a_3160_47472# a_2952_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3723 a_n2840_46634# a_n2661_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3724 VSS a_7705_45326# a_7639_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X3725 VSS a_167_45260# a_1423_45028# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3726 a_11967_42832# a_15682_43940# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3727 VDD a_9396_43370# a_5111_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3728 a_743_42282# a_13661_43548# a_20301_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3729 a_n3420_39616# a_n3690_39616# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3730 a_133_43172# a_n357_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.10075 ps=0.96 w=0.65 l=0.15
X3731 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3732 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3733 VSS a_n2946_37690# a_n3565_37414# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3734 VDD a_20512_43084# a_19987_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
X3735 a_1891_43646# a_1307_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.14825 ps=1.34 w=0.42 l=0.15
X3736 VSS a_526_44458# a_2075_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3737 a_14485_44260# a_5807_45002# a_12465_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3738 a_n4318_39304# a_n2840_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3739 VIN_P EN_VIN_BSTR_P C8_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3740 VSS a_n357_42282# a_17141_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X3741 a_11453_44696# a_17719_45144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
X3742 VSS a_n1059_45260# a_8945_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X3743 a_17701_42308# a_17531_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3744 a_13657_42558# a_11823_42460# a_13575_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3745 a_10545_42558# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3746 a_8292_43218# a_7765_42852# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3747 a_16751_46987# a_5807_45002# a_16292_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X3748 a_10586_45546# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3749 a_n1243_44484# a_n2433_44484# a_n1352_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3750 VSS a_16855_45546# a_16789_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X3751 a_45_45144# a_n143_45144# a_n37_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X3752 VDD a_3537_45260# a_4223_44672# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3753 a_3626_43646# a_1414_42308# a_3540_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3754 VSS a_n2946_37984# a_n3565_38216# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3755 VDD a_20107_42308# a_7174_31319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X3756 a_3815_47204# a_3785_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3757 a_n1917_44484# a_n2267_44484# a_n2012_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3758 VCM a_5342_30871# C8_N_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3759 a_15567_42826# a_15743_43084# a_15953_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3760 VSS a_10341_42308# a_11554_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X3761 VSS a_4791_45118# a_6640_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X3762 a_6755_46942# a_15015_46420# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X3763 a_2437_43646# a_1568_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3764 VDAC_Pi a_7754_39632# VSS sky130_fd_pr__res_high_po_0p35 l=18
X3765 a_n3420_38528# a_n3690_38528# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3766 a_n4209_39590# a_n2302_39866# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3767 a_9823_46155# a_9804_47204# a_9823_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3768 a_1990_45899# a_167_45260# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3769 a_15743_43084# a_19339_43156# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X3770 a_5129_47502# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X3771 VDD a_5385_46902# a_5275_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3772 a_9145_43396# a_8791_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X3773 VDD a_20841_46902# a_20731_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3774 a_n2438_43548# a_949_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3775 VIN_P EN_VIN_BSTR_P C10_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3776 VDD a_n785_47204# a_327_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X3777 a_7276_45260# a_n1151_42308# a_7418_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X3778 a_8103_44636# a_8375_44464# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3779 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3780 a_4915_47217# a_12991_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X3781 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3782 a_21753_35474# a_19998_34978# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3783 VDD a_8199_44636# a_8855_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X3784 VDD a_12549_44172# a_21115_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X3785 VDD a_2553_47502# a_2583_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3786 a_n327_42558# a_n357_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.155 ps=1.31 w=1 l=0.15
X3787 a_12800_43218# a_12089_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3788 VSS a_20623_43914# a_20365_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.5
X3789 VSS a_n743_46660# a_16501_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X3790 VSS a_22959_45036# a_19721_31679# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3791 VSS a_11967_42832# a_16243_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3792 VDD a_7754_40130# a_11206_38545# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3793 a_n4318_38680# a_n2472_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3794 a_3363_44484# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3795 a_13483_43940# a_13249_42308# a_13565_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X3796 a_7754_40130# RST_Z VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3797 VDD a_4235_43370# a_n2661_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3798 a_n4209_38502# a_n2302_38778# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3799 a_13249_42558# a_10903_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X3800 a_18504_43218# a_17333_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3801 a_n39_42308# a_n97_42460# a_n473_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3802 a_10210_45822# a_10180_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X3803 VSS a_11967_42832# a_20512_43084# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3804 VSS a_n443_46116# a_2813_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3805 VSS a_4646_46812# a_7411_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3806 a_20273_46660# a_20107_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3807 VDD a_11341_43940# a_22223_43948# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3808 a_n2312_38680# a_n2104_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3809 VDD a_12791_45546# a_12427_45724# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0987 ps=0.89 w=0.42 l=0.15
X3810 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3811 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X3812 a_19237_31679# a_22959_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3813 VSS a_18194_34908# a_19250_34978# VSS sky130_fd_pr__nfet_01v8 ad=1.24 pd=8.62 as=0.66 ps=4.33 w=4 l=0.15
X3814 VDD a_19328_44172# a_19279_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16675 pd=1.435 as=0.26 ps=2.52 w=1 l=0.15
X3815 VDD SMPL_ON_P a_n1605_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3816 VSS a_11967_42832# a_12379_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3817 VSS a_15227_44166# a_17719_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3818 VDD a_18315_45260# a_18189_46348# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X3819 a_10951_45334# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X3820 VREF a_n4315_30879# C10_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3821 VDD a_2123_42473# a_1184_42692# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3822 a_4791_45118# a_4743_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X3823 a_21195_42852# a_20922_43172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25675 ps=1.44 w=0.65 l=0.15
X3824 a_4156_43218# a_3905_42865# a_3935_42891# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X3825 a_15227_44166# a_22000_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3826 a_n3420_37440# a_n3690_37440# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3827 a_n1899_43946# a_n2065_43946# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3828 VDD a_17591_47464# a_16327_47482# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X3829 a_n743_46660# a_n1021_46688# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3830 a_n2293_45546# a_2274_45254# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X3831 a_11633_42308# a_9290_44172# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X3832 a_15682_46116# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3833 a_20205_31679# a_22223_46124# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3834 a_n2472_46634# a_n2293_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3835 a_2698_46116# a_2521_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X3836 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X3837 VDD a_10193_42453# a_11682_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X3838 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3839 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X3840 VDD a_n3565_38502# a_n3690_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X3841 a_5342_30871# a_14456_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3842 VDD a_8325_42308# a_8791_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3843 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3844 a_548_43396# a_n863_45724# a_458_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.195 ps=1.9 w=0.65 l=0.15
X3845 VDD a_n4334_39616# a_n4064_39616# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X3846 VSS a_1756_43548# a_1467_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.182 ps=1.86 w=0.65 l=0.15
X3847 a_288_46660# a_171_46873# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X3848 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3849 VDD a_17517_44484# a_22591_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3850 VSS a_n913_45002# a_19511_42282# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3851 a_20894_47436# a_20990_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3852 a_15312_46660# a_14976_45028# a_15009_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X3853 a_n2472_46090# a_n2293_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3854 VDD a_n2438_43548# a_n2157_46122# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X3855 VSS a_22959_43948# a_17538_32519# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X3856 a_18194_34908# a_n1794_35082# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3857 C9_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X3858 VDD a_n4064_38528# a_n2216_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X3859 a_8037_42858# a_7871_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3860 a_n1736_43218# a_n1853_43023# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X3861 a_n4209_37414# a_n2302_37690# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3862 a_13527_45546# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3863 VDD a_n2472_42282# a_n4318_38216# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3864 a_n2661_43370# a_11415_45002# a_11361_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3865 VSS a_1273_38525# a_2113_38308# VSS sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X3866 VDD a_22165_42308# a_22223_42860# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3867 VDD a_n2840_42826# a_n3674_39304# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3868 VSS a_14180_45002# a_13017_45260# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X3869 a_15681_43442# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3870 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3871 C8_N_btm a_21076_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3872 VSS a_n2302_40160# a_n4315_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3873 a_8488_45348# a_8199_44636# a_8191_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.39325 ps=2.51 w=0.65 l=0.15
X3874 a_16588_47582# a_15673_47210# a_16241_47178# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3875 a_18220_42308# a_18184_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.167375 ps=1.165 w=0.65 l=0.15
X3876 a_n1423_46090# a_n1641_46494# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3877 VDD a_n1794_35082# a_18194_34908# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3878 VSS a_n4334_38528# a_n4064_38528# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X3879 VDD a_18143_47464# a_12861_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3880 a_17609_46634# a_12549_44172# a_18280_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3881 a_16115_45572# a_15599_45572# a_16020_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3882 VSS a_19700_43370# a_n97_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3883 VSS a_2124_47436# a_1209_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X3884 VREF_GND a_17730_32519# C9_N_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3885 a_15595_45028# a_15415_45028# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X3886 VDD a_6755_46942# a_12741_44636# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3887 VSS a_19615_44636# a_18579_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X3888 a_12545_42858# a_12379_42858# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3889 a_16942_47570# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X3890 a_8791_45572# a_7499_43078# a_8697_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3891 a_14853_42852# a_n913_45002# a_14635_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3892 a_n2438_43548# a_949_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3893 a_8333_44056# a_4223_44672# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3894 VSS a_4958_30871# a_17531_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3895 a_6511_45714# a_4646_46812# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3896 VDD a_10949_43914# a_10867_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.29 pd=2.58 as=0.205 ps=1.41 w=1 l=0.15
X3897 a_17973_43940# a_17737_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X3898 a_18494_42460# a_18907_42674# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X3899 a_17061_44734# a_15227_44166# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X3900 a_n2472_46634# a_n2293_46634# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3901 C2_P_btm a_3080_42308# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X3902 VSS a_5267_42460# a_4905_42826# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X3903 VSS a_n2438_43548# a_n2065_43946# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3904 VDD a_7754_40130# a_3754_38470# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3905 a_22629_38406# a_22537_39537# CAL_N VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1302 ps=1.46 w=0.42 l=0.15
X3906 VDD a_n357_42282# a_5837_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3907 a_9159_45572# a_5937_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X3908 a_3483_46348# a_4099_45572# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3909 a_8238_44734# a_8199_44636# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X3910 VSS a_17517_44484# a_22591_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3911 VDD a_n3565_37414# a_n3690_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X3912 VDD a_3381_47502# a_3411_47243# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3913 VSS a_21613_42308# a_22775_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X3914 COMP_P a_1169_39587# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3915 a_10150_46912# a_10467_46802# a_10425_46660# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X3916 a_526_44458# a_3147_46376# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3917 a_n2810_45572# a_n2840_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3918 a_13675_47204# a_n1435_47204# a_13569_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X3919 VSS a_11827_44484# a_22223_45036# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3920 a_5518_44484# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.175 ps=1.35 w=1 l=0.15
X3921 VDD a_n4064_37440# a_n2216_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X3922 a_22165_42308# a_21887_42336# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X3923 a_n3565_38502# a_n2946_38778# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X3924 a_5891_43370# a_9127_43156# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3925 a_13678_32519# a_21855_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3926 a_n2312_40392# a_n2288_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3927 VDD a_8605_42826# a_8495_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X3928 a_7499_43078# a_10083_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X3929 VDD a_20193_45348# a_21887_42336# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3930 a_18691_45572# a_18341_45572# a_18596_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3931 a_13076_44458# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X3932 a_3600_43914# a_1307_43914# a_3992_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X3933 VSS a_n4334_37440# a_n4064_37440# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X3934 a_4743_43172# a_3537_45260# a_4649_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3935 a_11387_46155# a_11309_47204# a_11387_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3936 a_n755_45592# a_n809_44244# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3937 a_15682_43940# a_2324_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X3938 VDD a_1666_39587# a_1169_39587# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3939 a_n1177_44458# a_n1352_44484# a_n998_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3940 a_11554_42852# a_10835_43094# a_10991_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X3941 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3942 VDD a_2680_45002# a_2274_45254# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X3943 C10_N_btm a_4190_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3944 VSS a_9313_44734# a_22959_42860# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3945 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X3946 VDD a_n1177_43370# a_n1190_43762# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3947 VDD a_6755_46942# a_13556_45296# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3948 a_n785_47204# a_n815_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3949 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3950 VDD a_n971_45724# a_8147_43396# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X3951 a_n4251_40480# a_n4318_40392# a_n4334_40480# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X3952 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X3953 VDD a_7754_40130# a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.5
X3954 a_19900_46494# a_18819_46122# a_19553_46090# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X3955 C9_P_btm a_n4209_39590# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X3956 a_12359_47026# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X3957 a_12561_45572# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1034 ps=1 w=0.42 l=0.15
X3958 a_10083_42826# a_10518_42984# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X3959 VSS a_10355_46116# a_8199_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3960 a_3422_30871# a_21671_42860# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X3961 a_5937_45572# a_5907_45546# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3962 a_21005_45260# a_21101_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.5
X3963 VDD a_16327_47482# a_17767_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X3964 a_12649_45572# a_10903_43370# a_12561_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0609 ps=0.71 w=0.42 l=0.15
X3965 VSS a_19321_45002# a_19113_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3966 a_5111_44636# a_9396_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3967 a_12469_46902# a_12251_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X3968 a_21297_45572# a_20107_45572# a_21188_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X3969 a_376_46348# a_584_46384# a_518_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X3970 a_15146_44484# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X3971 VIN_P EN_VIN_BSTR_P C6_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X3972 a_n1696_34930# a_n1794_35082# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3973 VDD a_n971_45724# a_n327_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2529 pd=2.52 as=0.16 ps=1.32 w=1 l=0.15
X3974 a_n3565_37414# a_n2946_37690# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X3975 a_14180_45002# a_14537_43396# a_14309_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X3976 VDD a_10193_42453# a_16237_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X3977 a_18681_44484# a_16327_47482# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X3978 VSS a_15009_46634# a_14180_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X3979 a_17829_46910# a_12549_44172# a_765_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1525 ps=1.305 w=1 l=0.15
X3980 a_2304_45348# a_2274_45254# a_2232_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.06825 ps=0.86 w=0.65 l=0.15
X3981 VDD a_1169_39043# comp_n VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3982 a_6598_45938# a_6511_45714# a_6194_45824# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X3983 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3984 a_n3565_38216# a_n2946_37984# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3985 a_5745_43940# a_5013_44260# a_5663_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X3986 VDD a_10193_42453# a_18533_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X3987 SMPL_ON_P a_n2002_35448# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3988 a_5742_30871# a_10723_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X3989 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3990 a_19478_44056# a_3090_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.16675 ps=1.435 w=0.42 l=0.15
X3991 a_10890_34112# EN_VIN_BSTR_N VIN_N VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X3992 VSS a_15051_42282# a_11823_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3993 a_10185_46660# a_10150_46912# a_9863_46634# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X3994 a_8192_45572# a_8199_44636# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.12675 ps=1.04 w=0.65 l=0.15
X3995 a_15890_42674# a_15764_42576# a_15486_42560# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X3996 a_10835_43094# a_11967_42832# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3997 VSS a_15682_43940# a_11967_42832# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3998 a_n699_43396# a_n1177_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X3999 a_14033_45822# a_3483_46348# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X4000 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4001 a_6101_44260# a_1307_43914# a_5663_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X4002 a_7927_46660# a_7577_46660# a_7832_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4003 a_21496_47436# a_4883_46098# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14075 ps=1.325 w=0.42 l=0.15
X4004 a_16721_46634# a_16388_46812# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4005 a_5826_44734# a_5147_45002# a_5518_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.22 ps=1.44 w=1 l=0.15
X4006 VDD a_16763_47508# a_16750_47204# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4007 VSS a_6298_44484# a_4646_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4008 VDD a_n746_45260# a_175_44278# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X4009 a_n443_46116# a_n901_46420# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4010 a_2813_43396# a_3232_43370# a_2982_43646# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4011 a_6171_42473# a_5932_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4012 VDD a_601_46902# a_491_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X4013 VSS a_4646_46812# a_6031_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4014 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4015 VDD a_1123_46634# a_1110_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4016 VSS a_13059_46348# a_12638_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.091 ps=0.93 w=0.65 l=0.15
X4017 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4018 a_11787_45002# a_11963_45334# a_11915_45394# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X4019 VSS a_584_46384# a_2998_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4020 a_8292_43218# a_7765_42852# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4021 VDD a_n2472_42826# a_n4318_38680# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4022 a_1667_45002# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X4023 VDD a_n3690_38528# a_n3420_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4024 a_20731_47026# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X4025 a_8062_46482# a_8016_46348# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4026 VDD a_6298_44484# a_4646_46812# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4027 a_n2216_38778# a_n2312_38680# a_n2302_38778# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X4028 VSS a_11599_46634# a_20107_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4029 a_13925_46122# a_13759_46122# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4030 VSS CLK a_8953_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X4031 VSS a_n2104_46634# a_n2312_38680# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4032 a_5385_46902# a_5167_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4033 a_n1177_44458# a_n1613_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4034 VDD a_7499_43078# a_10729_43914# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X4035 a_9803_43646# a_8953_45546# a_9885_43646# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4036 VDD a_19256_45572# a_19431_45546# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4037 a_7911_44260# a_7845_44172# a_7542_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.182 ps=1.86 w=0.65 l=0.15
X4038 VDD a_5111_44636# a_7542_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.135 ps=1.27 w=1 l=0.15
X4039 VDD a_6761_42308# a_7227_42308# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X4040 VDD a_19553_46090# a_19443_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X4041 a_n1641_43230# a_n2157_42858# a_n1736_43218# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4042 a_5205_44484# a_5343_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4043 a_22400_42852# a_22223_42860# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4044 a_12603_44260# a_12549_44172# a_12495_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.12675 ps=1.04 w=0.65 l=0.15
X4045 a_3638_45822# a_1823_45246# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X4046 a_17324_43396# a_16243_43396# a_16977_43638# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X4047 a_19452_47524# a_19386_47436# a_13747_46662# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4048 a_5275_47026# a_4651_46660# a_5167_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4049 VSS a_327_47204# DATA[0] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4050 a_11915_45394# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X4051 a_14447_46660# a_n1151_42308# a_14084_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4052 a_20731_47026# a_20107_46660# a_20623_46660# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4053 VSS a_n1613_43370# a_n1655_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X4054 a_12800_43218# a_12089_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4055 VDD a_8953_45002# a_2324_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4056 VDAC_N a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4057 VSS a_20712_42282# a_10193_42453# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4058 a_15720_42674# a_15051_42282# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4059 VSS a_n443_42852# a_421_43172# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X4060 a_14493_46090# a_14275_46494# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4061 VDD a_11599_46634# a_15599_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4062 a_n659_45366# a_n746_45260# a_n745_45366# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4063 a_15682_46116# a_2324_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X4064 a_n881_46662# a_14495_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X4065 a_8685_43396# a_8147_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X4066 C7_P_btm a_n4209_39304# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4067 a_765_45546# a_17609_46634# a_17639_46660# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4068 a_8912_37509# VDAC_N a_5700_37509# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=0.2
X4069 a_11554_42852# a_10796_42968# a_10991_42826# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X4070 a_19386_47436# a_19321_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4071 a_8492_46660# a_7411_46660# a_8145_46902# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X4072 a_2063_45854# a_9863_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4073 VDD a_15803_42450# a_15764_42576# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4074 a_1337_46436# a_1176_45822# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4075 VSS a_949_44458# a_n2438_43548# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4076 VSS a_4419_46090# a_4365_46436# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4077 a_n1549_44318# a_n1899_43946# a_n1644_44306# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4078 VDD a_9067_47204# DATA[4] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4079 VSS a_6575_47204# a_9067_47204# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X4080 a_n1331_43914# a_n1549_44318# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4081 VDD a_3537_45260# a_5093_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1575 pd=1.315 as=0.165 ps=1.33 w=1 l=0.15
X4082 VSS a_11189_46129# a_11608_46482# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X4083 a_20835_44721# a_20640_44752# a_21145_44484# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X4084 w_10694_33990# a_10890_34112# w_10694_33990# w_10694_33990# sky130_fd_pr__pfet_01v8 ad=0.986 pd=7.38 as=0 ps=0 w=3.4 l=16.6
X4085 a_n327_42558# a_n97_42460# a_n473_42460# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.25285 ps=2.52 w=1 l=0.15
X4086 a_8147_43396# a_7499_43078# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X4087 VDD a_n3690_37440# a_n3420_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4088 a_19431_46494# a_18985_46122# a_19335_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4089 VDD a_12607_44458# a_n2661_43922# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4090 VDD a_17324_43396# a_17499_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4091 a_8685_42308# a_8515_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4092 a_1414_42308# a_1067_42314# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X4093 VDD a_4883_46098# a_10355_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4094 a_n2216_37690# a_n2810_45028# a_n2302_37690# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X4095 VDD a_10193_42453# a_9885_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4096 VDD a_21356_42826# a_n357_42282# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4097 a_16977_43638# a_16759_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4098 VSS a_n4334_40480# a_n4064_40160# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X4099 VSS a_n237_47217# a_8270_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4100 a_10555_43940# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4101 a_1049_43396# a_458_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4102 VSS a_22775_42308# a_22485_38105# VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4103 VDD a_n443_42852# a_742_44458# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4104 a_8145_46902# a_7927_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4105 a_21613_42308# a_21335_42336# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X4106 VDD a_n23_45546# a_7_45899# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4107 VSS a_16019_45002# a_15903_45785# VSS sky130_fd_pr__nfet_01v8 ad=0.160875 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X4108 VCM a_5342_30871# C8_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4109 VDD a_2698_46116# a_2804_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X4110 a_20935_43940# a_18479_47436# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4111 a_18194_34908# a_n1794_35082# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4112 a_2713_42308# a_n755_45592# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4113 VDD a_n699_43396# a_4743_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4114 DATA[1] a_1431_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4115 a_17591_47464# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.07035 ps=0.755 w=0.42 l=0.15
X4116 a_9223_42460# a_5891_43370# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X4117 a_12741_44636# a_14537_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4118 a_2684_37794# a_1666_39587# a_1666_39043# VSS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X4119 VDD a_20202_43084# a_21335_42336# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X4120 a_564_42282# a_743_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4121 a_15367_44484# a_13556_45296# a_15004_44636# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4122 VSS a_n2302_40160# a_n4315_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4123 VSS a_n452_47436# a_n815_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4124 VDD a_2063_45854# a_9863_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X4125 a_2981_46116# a_2804_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X4126 VSS a_6511_45714# a_6472_45840# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4127 VSS a_13159_45002# a_13105_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4128 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4129 EN_VIN_BSTR_P a_n1696_34930# w_1575_34786# w_1575_34786# sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X4130 a_9223_42460# a_5891_43370# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X4131 VSS a_19987_42826# a_n2017_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.203125 pd=1.275 as=0.08775 ps=0.92 w=0.65 l=0.15
X4132 a_20692_30879# a_22959_46124# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4133 a_21188_45572# a_20273_45572# a_20841_45814# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4134 a_9028_43914# a_9482_43914# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X4135 VDD a_17715_44484# a_17737_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4136 VSS a_n2840_44458# a_n4318_40392# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4137 VSS a_15004_44636# a_14815_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4138 a_16759_43396# a_16243_43396# a_16664_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4139 a_4574_45260# a_4791_45118# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X4140 a_17829_46910# a_12861_44030# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X4141 VSS a_n443_46116# a_4880_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X4142 a_n4064_38528# a_n4334_38528# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4143 VDD a_1799_45572# a_1983_46706# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X4144 VDD a_21363_45546# a_21350_45938# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4145 SMPL_ON_P a_n2002_35448# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4146 a_n4064_40160# a_n4334_40480# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.138125 ps=1.075 w=0.65 l=0.15
X4147 VDD a_22775_42308# a_22485_38105# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4148 a_13259_45724# a_17583_46090# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4149 w_1575_34786# a_n1057_35014# w_1575_34786# w_1575_34786# sky130_fd_pr__pfet_01v8 ad=0.493 pd=3.69 as=0 ps=0 w=3.4 l=16.6
X4150 VDAC_P a_3422_30871# VCM VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4151 C1_P_btm a_n4064_37440# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4152 VIN_P EN_VIN_BSTR_P C4_P_btm VSS sky130_fd_pr__nfet_01v8 ad=0.31 pd=2.62 as=0.31 ps=2.62 w=1 l=0.15
X4153 a_6575_47204# a_6545_47178# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4154 VSS a_765_45546# a_380_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X4155 VSS a_327_44734# a_501_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4156 a_104_43370# a_n699_43396# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4157 VDD a_22959_42860# a_14097_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4158 a_n2293_42282# a_3357_43084# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4159 VSS a_6171_42473# a_5379_42460# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4160 a_3935_42891# a_2382_45260# a_3935_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4161 VSS a_9067_47204# DATA[4] VSS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X4162 VDD a_8145_46902# a_8035_47026# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X4163 VDD a_n863_45724# a_327_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X4164 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4165 a_17141_43172# a_n1059_45260# a_16795_42852# VSS sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X4166 VDD a_9127_43156# a_5891_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4167 a_15433_44458# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4168 VSS a_10193_42453# a_11897_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X4169 VSS a_4791_45118# a_5066_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4170 VDD a_5691_45260# a_n2109_47186# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.26 ps=2.52 w=1 l=0.15
X4171 VDD a_n1550_35448# a_n2002_35448# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4172 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X4173 VDD a_1983_46706# a_n2661_46098# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4174 a_15227_46910# a_15368_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X4175 a_18753_44484# a_18374_44850# a_18681_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X4176 a_15486_42560# a_15803_42450# a_15761_42308# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X4177 a_n1641_43230# a_n1991_42858# a_n1736_43218# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X4178 a_6682_46987# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X4179 a_n1079_45724# a_n755_45592# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.14575 ps=1.335 w=0.42 l=0.15
X4180 a_12429_44172# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.118125 ps=1.04 w=0.42 l=0.15
X4181 a_1568_43370# a_1847_42826# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4182 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X4183 VSS a_n1794_35082# a_n1696_34930# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4184 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4185 a_10890_34112# a_18194_34908# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=1.24 ps=8.62 w=4 l=0.15
X4186 VDD a_7227_42308# a_6123_31319# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4187 VSS a_1123_46634# a_584_46384# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4188 a_3457_43396# a_3232_43370# a_3626_43646# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X4189 a_7174_31319# a_20107_42308# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4190 a_8952_43230# a_8037_42858# a_8605_42826# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4191 VSS a_167_45260# a_n37_45144# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X4192 a_13490_45067# a_9482_43914# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X4193 a_4181_44734# a_3090_45724# a_n2497_47436# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4194 VSS a_6171_45002# a_11909_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4195 VSS a_n2302_39866# a_n4209_39590# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4196 a_33_46660# a_n133_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4197 a_16388_46812# a_17957_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.112125 ps=0.995 w=0.65 l=0.15
X4198 VDD a_3218_45724# a_3175_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X4199 a_8283_46482# a_n1151_42308# a_7920_46348# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4200 a_8953_45002# CLK VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4201 VSS a_n809_44244# a_n755_45592# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4202 VDD a_15279_43071# a_14579_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4203 VDD a_16763_47508# a_5807_45002# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4204 VDD a_310_45028# a_509_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X4205 a_n23_47502# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4206 a_n1099_45572# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1925 ps=1.385 w=1 l=0.15
X4207 VDD a_10903_43370# a_10907_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.635 ps=3.27 w=1 l=0.15
X4208 a_3935_43218# a_3681_42891# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1449 ps=1.11 w=0.42 l=0.15
X4209 a_14949_46494# a_13759_46122# a_14840_46494# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X4210 a_11599_46634# a_15682_46116# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4211 a_6851_47204# a_6491_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4212 a_13556_45296# a_6755_46942# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4213 VDD a_n4315_30879# a_n4334_40480# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X4214 VSS a_15227_44166# a_14539_43914# VSS sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.08775 ps=0.92 w=0.65 l=0.15
X4215 a_19987_42826# a_18494_42460# a_20356_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
X4216 a_n2833_47464# a_n2497_47436# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.165 ps=1.33 w=1 l=0.15
X4217 a_3524_46660# a_2609_46660# a_3177_46902# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X4218 a_n4209_39304# a_n2302_39072# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.115375 ps=1.005 w=0.65 l=0.15
X4219 VSS a_22223_47212# a_21588_30879# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4220 VSS a_6151_47436# a_6229_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X4221 a_18533_43940# a_13661_43548# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X4222 a_14205_43396# a_13667_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X4223 VREF a_n3565_39590# C8_P_btm VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4224 VCM a_3422_30871# VDAC_N VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4225 VDD a_949_44458# a_n2438_43548# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4226 a_n4064_37440# a_n4334_37440# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4227 a_16377_45572# a_16333_45814# a_16211_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X4228 a_4646_46812# a_6298_44484# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X4229 a_10044_46482# a_n743_46660# a_9823_46155# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4230 a_19113_45348# a_18911_45144# a_3090_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4231 VSS a_13720_44458# a_12607_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X4232 a_n2860_37984# a_n2956_38216# a_n2946_37984# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X4233 a_2266_47570# a_n971_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4234 a_5837_43396# a_5111_44636# a_5147_45002# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4235 a_5934_30871# a_8791_42308# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X4236 a_10861_46660# a_10227_46804# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X4237 VSS a_7920_46348# a_7715_46873# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4238 a_14383_46116# a_10227_46804# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X4239 a_2809_45348# a_526_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4240 a_2905_42968# a_742_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4241 a_6540_46812# a_6755_46942# a_6682_46987# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X4242 a_6709_45028# a_6431_45366# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X4243 a_8953_45002# CLK VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4244 VSS a_18494_42460# a_20193_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4245 a_n2442_46660# a_n2472_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4246 C7_P_btm EN_VIN_BSTR_P VIN_P VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X4247 a_13249_42308# a_13070_42354# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X4248 a_n1991_42858# a_n2157_42858# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4249 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X4250 VDD a_15682_46116# a_11599_46634# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4251 a_13348_45260# a_12891_46348# a_13490_45067# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X4252 VREF_GND a_n4064_39616# C9_P_btm VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4253 a_17061_44484# a_11691_44458# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X4254 comp_n a_1169_39043# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4255 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X4256 VDD a_18443_44721# a_18374_44850# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X4257 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4258 a_1512_43396# a_n443_46116# a_1209_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X4259 VDD a_n3565_39304# a_n3690_39392# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.14 ps=1.28 w=1 l=0.15
X4260 VDD a_22591_44484# a_17730_32519# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4261 VDD a_22581_37893# a_22537_39537# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4262 VDD a_n2002_35448# SMPL_ON_P VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4263 VSS a_15803_42450# a_15764_42576# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4264 a_11901_46660# a_11735_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4265 a_21076_30879# a_22959_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4266 a_3877_44458# a_3699_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X4267 VDD a_n4064_39072# a_n2216_39072# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1775 pd=1.355 as=0.105 ps=1.21 w=1 l=0.15
X4268 a_11599_46634# a_15682_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4269 a_11691_44458# a_5807_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4270 a_15368_46634# a_15143_45578# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X4271 VSS a_9028_43914# a_8975_43940# VSS sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X4272 a_2813_43396# a_n443_46116# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.12675 ps=1.04 w=0.65 l=0.15
X4273 C8_N_btm a_17538_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4274 a_5093_45028# a_4558_45348# a_5009_45028# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4275 VSS a_10193_42453# a_13921_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X4276 a_15597_42852# a_15567_42826# a_15095_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X4277 a_2553_47502# a_n971_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4278 VDD a_13059_46348# a_12839_46116# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4279 C10_N_btm a_22612_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4280 a_3823_42558# a_3065_45002# a_3905_42308# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X4281 VDD a_526_44458# a_5193_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4282 VSS a_1667_45002# a_n863_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X4283 a_1307_43914# a_2779_44458# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4284 VDD a_n3690_38528# a_n3420_38528# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X4285 VDD a_21177_47436# a_20990_47178# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X4286 a_16855_45546# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4287 a_5495_43940# a_5244_44056# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X4288 VDD a_5815_47464# a_n1613_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.14 ps=1.28 w=1 l=0.15
X4289 VSS a_19787_47423# a_19594_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4290 VDD a_22365_46825# a_20202_43084# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4291 a_5063_47570# a_4915_47217# a_4700_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4292 a_n1736_46482# a_n1853_46287# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4293 VDD a_11459_47204# DATA[5] VDD sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X4294 a_11322_45546# a_11823_42460# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4295 a_19787_47423# START VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4296 a_3754_39466# a_7754_39632# VSS sky130_fd_pr__res_high_po_0p35 l=18
X4297 a_n4251_39616# a_n4318_39768# a_n4334_39616# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.17225 ps=1.83 w=0.65 l=0.15
X4298 VDD a_9127_43156# a_9114_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4299 a_10384_47026# a_9863_46634# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4300 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X4301 VSS a_11525_45546# a_11189_46129# VSS sky130_fd_pr__nfet_01v8 ad=0.167375 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X4302 SMPL_ON_N a_21753_35474# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4303 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X4304 a_10729_43914# a_11750_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4305 a_4921_42308# a_n913_45002# a_4933_42558# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4306 VSS a_n23_47502# a_n89_47570# VSS sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4307 a_20528_46660# a_20411_46873# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X4308 VSS a_8568_45546# a_8162_45546# VSS sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X4309 a_13657_42558# a_13259_45724# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X4310 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X4311 VSS a_4223_44672# a_5205_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4312 a_18005_44484# a_17970_44736# a_17767_44458# VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X4313 a_13837_43396# a_13259_45724# a_13749_43396# VSS sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X4314 a_19177_43646# a_17339_46660# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X4315 a_196_42282# a_375_42282# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4316 a_791_42968# a_n1059_45260# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4317 VSS a_327_47204# DATA[0] VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4318 a_11309_47204# a_11031_47542# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X4319 VSS a_4646_46812# a_7871_42858# VSS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4320 VSS a_5815_47464# a_n1613_43370# VSS sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.0588 ps=0.7 w=0.42 l=0.15
X4321 a_n23_45546# a_n356_45724# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X4322 a_18691_45572# a_18175_45572# a_18596_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X4323 a_9885_42558# a_9290_44172# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X4324 VSS a_4700_47436# a_3785_47178# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4325 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X4326 a_4361_42308# a_3823_42558# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X4327 VDD a_n2840_46634# a_n2956_39768# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X4328 a_4817_46660# a_4651_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4329 VDD a_13635_43156# a_13622_42852# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X4330 VDD a_n2438_43548# a_n2157_42858# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4331 a_8415_44056# a_5343_44458# a_8333_44056# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X4332 a_8912_37509# VDAC_P a_5088_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.2
X4333 VSS a_1307_43914# a_4156_43218# VSS sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.0693 ps=0.75 w=0.42 l=0.15
X4334 a_n1699_44726# a_n1917_44484# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X4335 a_1525_44260# a_1467_44172# a_1115_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X4336 VDD a_n2946_39866# a_n3565_39590# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4337 a_14976_45028# a_14797_45144# a_15060_45348# VSS sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.125125 ps=1.035 w=0.65 l=0.15
X4338 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X4339 a_2324_44458# a_8953_45002# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4340 VSS VDD VSS VSS sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X4341 a_n3565_39304# a_n2946_39072# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1775 ps=1.355 w=1 l=0.15
X4342 VSS a_15959_42545# a_15890_42674# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X4343 a_n2312_39304# a_n1920_47178# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X4344 VDD a_15682_43940# a_11967_42832# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4345 VIN_N EN_VIN_BSTR_N C7_N_btm VSS sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X4346 VDD a_1666_39587# a_1666_39043# VDD sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X4347 VDD a_n3690_37440# a_n3420_37440# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.285 pd=2.57 as=0.14 ps=1.28 w=1 l=0.15
X4348 VSS a_21363_45546# a_21297_45572# VSS sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X4349 VDD a_n452_44636# a_n2129_44697# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X4350 a_19443_46116# a_18819_46122# a_19335_46494# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4351 VDD a_7112_43396# a_7287_43370# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X4352 a_310_45028# a_n37_45144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X4353 VDD a_5111_44636# a_5518_44484# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.3 ps=2.6 w=1 l=0.15
X4354 a_17719_45144# a_17613_45144# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X4355 a_17499_43370# a_16327_47482# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X4356 VDD a_12563_42308# a_5534_30871# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X4357 VSS a_13747_46662# a_19466_46812# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4358 a_14112_44734# a_768_44030# a_13857_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X4359 VSS a_n2946_38778# a_n3565_38502# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4360 a_n357_42282# a_21356_42826# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4361 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X4362 VDD a_3483_46348# a_15037_43940# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X4363 VCM a_4190_30871# C10_P_btm VSS sky130_fd_pr__nfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4364 a_5700_37509# VDAC_N a_8912_37509# VDD sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=0.2
X4365 VDD a_13635_43156# a_9290_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=2.61 as=0.135 ps=1.27 w=1 l=0.15
X4366 VDD a_13487_47204# a_768_44030# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4367 a_14097_32519# a_22959_42860# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4368 a_3094_47570# a_2905_45572# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4369 a_8270_45546# a_n237_47217# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4370 a_8781_46436# a_8199_44636# a_8034_45724# VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4371 VDD VSS VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X4372 VSS a_3232_43370# a_11541_44484# VSS sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X4373 DATA[4] a_9067_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X4374 a_20841_46902# a_20623_46660# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4375 a_13527_45546# a_12861_44030# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4376 a_10533_42308# a_7499_43078# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4377 a_17896_45144# a_16922_45042# a_17801_45144# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
X4378 DATA[1] a_1431_47204# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X4379 a_18817_42826# a_18599_43230# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X4380 a_104_43370# a_n699_43396# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X4381 C10_P_btm a_n4315_30879# VREF VDD sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=0.35
X4382 a_16211_45572# a_15765_45572# a_16115_45572# VSS sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X4383 VDD a_4223_44672# a_4181_44734# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X4384 VSS a_20835_44721# a_20766_44850# VSS sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X4385 a_19741_43940# a_19478_44306# a_19328_44172# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4386 VDD a_13747_46662# a_14495_45572# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X4387 a_2487_47570# a_2063_45854# a_2124_47436# VSS sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4388 VSS a_10809_44734# a_22959_46124# VSS sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4389 a_11967_42832# a_15682_43940# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4390 C10_N_btm a_18114_32519# VREF_GND VSS sky130_fd_pr__nfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4391 VSS a_7754_38470# a_6886_37412# VSS sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.62 ps=4.62 w=2 l=0.15
X4392 VSS a_20567_45036# a_12549_44172# VSS sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4393 a_21359_45002# a_21513_45002# VDD VDD sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X4394 a_18451_43940# a_18579_44172# a_18533_44260# VSS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X4395 a_13904_45546# a_13249_42308# a_14033_45822# VDD sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X4396 VSS a_13661_43548# a_18587_45118# VSS sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X4397 a_6547_43396# a_6031_43396# a_6452_43396# VSS sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
C0 a_n237_47217# a_5257_43370# 0.022234f
C1 a_n1151_42308# a_4955_46873# 0.261025f
C2 a_n971_45724# a_7715_46873# 0.029319f
C3 a_n4318_37592# a_n4064_37440# 0.04779f
C4 a_13258_32519# a_7174_31319# 0.02542f
C5 a_16327_47482# a_18083_42858# 0.591108f
C6 a_21588_30879# a_13467_32519# 0.057457f
C7 a_8199_44636# a_9672_43914# 0.043804f
C8 a_3537_45260# a_4574_45260# 0.234297f
C9 a_11453_44696# a_3483_46348# 0.027804f
C10 a_768_44030# a_11415_45002# 0.021062f
C11 a_4883_46098# a_5164_46348# 0.01685f
C12 a_4646_46812# a_3090_45724# 0.199722f
C13 a_n1613_43370# a_n1853_46287# 0.354256f
C14 a_11599_46634# a_13351_46090# 0.105205f
C15 a_n4209_39590# VIN_P 0.10512f
C16 a_n4064_40160# VCM 0.121302f
C17 a_7754_38636# a_5088_37509# 0.288061f
C18 VDAC_Ni a_4338_37500# 0.640521f
C19 a_n4209_37414# a_n2302_37690# 0.407594f
C20 a_n3565_37414# a_n2946_37690# 0.407439f
C21 a_n3690_37440# a_n3420_37440# 0.431074f
C22 a_n4334_37440# a_n4064_37440# 0.448688f
C23 a_16019_45002# VDD 0.174085f
C24 a_n97_42460# a_19339_43156# 0.012502f
C25 a_n2661_42282# a_n3674_37592# 0.12829f
C26 a_7229_43940# a_n2661_43922# 0.030151f
C27 a_4185_45028# a_14209_32519# 0.091175f
C28 a_8199_44636# a_743_42282# 0.036554f
C29 a_n2017_45002# a_11967_42832# 0.086561f
C30 a_9482_43914# a_9313_44734# 0.060868f
C31 a_4791_45118# a_5932_42308# 0.212275f
C32 a_n743_46660# a_n23_45546# 0.070296f
C33 a_15227_44166# a_6945_45028# 0.548194f
C34 a_17609_46634# a_10809_44734# 0.018125f
C35 a_12861_44030# a_15765_45572# 0.026773f
C36 a_n2293_46098# a_n1853_46287# 0.02738f
C37 a_17364_32525# a_14097_32519# 0.059348f
C38 a_2982_43646# a_17303_42282# 0.139588f
C39 a_4223_44672# a_6453_43914# 0.019918f
C40 a_2437_43646# a_2813_43396# 0.012852f
C41 a_n1613_43370# a_n2661_43370# 0.05744f
C42 a_1823_45246# a_3775_45552# 0.070347f
C43 a_11415_45002# a_11652_45724# 0.128811f
C44 a_11453_44696# a_17719_45144# 0.105851f
C45 a_8953_45546# a_n443_42852# 0.134632f
C46 a_3877_44458# a_2382_45260# 0.395451f
C47 a_3090_45724# a_18479_45785# 0.259218f
C48 a_18479_47436# a_20193_45348# 0.021013f
C49 a_4185_45028# a_4099_45572# 0.025863f
C50 a_8791_43396# VDD 0.191045f
C51 a_4190_30871# a_n3420_37440# 0.034998f
C52 a_n2293_42282# a_1606_42308# 0.192228f
C53 a_20193_45348# a_4190_30871# 0.02125f
C54 a_10428_46928# VDD 0.278873f
C55 a_n755_45592# a_1606_42308# 0.104938f
C56 a_8049_45260# a_2437_43646# 0.041161f
C57 a_n2293_46098# a_n2661_43370# 0.027372f
C58 a_2324_44458# a_8953_45002# 1.65784f
C59 a_3090_45724# a_10057_43914# 0.230475f
C60 a_10227_46804# a_10405_44172# 0.011223f
C61 a_10227_46804# a_19386_47436# 0.041193f
C62 a_18479_47436# a_18780_47178# 0.056304f
C63 a_n237_47217# a_5807_45002# 0.082779f
C64 a_n443_46116# a_n881_46662# 0.114922f
C65 a_4915_47217# a_n1613_43370# 0.195064f
C66 a_16327_47482# a_13507_46334# 0.043159f
C67 a_n4318_37592# a_n3420_39072# 0.02033f
C68 a_n3674_38216# a_n4064_39072# 0.019725f
C69 a_15493_43396# a_19268_43646# 0.024436f
C70 a_4185_45028# a_17730_32519# 0.097949f
C71 a_n357_42282# a_n2661_44458# 0.031616f
C72 a_3090_45724# a_14021_43940# 0.049176f
C73 a_12549_44172# a_10341_43396# 0.0385f
C74 a_21513_45002# a_3357_43084# 0.04265f
C75 a_5807_45002# a_8270_45546# 0.029164f
C76 a_12891_46348# a_12816_46660# 0.024711f
C77 a_12549_44172# a_12991_46634# 0.010497f
C78 a_12861_44030# a_18280_46660# 0.140921f
C79 a_n2661_46634# a_6755_46942# 1.40968f
C80 a_n237_47217# a_3699_46348# 0.044064f
C81 a_4883_46098# a_16388_46812# 0.041939f
C82 a_584_46384# a_1823_45246# 0.094654f
C83 a_14456_42282# VDD 0.265543f
C84 a_22485_38105# a_22581_37893# 0.902394f
C85 a_19237_31679# a_14097_32519# 0.052198f
C86 a_3537_45260# a_5883_43914# 0.018824f
C87 a_5111_44636# a_5518_44484# 0.124556f
C88 SMPL_ON_P a_n3674_38680# 0.038963f
C89 a_3232_43370# a_n699_43396# 0.074855f
C90 a_768_44030# a_13259_45724# 0.315247f
C91 a_2063_45854# a_11962_45724# 0.011034f
C92 a_n2661_46634# a_8049_45260# 0.027919f
C93 C4_N_btm VDD 0.265463f
C94 C9_P_btm VREF_GND 5.18245f
C95 C10_P_btm VCM 10.5945f
C96 C8_P_btm VREF 3.6701f
C97 C6_N_btm C10_N_btm 0.895671f
C98 C7_N_btm C9_N_btm 0.22201f
C99 C6_P_btm VIN_P 0.391898f
C100 a_11827_44484# a_3422_30871# 0.076229f
C101 a_1307_43914# a_10405_44172# 0.010378f
C102 a_13076_44458# a_13213_44734# 0.126609f
C103 a_11823_42460# a_14205_43396# 0.176571f
C104 a_12465_44636# a_9482_43914# 0.069673f
C105 a_8199_44636# a_8049_45260# 0.069189f
C106 a_22612_30879# a_19963_31679# 0.078731f
C107 a_4791_45118# a_n2661_43370# 0.408007f
C108 a_21588_30879# RST_Z 0.052092f
C109 a_11967_42832# a_18079_43940# 0.052453f
C110 a_2675_43914# a_2998_44172# 0.173844f
C111 a_n913_45002# a_8952_43230# 0.04786f
C112 a_22612_30879# VDD 3.23752f
C113 a_9290_44172# a_13070_42354# 0.140007f
C114 a_2957_45546# a_2711_45572# 0.056166f
C115 a_12741_44636# a_6171_45002# 0.08387f
C116 a_n2438_43548# a_n356_44636# 0.082195f
C117 a_768_44030# a_n2661_43922# 1.9176f
C118 a_12891_46348# a_13213_44734# 0.052195f
C119 a_12549_44172# a_n2293_43922# 0.194293f
C120 a_5342_30871# C6_N_btm 0.012f
C121 a_4791_45118# a_4915_47217# 0.226891f
C122 a_2063_45854# a_9863_47436# 0.12173f
C123 a_12895_43230# VDD 0.212352f
C124 a_5755_42308# a_6171_42473# 0.017801f
C125 a_7920_46348# VDD 0.100184f
C126 a_2711_45572# a_9482_43914# 0.01017f
C127 a_1138_42852# a_n2661_42834# 0.024191f
C128 a_13249_42308# a_n913_45002# 0.019571f
C129 a_12741_44636# a_14673_44172# 0.178572f
C130 a_11459_47204# a_11735_46660# 0.010464f
C131 a_n2661_46634# a_n2442_46660# 0.063483f
C132 a_n3674_38216# VDD 0.309006f
C133 a_n3565_39590# a_n4209_38502# 0.0315f
C134 a_n4209_39304# a_n3690_39392# 0.045342f
C135 a_n4209_39590# a_n3565_38502# 0.031792f
C136 a_n4064_40160# a_n4064_38528# 0.055466f
C137 a_6171_45002# a_n2293_42834# 0.035829f
C138 a_9290_44172# a_9801_43940# 0.091547f
C139 a_4185_45028# a_17538_32519# 0.043989f
C140 a_n237_47217# a_n755_45592# 0.286948f
C141 a_584_46384# a_n2293_45546# 0.029113f
C142 a_2107_46812# a_3147_46376# 0.010901f
C143 a_n2661_46098# a_1208_46090# 0.023477f
C144 a_5807_45002# a_13759_46122# 0.022269f
C145 a_8530_39574# VDD 0.346613f
C146 a_22629_37990# a_22737_36887# 0.08947f
C147 VDAC_P C5_P_btm 27.6071f
C148 a_7754_38470# RST_Z 0.034995f
C149 a_11827_44484# VDD 0.615802f
C150 a_3065_45002# a_3600_43914# 0.011102f
C151 a_n2312_38680# a_n3674_38216# 0.023419f
C152 a_n2442_46660# COMP_P 0.024155f
C153 a_10227_46804# a_15486_42560# 0.227612f
C154 a_10227_46804# a_3357_43084# 0.305304f
C155 a_8199_44636# a_8953_45546# 0.71291f
C156 a_8016_46348# a_9569_46155# 0.044705f
C157 a_n2840_46090# a_n2956_39304# 0.158668f
C158 a_4791_45118# a_4574_45260# 0.091783f
C159 a_5649_42852# a_5742_30871# 0.059614f
C160 a_18287_44626# a_19328_44172# 0.011011f
C161 a_n2661_42834# a_n4318_39768# 0.031793f
C162 a_16588_47582# VDD 0.282243f
C163 a_n1613_43370# a_5883_43914# 0.352323f
C164 a_3090_45724# a_4927_45028# 0.088804f
C165 a_n3674_38680# a_n1794_35082# 0.020981f
C166 a_n4318_38216# a_n3674_37592# 0.077253f
C167 a_10405_44172# a_10867_43940# 0.022925f
C168 a_n913_45002# a_22223_42860# 0.011179f
C169 a_n2017_45002# a_n2293_42282# 0.095773f
C170 a_12741_44636# a_12607_44458# 0.134974f
C171 a_n755_45592# a_n2017_45002# 0.088948f
C172 a_n357_42282# a_n1059_45260# 7.3759f
C173 a_1609_45822# a_2437_43646# 0.189329f
C174 a_n443_46116# a_1049_43396# 0.085877f
C175 a_n2293_46098# a_5883_43914# 0.069185f
C176 a_16375_45002# a_6171_45002# 0.026914f
C177 a_13661_43548# a_17973_43940# 0.031319f
C178 a_12549_44172# a_21115_43940# 0.211261f
C179 a_16327_47482# a_n743_46660# 0.53683f
C180 a_10227_46804# a_n2293_46634# 0.032913f
C181 a_n971_45724# a_7411_46660# 0.567031f
C182 a_12465_44636# a_13747_46662# 0.039773f
C183 a_n1613_43370# a_n881_46662# 1.06426f
C184 a_4883_46098# a_19321_45002# 0.026904f
C185 a_n1151_42308# a_4651_46660# 0.028941f
C186 a_19511_42282# a_21335_42336# 0.011904f
C187 a_13258_32519# a_20712_42282# 0.016015f
C188 a_6547_43396# a_6643_43396# 0.013793f
C189 a_13259_45724# a_17517_44484# 0.028602f
C190 a_8016_46348# a_10405_44172# 0.098226f
C191 a_3357_43084# a_1307_43914# 0.197864f
C192 a_10227_46804# a_5342_30871# 0.163388f
C193 a_12549_44172# a_11415_45002# 0.028008f
C194 a_4883_46098# a_5068_46348# 0.031466f
C195 a_7927_46660# a_8035_47026# 0.057222f
C196 a_3877_44458# a_3090_45724# 0.23348f
C197 a_11599_46634# a_12594_46348# 0.085826f
C198 a_n1613_43370# a_n2157_46122# 0.296124f
C199 a_4915_47217# a_6945_45028# 0.207881f
C200 a_n881_46662# a_n2293_46098# 0.291354f
C201 a_10554_47026# a_10249_46116# 0.023301f
C202 a_n4064_40160# VREF_GND 0.493568f
C203 VDAC_Ni a_3726_37500# 1.5261f
C204 a_n3565_37414# a_n3420_37440# 0.307576f
C205 a_n4209_37414# a_n4064_37440# 0.265895f
C206 a_4190_30871# a_5534_30871# 0.020828f
C207 a_16823_43084# a_16795_42852# 0.065873f
C208 a_15595_45028# VDD 0.156299f
C209 a_7229_43940# a_n2661_42834# 0.023622f
C210 a_7499_43078# a_10555_44260# 0.03816f
C211 a_n2661_45546# a_n97_42460# 0.038952f
C212 SMPL_ON_N a_14097_32519# 0.029158f
C213 a_n743_46660# a_n356_45724# 0.223429f
C214 a_13747_46662# a_2711_45572# 0.032065f
C215 a_15227_44166# a_21137_46414# 0.081665f
C216 a_n2293_46098# a_n2157_46122# 0.015455f
C217 a_12861_44030# a_15903_45785# 0.156145f
C218 a_11453_44696# a_13249_42308# 0.026348f
C219 a_13059_46348# a_10903_43370# 0.11738f
C220 a_n2661_46098# a_n2661_45546# 0.011799f
C221 a_2982_43646# a_4958_30871# 0.136637f
C222 a_4223_44672# a_5663_43940# 0.01368f
C223 a_2324_44458# a_n863_45724# 0.01106f
C224 a_4419_46090# a_2711_45572# 0.026096f
C225 a_n2293_46634# a_1307_43914# 0.184387f
C226 a_3090_45724# a_18175_45572# 0.130163f
C227 a_8147_43396# VDD 0.393534f
C228 a_10150_46912# VDD 0.284144f
C229 a_18184_42460# a_5649_42852# 0.028842f
C230 a_19279_43940# a_19319_43548# 0.023499f
C231 a_2324_44458# a_8191_45002# 0.120399f
C232 a_12861_44030# a_11453_44696# 0.173308f
C233 a_10227_46804# a_18597_46090# 0.07604f
C234 a_n2833_47464# a_n2840_46634# 0.019713f
C235 a_2063_45854# a_768_44030# 0.027746f
C236 a_4791_45118# a_n881_46662# 0.429542f
C237 a_n443_46116# a_n1613_43370# 0.410263f
C238 a_11599_46634# a_12465_44636# 0.018625f
C239 a_n97_42460# a_1427_43646# 0.047018f
C240 a_15493_43396# a_15743_43084# 0.517624f
C241 a_10227_46804# a_743_42282# 0.045325f
C242 a_4185_45028# a_22591_44484# 0.013394f
C243 a_16327_47482# a_4361_42308# 0.029635f
C244 a_13259_45724# a_13720_44458# 0.016851f
C245 a_n2293_46634# a_9396_43370# 0.012588f
C246 a_2437_43646# a_22223_45572# 0.165664f
C247 a_12891_46348# a_12991_46634# 0.018656f
C248 a_584_46384# a_1138_42852# 0.491749f
C249 a_n1151_42308# a_n1076_46494# 0.023834f
C250 a_12861_44030# a_17639_46660# 0.033515f
C251 a_3699_46634# a_3877_44458# 0.087244f
C252 a_n2661_46634# a_10249_46116# 0.055133f
C253 a_n237_47217# a_3483_46348# 0.090759f
C254 a_4883_46098# a_13059_46348# 0.097406f
C255 a_18597_46090# a_17339_46660# 0.018491f
C256 a_n443_46116# a_n2293_46098# 0.251135f
C257 a_n4209_39304# a_n3420_37440# 0.033347f
C258 a_13575_42558# VDD 0.182133f
C259 a_n3565_39304# a_n3565_37414# 0.029571f
C260 a_n3420_39072# a_n4209_37414# 0.030579f
C261 a_n4064_37984# a_n2302_37984# 0.250408f
C262 a_19963_31679# C3_N_btm 0.041776f
C263 a_5111_44636# a_5343_44458# 0.477401f
C264 a_5147_45002# a_5518_44484# 0.064422f
C265 a_1307_43914# a_16237_45028# 0.056593f
C266 a_3232_43370# a_4223_44672# 0.033907f
C267 a_12549_44172# a_13259_45724# 0.110646f
C268 a_8270_45546# a_3483_46348# 0.058754f
C269 a_n1151_42308# a_10193_42453# 0.238612f
C270 a_11599_46634# a_2711_45572# 0.018466f
C271 C3_N_btm VDD 0.26836f
C272 C10_P_btm VREF_GND 10.3207f
C273 C9_P_btm VREF 7.369471f
C274 C5_N_btm C10_N_btm 0.51798f
C275 C6_N_btm C9_N_btm 0.165353f
C276 C7_N_btm C8_N_btm 31.072699f
C277 C7_P_btm VIN_P 1.52449f
C278 a_22959_43396# a_22959_42860# 0.026152f
C279 a_11823_42460# a_14358_43442# 0.122636f
C280 a_13249_42308# a_9145_43396# 0.072489f
C281 a_13556_45296# a_14955_43940# 0.059957f
C282 a_6945_45028# a_10809_44734# 0.953135f
C283 a_765_45546# a_1609_45822# 0.021736f
C284 a_21076_30879# a_20692_30879# 0.117886f
C285 a_21588_30879# a_19963_31679# 0.055898f
C286 a_n1613_43370# a_3537_45260# 0.095192f
C287 a_11967_42832# a_17973_43940# 0.070514f
C288 a_2675_43914# a_2889_44172# 0.083573f
C289 a_n1899_43946# a_n1644_44306# 0.06121f
C290 a_n913_45002# a_9127_43156# 0.038139f
C291 a_n1059_45260# a_8952_43230# 0.010945f
C292 a_21588_30879# VDD 1.79397f
C293 a_9290_44172# a_12563_42308# 0.052279f
C294 a_n2293_46098# a_3537_45260# 0.019207f
C295 a_n443_46116# a_2675_43914# 0.011921f
C296 a_768_44030# a_n2661_42834# 4.99505f
C297 a_12549_44172# a_n2661_43922# 0.061277f
C298 a_5534_30871# C7_N_btm 0.060228f
C299 a_4791_45118# a_n443_46116# 0.115639f
C300 a_4700_47436# a_4915_47217# 0.07122f
C301 a_13113_42826# VDD 0.217254f
C302 a_9313_44734# a_10835_43094# 0.050385f
C303 a_n356_44636# a_17701_42308# 0.065679f
C304 a_6419_46155# VDD 0.094119f
C305 a_10193_42453# a_18214_42558# 0.028997f
C306 a_20202_43084# a_17517_44484# 0.021286f
C307 a_7227_45028# a_6709_45028# 0.115677f
C308 a_13249_42308# a_n1059_45260# 0.026496f
C309 a_4185_45028# a_9313_44734# 0.078424f
C310 a_n443_42852# a_375_42282# 0.075658f
C311 a_10227_46804# a_6755_46942# 0.778648f
C312 a_n2661_46634# a_n2472_46634# 0.0842f
C313 a_n2956_39768# a_n2442_46660# 6.5214f
C314 a_n2104_42282# VDD 0.280329f
C315 a_n4209_39304# a_n3565_39304# 6.82668f
C316 a_10341_43396# a_16409_43396# 0.028466f
C317 a_10907_45822# VDD 0.352181f
C318 a_4185_45028# a_20974_43370# 0.184625f
C319 a_3232_43370# a_n2293_42834# 0.041207f
C320 a_19479_31679# a_22959_45036# 0.018372f
C321 a_3065_45002# a_n2661_43370# 0.356646f
C322 a_n881_46662# a_6945_45028# 0.239384f
C323 a_n746_45260# a_n755_45592# 0.172774f
C324 a_n743_46660# a_5204_45822# 0.034798f
C325 a_n2661_46098# a_805_46414# 0.044109f
C326 a_10227_46804# a_8049_45260# 0.058336f
C327 a_7754_38470# VDD 0.302129f
C328 VDAC_P C6_P_btm 55.214397f
C329 a_14543_43071# a_5534_30871# 0.196814f
C330 a_21359_45002# VDD 0.319372f
C331 a_n97_42460# a_16877_42852# 0.011527f
C332 a_n2442_46660# a_n4318_37592# 0.023729f
C333 a_2382_45260# a_3905_42865# 0.291572f
C334 a_9290_44172# a_12089_42308# 0.047614f
C335 a_10227_46804# a_15051_42282# 0.361922f
C336 a_3065_45002# a_2998_44172# 0.024536f
C337 a_18479_47436# a_2437_43646# 0.041425f
C338 a_8016_46348# a_9625_46129# 0.128435f
C339 a_8199_44636# a_5937_45572# 0.573373f
C340 a_13747_46662# a_14033_45822# 0.021007f
C341 a_17339_46660# a_8049_45260# 0.023006f
C342 a_4791_45118# a_3537_45260# 0.33264f
C343 a_5534_30871# COMP_P 0.027557f
C344 a_16137_43396# a_18214_42558# 0.0459f
C345 a_n2661_42282# VDD 0.406474f
C346 a_n2293_42834# a_4905_42826# 0.046599f
C347 a_19279_43940# a_3422_30871# 0.02352f
C348 a_13717_47436# CLK 0.057477f
C349 a_16763_47508# VDD 0.392885f
C350 a_3090_45724# a_5111_44636# 0.063636f
C351 a_2324_44458# a_11823_42460# 0.058835f
C352 a_6755_46942# a_1307_43914# 0.076439f
C353 a_16823_43084# VDD 0.159922f
C354 a_13467_32519# C1_N_btm 0.031032f
C355 COMP_P a_n1329_42308# 0.232443f
C356 a_n2840_42282# a_n1794_35082# 0.040623f
C357 a_n356_44636# a_4361_42308# 0.030056f
C358 a_10405_44172# a_10651_43940# 0.014272f
C359 a_n913_45002# a_22165_42308# 0.074472f
C360 a_n357_42282# a_n2017_45002# 0.580077f
C361 a_n2293_45546# a_n967_45348# 0.119714f
C362 a_n443_46116# a_1209_43370# 0.061682f
C363 a_4185_45028# a_18114_32519# 0.080343f
C364 a_13661_43548# a_17737_43940# 0.031811f
C365 a_12549_44172# a_20935_43940# 0.110704f
C366 a_n1151_42308# a_4646_46812# 0.330834f
C367 a_12465_44636# a_13661_43548# 0.106973f
C368 a_13258_32519# a_20107_42308# 0.021019f
C369 a_19511_42282# a_7174_31319# 0.240861f
C370 a_n2956_37592# a_n4064_40160# 0.012264f
C371 a_n1613_43370# a_n1533_42852# 0.012196f
C372 a_n2661_45546# a_n2661_43922# 0.028803f
C373 a_3429_45260# a_3537_45260# 0.138977f
C374 a_8016_46348# a_9672_43914# 0.074243f
C375 a_12861_44030# a_13925_46122# 0.012485f
C376 a_11599_46634# a_12005_46116# 0.27095f
C377 a_12891_46348# a_11415_45002# 0.059955f
C378 a_12549_44172# a_20202_43084# 0.028142f
C379 a_8145_46902# a_8035_47026# 0.097745f
C380 a_7927_46660# a_7832_46660# 0.049827f
C381 a_n743_46660# a_16721_46634# 0.038286f
C382 a_n1613_43370# a_n2293_46098# 0.037934f
C383 a_10623_46897# a_10249_46116# 0.032312f
C384 a_10467_46802# a_6755_46942# 0.256039f
C385 a_4883_46098# a_4704_46090# 0.1774f
C386 a_n4209_38502# C5_P_btm 0.040445f
C387 a_n4315_30879# VCM 0.473529f
C388 a_1666_39587# VDD 3.12922f
C389 a_n3565_37414# a_n3690_37440# 0.247968f
C390 a_n4334_37440# a_n3420_37440# 0.015567f
C391 a_n4209_37414# a_n2946_37690# 0.023544f
C392 a_16823_43084# a_16414_43172# 0.024882f
C393 a_n2661_42282# a_n784_42308# 0.062364f
C394 a_15415_45028# VDD 0.191729f
C395 a_5205_44484# a_n2661_43922# 0.032439f
C396 a_4185_45028# a_13887_32519# 0.044689f
C397 a_10193_42453# a_15493_43940# 0.597095f
C398 a_13661_43548# a_2711_45572# 0.552383f
C399 a_15227_44166# a_20708_46348# 0.106656f
C400 a_n2472_46090# a_n2157_46122# 0.080495f
C401 a_12861_44030# a_15599_45572# 0.025507f
C402 a_14209_32519# a_14097_32519# 10.7606f
C403 a_8387_43230# a_8495_42852# 0.057222f
C404 a_4190_30871# COMP_P 0.027242f
C405 a_19279_43940# VDD 0.302681f
C406 a_9313_44734# a_11967_42832# 0.216837f
C407 a_4223_44672# a_5495_43940# 0.06577f
C408 en_comp a_2982_43646# 0.021697f
C409 a_4185_45028# a_2711_45572# 0.102913f
C410 a_4791_45118# a_8701_44490# 0.138973f
C411 a_8034_45724# a_8049_45260# 0.141057f
C412 a_8199_44636# a_n443_42852# 0.021145f
C413 a_13507_46334# a_18494_42460# 0.234442f
C414 a_11415_45002# a_11322_45546# 0.527707f
C415 a_3090_45724# a_16147_45260# 0.076341f
C416 a_12741_44636# a_10193_42453# 0.078619f
C417 a_3483_46348# a_4099_45572# 0.15767f
C418 a_7112_43396# VDD 0.273193f
C419 a_n2293_42834# a_2905_42968# 0.010834f
C420 a_9863_46634# VDD 0.411318f
C421 a_16922_45042# a_20749_43396# 0.106779f
C422 a_18184_42460# a_13678_32519# 0.019189f
C423 a_8953_45546# a_1307_43914# 0.022061f
C424 a_n1925_42282# a_n913_45002# 0.017956f
C425 a_1823_45246# a_2809_45028# 0.076288f
C426 a_10903_43370# a_9482_43914# 1.20611f
C427 a_2324_44458# a_7705_45326# 0.029419f
C428 a_13717_47436# a_11453_44696# 0.041574f
C429 a_n971_45724# a_5807_45002# 0.0339f
C430 a_584_46384# a_768_44030# 0.105366f
C431 a_n1151_42308# a_9804_47204# 0.108722f
C432 a_4791_45118# a_n1613_43370# 0.223884f
C433 a_10227_46804# a_18780_47178# 0.050298f
C434 a_18143_47464# a_18479_47436# 0.238309f
C435 a_n3674_38216# a_n3420_39072# 0.020386f
C436 a_n4318_38216# a_n4064_39072# 0.023072f
C437 a_1209_43370# a_1049_43396# 0.194938f
C438 a_n97_42460# a_n1557_42282# 0.149645f
C439 a_15493_43940# a_16137_43396# 0.043956f
C440 a_15493_43396# a_18783_43370# 0.029898f
C441 a_526_44458# a_3363_44484# 0.119556f
C442 a_17715_44484# a_17517_44484# 0.163303f
C443 a_13059_46348# a_13483_43940# 0.124566f
C444 a_13259_45724# a_13076_44458# 0.188498f
C445 a_4185_45028# a_22485_44484# 0.080982f
C446 a_n2293_46634# a_8791_43396# 0.010288f
C447 a_n2109_47186# a_5497_46414# 0.017063f
C448 a_584_46384# a_1176_45822# 0.039976f
C449 a_13507_46334# a_16388_46812# 0.083261f
C450 a_n237_47217# a_3147_46376# 0.052931f
C451 a_n971_45724# a_3699_46348# 0.013334f
C452 a_4791_45118# a_n2293_46098# 0.411939f
C453 a_13070_42354# VDD 0.18656f
C454 a_22485_38105# a_22527_39145# 0.984424f
C455 a_21259_43561# a_4190_30871# 0.198353f
C456 a_17730_32519# a_14097_32519# 0.053763f
C457 a_n2293_43922# a_5934_30871# 0.079987f
C458 a_19862_44208# a_20922_43172# 0.164553f
C459 a_5111_44636# a_4743_44484# 0.02485f
C460 a_5147_45002# a_5343_44458# 0.063193f
C461 a_16019_45002# a_16237_45028# 0.053167f
C462 a_3537_45260# a_8103_44636# 0.140404f
C463 a_12891_46348# a_13259_45724# 1.04614f
C464 a_4791_45118# a_7230_45938# 0.010716f
C465 a_765_45546# a_17829_46910# 0.069261f
C466 a_17339_46660# a_18285_46348# 0.184197f
C467 C2_N_btm VDD 0.268945f
C468 C10_P_btm VREF 14.773f
C469 C5_N_btm C9_N_btm 0.150576f
C470 C4_N_btm C10_N_btm 0.703336f
C471 C6_N_btm C8_N_btm 0.163943f
C472 C8_P_btm VIN_P 0.907642f
C473 a_4905_42826# a_5379_42460# 0.077171f
C474 a_n97_42460# a_5934_30871# 0.221607f
C475 a_n2312_40392# a_n2302_40160# 0.151095f
C476 a_1307_43914# a_9028_43914# 0.010468f
C477 a_12883_44458# a_n2293_43922# 0.06281f
C478 a_11823_42460# a_14579_43548# 0.106967f
C479 a_6945_45028# a_22223_46124# 0.17119f
C480 a_8016_46348# a_8049_45260# 0.09608f
C481 a_765_45546# a_n443_42852# 0.232932f
C482 a_21076_30879# a_20205_31679# 0.055235f
C483 a_n2661_46634# a_2437_43646# 0.02989f
C484 a_4883_46098# a_9482_43914# 0.025151f
C485 a_5342_30871# a_14456_42282# 0.160195f
C486 a_9801_43940# VDD 0.19512f
C487 a_n1761_44111# a_n1644_44306# 0.170098f
C488 a_11967_42832# a_17737_43940# 0.054562f
C489 a_n913_45002# a_8387_43230# 0.024148f
C490 a_22612_30879# C10_N_btm 1.5848f
C491 a_20916_46384# VDD 0.302226f
C492 a_9290_44172# a_11633_42558# 0.014294f
C493 a_n1925_42282# a_1755_42282# 0.019802f
C494 a_526_44458# a_2123_42473# 0.012631f
C495 a_8049_45260# a_11682_45822# 0.011453f
C496 a_3877_44458# a_n699_43396# 0.061672f
C497 a_4646_46812# a_4223_44672# 0.018453f
C498 a_n443_46116# a_895_43940# 0.163929f
C499 a_12549_44172# a_n2661_42834# 0.04571f
C500 a_n755_45592# a_3175_45822# 0.046968f
C501 a_509_45822# a_n443_42852# 0.035689f
C502 a_16375_45002# a_10193_42453# 0.125364f
C503 a_5534_30871# C6_N_btm 0.01116f
C504 a_4700_47436# a_n443_46116# 0.255594f
C505 a_n1151_42308# a_6545_47178# 0.01616f
C506 a_12545_42858# VDD 0.285703f
C507 a_5379_42460# a_6123_31319# 0.011994f
C508 a_4921_42308# a_5932_42308# 0.194195f
C509 a_n1794_35082# a_5742_30871# 1.85696f
C510 a_6165_46155# VDD 0.204296f
C511 a_13747_46662# a_21381_43940# 0.030122f
C512 a_n1925_42282# a_n2661_44458# 0.029506f
C513 a_2324_44458# a_14539_43914# 0.028976f
C514 a_3090_45724# a_3905_42865# 0.025179f
C515 a_7227_45028# a_7229_43940# 0.019397f
C516 a_13249_42308# a_n2017_45002# 0.030327f
C517 a_4883_46098# a_7715_46873# 0.01159f
C518 a_10227_46804# a_10249_46116# 0.137273f
C519 a_n4064_40160# a_n3420_38528# 0.057096f
C520 a_n4209_39304# a_n4334_39392# 0.253307f
C521 a_n4315_30879# a_n4064_38528# 0.034153f
C522 a_n4318_38216# VDD 0.538766f
C523 a_n4209_39590# a_n4209_38502# 0.031979f
C524 a_10341_43396# a_16547_43609# 0.026476f
C525 a_10210_45822# VDD 0.323342f
C526 a_4185_45028# a_14401_32519# 0.040395f
C527 a_2711_45572# a_11967_42832# 0.068241f
C528 a_9290_44172# a_9165_43940# 0.01396f
C529 a_19479_31679# a_22223_45036# 0.01502f
C530 a_n1613_43370# a_6945_45028# 0.049203f
C531 a_n971_45724# a_n755_45592# 0.347347f
C532 a_2063_45854# a_n2661_45546# 0.038547f
C533 a_12251_46660# a_12359_47026# 0.057222f
C534 a_14976_45028# a_15227_44166# 0.035507f
C535 a_13747_46662# a_10903_43370# 0.027209f
C536 a_n743_46660# a_5164_46348# 0.031878f
C537 a_12549_44172# a_17715_44484# 0.03426f
C538 a_n2661_46098# a_472_46348# 0.065456f
C539 a_22629_37990# a_22725_37990# 0.087835f
C540 VDAC_P C7_P_btm 0.11042p
C541 a_3754_38470# RST_Z 0.203816f
C542 a_13460_43230# a_5534_30871# 0.052631f
C543 a_21101_45002# VDD 0.2903f
C544 a_17538_32519# a_14097_32519# 0.050981f
C545 a_n97_42460# a_16245_42852# 0.088473f
C546 en_comp a_n3674_39768# 0.036087f
C547 a_18479_45785# a_15493_43940# 0.016583f
C548 a_n2312_38680# a_n4318_38216# 0.023247f
C549 a_10227_46804# a_14113_42308# 0.627404f
C550 a_2382_45260# a_3600_43914# 0.158274f
C551 a_768_44030# a_8696_44636# 0.031444f
C552 a_1823_45246# a_2324_44458# 0.069409f
C553 a_8016_46348# a_8953_45546# 0.060003f
C554 a_14035_46660# a_14180_46482# 0.157972f
C555 a_18143_47464# a_2437_43646# 0.013364f
C556 a_5257_43370# a_2711_45572# 0.082068f
C557 a_4361_42308# a_11551_42558# 0.011423f
C558 a_3935_42891# a_3823_42558# 0.012124f
C559 a_n2293_42834# a_3080_42308# 0.021566f
C560 a_19778_44110# a_19741_43940# 0.054731f
C561 a_n2661_42834# a_7542_44172# 0.019328f
C562 a_19279_43940# a_21398_44850# 0.183186f
C563 a_n1435_47204# CLK 1.41989f
C564 a_16023_47582# VDD 0.201413f
C565 a_3090_45724# a_5147_45002# 0.023629f
C566 a_765_45546# a_2437_43646# 0.030322f
C567 a_12741_44636# a_18479_45785# 0.035678f
C568 a_4646_46812# a_n2293_42834# 0.152973f
C569 a_8199_44636# a_8192_45572# 0.04905f
C570 a_n3674_38680# a_n3674_37592# 0.028019f
C571 a_15493_43940# a_14021_43940# 0.08284f
C572 a_10405_44172# a_10555_43940# 0.018661f
C573 a_n755_45592# a_n2293_45010# 0.159033f
C574 a_15143_45578# a_15037_45618# 0.13675f
C575 a_12549_44172# a_20623_43914# 0.033887f
C576 a_13661_43548# a_15682_43940# 0.055235f
C577 a_15227_44166# a_15433_44458# 0.026124f
C578 a_16327_47482# a_19319_43548# 0.021453f
C579 a_n1151_42308# a_3877_44458# 0.019733f
C580 a_n443_46116# a_3067_47026# 0.030121f
C581 a_13507_46334# a_19321_45002# 0.034054f
C582 a_12465_44636# a_5807_45002# 0.59474f
C583 a_4883_46098# a_13747_46662# 0.050962f
C584 a_19511_42282# a_20712_42282# 0.05034f
C585 a_n97_42460# a_16547_43609# 0.066612f
C586 a_19721_31679# a_14097_32519# 0.051111f
C587 a_n23_45546# VDD 0.150941f
C588 a_n2661_45546# a_n2661_42834# 0.029567f
C589 a_10227_46804# a_5534_30871# 0.304847f
C590 a_3065_45002# a_3537_45260# 0.162384f
C591 a_7499_43078# a_5343_44458# 0.050528f
C592 a_4791_45118# a_6945_45028# 0.493927f
C593 a_12861_44030# a_13759_46122# 0.032694f
C594 a_11599_46634# a_10903_43370# 0.439916f
C595 a_7577_46660# a_8035_47026# 0.027606f
C596 a_n743_46660# a_16388_46812# 0.035819f
C597 a_n2661_46634# a_765_45546# 1.82448f
C598 a_10467_46802# a_10249_46116# 0.12624f
C599 a_10428_46928# a_6755_46942# 0.155315f
C600 a_10623_46897# a_10554_47026# 0.209641f
C601 a_n4315_30879# VREF_GND 0.168163f
C602 a_1169_39587# VDD 0.531695f
C603 a_n4209_37414# a_n3420_37440# 0.245806f
C604 a_14797_45144# VDD 0.124624f
C605 a_10775_45002# CLK 0.058141f
C606 a_5205_44484# a_n2661_42834# 0.030553f
C607 a_526_44458# a_9803_43646# 0.170855f
C608 a_5807_45002# a_2711_45572# 0.065611f
C609 a_15227_44166# a_19900_46494# 0.053335f
C610 a_14035_46660# a_13925_46122# 0.207108f
C611 a_n2472_46090# a_n2293_46098# 0.176709f
C612 a_19466_46812# a_19335_46494# 0.017838f
C613 a_8605_42826# a_8495_42852# 0.097745f
C614 a_20766_44850# VDD 0.197657f
C615 a_4223_44672# a_5013_44260# 0.07599f
C616 a_n913_45002# a_3539_42460# 0.359316f
C617 a_10227_46804# a_11691_44458# 0.012084f
C618 a_11453_44696# a_16922_45042# 0.07136f
C619 a_13507_46334# a_18184_42460# 0.505552f
C620 a_4791_45118# a_8103_44636# 0.048713f
C621 a_18597_46090# a_11827_44484# 0.039373f
C622 a_7287_43370# VDD 0.457521f
C623 a_18494_42460# a_4361_42308# 0.061307f
C624 a_8492_46660# VDD 0.273866f
C625 a_n863_45724# a_2351_42308# 0.038802f
C626 a_n755_45592# a_961_42354# 0.01273f
C627 a_5937_45572# a_1307_43914# 0.101589f
C628 a_526_44458# a_n913_45002# 0.250864f
C629 a_n1925_42282# a_n1059_45260# 0.023119f
C630 a_10903_43370# a_13348_45260# 0.011259f
C631 a_2324_44458# a_6709_45028# 0.076559f
C632 a_17339_46660# a_11691_44458# 0.018074f
C633 a_13717_47436# SMPL_ON_N 0.132417f
C634 a_11599_46634# a_4883_46098# 0.261488f
C635 a_n1151_42308# a_8128_46384# 0.328697f
C636 a_10227_46804# a_18479_47436# 1.40697f
C637 a_458_43396# a_1049_43396# 0.052073f
C638 a_15493_43396# a_18525_43370# 0.031354f
C639 a_526_44458# a_556_44484# 0.077901f
C640 a_n2293_46634# a_8147_43396# 0.011922f
C641 a_19692_46634# a_15493_43940# 0.16692f
C642 a_584_46384# a_1208_46090# 0.034313f
C643 a_13507_46334# a_13059_46348# 0.192049f
C644 a_n237_47217# a_2804_46116# 0.039625f
C645 a_n971_45724# a_3483_46348# 0.211534f
C646 a_n881_46662# a_15368_46634# 0.023127f
C647 a_n4209_39304# a_n3565_37414# 0.030571f
C648 a_12563_42308# VDD 0.254292f
C649 a_n3565_39304# a_n4209_37414# 0.028483f
C650 a_n2946_37984# a_n4064_37984# 0.053263f
C651 a_22485_38105# a_22589_40055# 0.212168f
C652 a_8953_45546# a_8791_43396# 0.012124f
C653 a_5111_44636# a_n699_43396# 0.016349f
C654 a_1307_43914# a_11691_44458# 0.024289f
C655 a_n743_46660# a_5066_45546# 0.124676f
C656 a_10227_46804# a_n443_42852# 0.043674f
C657 a_2063_45854# a_11322_45546# 0.105268f
C658 a_19692_46634# a_12741_44636# 0.022879f
C659 C1_N_btm VDD 0.264503f
C660 C6_N_btm C7_N_btm 26.0771f
C661 C5_N_btm C8_N_btm 0.145019f
C662 C3_N_btm C10_N_btm 0.321945f
C663 C4_N_btm C9_N_btm 0.154834f
C664 C9_P_btm VIN_P 1.82823f
C665 a_4905_42826# a_5267_42460# 0.146764f
C666 a_n23_44458# VDD 0.169093f
C667 a_3232_43370# a_11341_43940# 0.112367f
C668 a_n2312_40392# a_n4064_40160# 0.103899f
C669 a_12607_44458# a_n2293_43922# 0.078602f
C670 a_11823_42460# a_13667_43396# 0.107673f
C671 a_22612_30879# a_19479_31679# 0.064572f
C672 a_5937_45572# a_8034_45724# 0.052916f
C673 a_3090_45724# a_7499_43078# 0.23734f
C674 a_n2065_43946# a_n1644_44306# 0.090164f
C675 a_11967_42832# a_15682_43940# 1.63211f
C676 a_895_43940# a_2675_43914# 0.099822f
C677 a_n913_45002# a_8605_42826# 0.019641f
C678 a_19594_46812# START 0.020669f
C679 a_9290_44172# a_11551_42558# 0.123803f
C680 a_n1925_42282# a_1606_42308# 0.065478f
C681 a_n357_42282# a_7309_42852# 0.016177f
C682 a_n443_46116# a_2479_44172# 0.732848f
C683 a_11415_45002# a_6171_45002# 1.05801f
C684 a_16327_47482# a_3422_30871# 0.220296f
C685 a_6755_46942# a_11827_44484# 0.529579f
C686 a_n755_45592# a_2711_45572# 0.168218f
C687 a_4700_47436# a_4791_45118# 0.31818f
C688 a_n1151_42308# a_6151_47436# 0.026437f
C689 a_12089_42308# VDD 0.807892f
C690 a_9313_44734# a_10083_42826# 0.013808f
C691 a_18579_44172# a_4190_30871# 0.052036f
C692 a_5497_46414# VDD 0.200657f
C693 a_3483_46348# a_9313_44734# 0.015646f
C694 a_2711_45572# a_13017_45260# 0.050114f
C695 a_526_44458# a_n2661_44458# 0.087308f
C696 a_11415_45002# a_14673_44172# 0.229077f
C697 a_n443_42852# a_1307_43914# 0.05746f
C698 a_7227_45028# a_7276_45260# 0.098279f
C699 a_n1613_43370# a_3067_47026# 0.013046f
C700 a_10227_46804# a_10554_47026# 0.166977f
C701 a_n2472_42282# VDD 0.278905f
C702 a_n784_42308# C1_N_btm 0.027772f
C703 a_10341_43396# a_16243_43396# 0.058241f
C704 a_9313_44734# a_14097_32519# 0.053061f
C705 a_2382_45260# a_n2661_43370# 0.03415f
C706 a_19479_31679# a_11827_44484# 0.01397f
C707 a_22223_45572# a_22223_45036# 0.026152f
C708 a_n2661_46098# a_376_46348# 0.060405f
C709 a_n971_45724# a_n357_42282# 0.271282f
C710 a_584_46384# a_n2661_45546# 0.100439f
C711 a_12469_46902# a_12359_47026# 0.097745f
C712 a_12251_46660# a_12156_46660# 0.049827f
C713 a_3090_45724# a_15227_44166# 0.428743f
C714 a_n746_45260# a_310_45028# 0.378188f
C715 a_3754_38470# VDD 2.52245f
C716 VDAC_P C8_P_btm 0.220914p
C717 a_22629_38406# a_22737_37285# 0.08753f
C718 a_13635_43156# a_5534_30871# 0.078849f
C719 a_21005_45260# VDD 0.184261f
C720 a_n2956_37592# a_n3674_39768# 0.024317f
C721 a_3357_43084# a_n2661_42282# 0.028477f
C722 a_n443_42852# a_9396_43370# 0.039136f
C723 a_9290_44172# a_10341_42308# 0.051084f
C724 a_2382_45260# a_2998_44172# 0.045272f
C725 a_n2956_38680# a_n4318_38680# 0.023283f
C726 a_n2442_46660# a_n3674_38216# 0.023932f
C727 a_12549_44172# a_8696_44636# 0.035105f
C728 a_3483_46348# a_12594_46348# 0.011082f
C729 a_8016_46348# a_5937_45572# 0.021789f
C730 a_8349_46414# a_8199_44636# 0.032352f
C731 a_10227_46804# a_2437_43646# 0.150025f
C732 a_4361_42308# a_5742_30871# 0.071684f
C733 a_n1059_45260# a_15743_43084# 0.101833f
C734 a_n2661_42834# a_7281_43914# 0.010117f
C735 a_11967_42832# a_20512_43084# 0.106819f
C736 a_16327_47482# VDD 2.81451f
C737 a_3090_45724# a_4558_45348# 0.147318f
C738 a_6755_46942# a_15595_45028# 0.012879f
C739 a_n1613_43370# a_6298_44484# 0.02075f
C740 a_n1736_42282# a_n1329_42308# 0.050456f
C741 a_20692_30879# a_413_45260# 0.111034f
C742 a_n971_45724# a_n144_43396# 0.010576f
C743 a_13259_45724# a_6171_45002# 0.068737f
C744 a_n357_42282# a_n2293_45010# 0.020718f
C745 a_13661_43548# a_14955_43940# 0.010124f
C746 a_12549_44172# a_20365_43914# 0.069119f
C747 a_n2293_46634# a_n2661_42282# 0.039408f
C748 a_20894_47436# a_20843_47204# 0.134298f
C749 a_10227_46804# a_n2661_46634# 0.030546f
C750 a_4883_46098# a_13661_43548# 0.032161f
C751 a_19647_42308# a_13258_32519# 0.153411f
C752 a_19511_42282# a_20107_42308# 0.043647f
C753 a_17303_42282# a_22397_42558# 0.012536f
C754 a_10807_43548# a_10341_42308# 0.099222f
C755 a_18114_32519# a_14097_32519# 0.054468f
C756 a_9313_44734# a_22959_42860# 0.174475f
C757 a_n2956_37592# a_n4315_30879# 0.107228f
C758 a_n356_45724# VDD 0.719282f
C759 a_2437_43646# a_1307_43914# 0.160142f
C760 a_n357_42282# a_9313_44734# 5.02008f
C761 a_3065_45002# a_3429_45260# 0.037292f
C762 a_n237_47217# a_n1925_42282# 0.109762f
C763 a_11599_46634# a_11387_46155# 0.035936f
C764 a_12465_44636# a_3483_46348# 0.210833f
C765 a_7577_46660# a_7832_46660# 0.056391f
C766 a_n743_46660# a_13059_46348# 0.060636f
C767 a_10467_46802# a_10554_47026# 0.07009f
C768 a_10428_46928# a_10249_46116# 0.704177f
C769 a_10227_46804# a_8199_44636# 0.460391f
C770 a_n4064_40160# VIN_P 0.062574f
C771 a_n4315_30879# VREF 1.73216f
C772 a_n4209_37414# a_n3690_37440# 0.046103f
C773 a_14537_43396# VDD 0.779752f
C774 a_8953_45002# CLK 0.310391f
C775 a_4185_45028# a_5649_42852# 8.049951f
C776 a_11827_44484# a_20193_45348# 0.051742f
C777 a_10193_42453# a_11341_43940# 0.082222f
C778 a_6171_45002# a_n2661_43922# 0.020767f
C779 a_12465_44636# a_14495_45572# 0.019417f
C780 a_15227_44166# a_20075_46420# 0.060002f
C781 a_14035_46660# a_13759_46122# 0.162408f
C782 a_13887_32519# a_14097_32519# 10.5943f
C783 a_8037_42858# a_8495_42852# 0.027317f
C784 a_20835_44721# VDD 0.198384f
C785 a_3232_43370# a_n97_42460# 0.113391f
C786 a_n913_45002# a_3626_43646# 0.104422f
C787 a_n1059_45260# a_3539_42460# 0.021504f
C788 a_4223_44672# a_5244_44056# 0.019617f
C789 a_2107_46812# a_8953_45002# 0.016508f
C790 a_3483_46348# a_2711_45572# 0.167588f
C791 a_4791_45118# a_6298_44484# 0.033887f
C792 a_6547_43396# VDD 0.219105f
C793 a_18184_42460# a_4361_42308# 0.058569f
C794 a_n2293_42834# a_1847_42826# 0.078127f
C795 a_8667_46634# VDD 0.39254f
C796 a_n863_45724# a_2123_42473# 0.036254f
C797 a_n755_45592# a_1184_42692# 0.016193f
C798 a_8199_44636# a_1307_43914# 0.044343f
C799 a_526_44458# a_n1059_45260# 0.097646f
C800 a_n1925_42282# a_n2017_45002# 0.041988f
C801 a_n2312_39304# a_n3674_39768# 0.023328f
C802 a_13717_47436# a_22731_47423# 0.109987f
C803 a_10227_46804# a_18143_47464# 0.112443f
C804 a_2063_45854# a_11309_47204# 0.141276f
C805 a_14456_42282# a_14113_42308# 0.038993f
C806 a_n3674_38680# a_n4064_39072# 0.020036f
C807 a_n4318_38216# a_n3420_39072# 0.032825f
C808 a_3537_45260# a_4921_42308# 0.01091f
C809 a_458_43396# a_1209_43370# 0.0172f
C810 a_11967_42832# a_18249_42858# 0.018824f
C811 a_n97_42460# a_4905_42826# 0.147727f
C812 a_n2661_42282# a_743_42282# 0.043675f
C813 a_15493_43396# a_18429_43548# 0.045352f
C814 a_13259_45724# a_12607_44458# 0.132105f
C815 a_n2293_46634# a_7112_43396# 0.012325f
C816 a_10903_43370# a_11967_42832# 0.02192f
C817 a_12891_46348# a_11901_46660# 0.028795f
C818 a_n881_46662# a_14976_45028# 0.020069f
C819 a_n2109_47186# a_5164_46348# 0.603312f
C820 a_584_46384# a_805_46414# 0.135394f
C821 a_2959_46660# a_3055_46660# 0.013793f
C822 a_n2661_46634# a_10467_46802# 0.033928f
C823 a_n237_47217# a_2698_46116# 0.032015f
C824 a_12465_44636# a_14513_46634# 0.01549f
C825 a_10227_46804# a_765_45546# 0.038035f
C826 a_11633_42558# VDD 0.193501f
C827 a_n3420_37984# a_n4064_37984# 8.18485f
C828 a_n2293_43922# a_6123_31319# 0.080985f
C829 a_20731_45938# VDD 0.142103f
C830 a_n356_44636# a_15803_42450# 0.078793f
C831 a_5111_44636# a_4223_44672# 0.418299f
C832 a_17339_46660# a_765_45546# 0.244447f
C833 a_2063_45854# a_10490_45724# 0.082703f
C834 a_19466_46812# a_12741_44636# 0.043645f
C835 C0_N_btm VDD 1.02806f
C836 C10_P_btm VIN_P 3.66034f
C837 C4_N_btm C8_N_btm 0.145646f
C838 C3_N_btm C9_N_btm 0.137552f
C839 C2_N_btm C10_N_btm 0.327137f
C840 C5_N_btm C7_N_btm 0.151416f
C841 a_21753_35474# VIN_N 0.029412f
C842 a_13887_32519# a_22959_42860# 0.012735f
C843 a_3626_43646# a_1755_42282# 0.119352f
C844 a_n97_42460# a_6123_31319# 0.182488f
C845 a_n356_44636# VDD 1.17667f
C846 a_12607_44458# a_n2661_43922# 0.060913f
C847 a_10193_42453# a_10341_43396# 0.064616f
C848 a_9482_43914# a_12429_44172# 0.0636f
C849 a_n2312_39304# a_n4315_30879# 0.033437f
C850 a_20820_30879# a_20692_30879# 8.973741f
C851 a_21588_30879# a_19479_31679# 0.055797f
C852 a_21137_46414# a_6945_45028# 0.042885f
C853 a_8199_44636# a_8034_45724# 0.127067f
C854 a_2982_43646# CAL_N 0.181412f
C855 a_9165_43940# VDD 0.192035f
C856 a_1414_42308# a_3600_43914# 0.012293f
C857 a_2479_44172# a_2675_43914# 0.061502f
C858 a_n913_45002# a_8037_42858# 0.316376f
C859 a_19321_45002# START 0.10793f
C860 a_9290_44172# a_5742_30871# 0.118117f
C861 a_21588_30879# C9_N_btm 0.786375f
C862 a_20843_47204# VDD 0.188032f
C863 a_526_44458# a_1606_42308# 0.011179f
C864 a_n357_42282# a_5837_42852# 0.01329f
C865 a_8049_45260# a_10907_45822# 0.010337f
C866 a_n443_46116# a_2127_44172# 0.196411f
C867 a_18597_46090# a_19279_43940# 0.021978f
C868 a_3090_45724# a_n2661_43370# 0.101361f
C869 a_997_45618# a_1260_45572# 0.010598f
C870 a_n357_42282# a_2711_45572# 0.039058f
C871 a_12379_42858# VDD 0.484153f
C872 a_4921_42308# a_5755_42308# 0.175841f
C873 a_5204_45822# VDD 0.359177f
C874 a_n2840_46634# a_n2661_46634# 0.180867f
C875 a_n1613_43370# a_2864_46660# 0.014165f
C876 a_4883_46098# a_5257_43370# 0.026597f
C877 a_10227_46804# a_10623_46897# 0.180903f
C878 a_n3674_38680# VDD 0.503323f
C879 a_n2302_39866# a_n2302_39072# 0.052227f
C880 a_n4064_40160# a_n3565_38502# 0.028121f
C881 a_n4315_30879# a_n3420_38528# 0.034192f
C882 a_n784_42308# C0_N_btm 0.281635f
C883 a_10341_43396# a_16137_43396# 0.021507f
C884 a_8697_45822# VDD 0.189893f
C885 a_n356_44636# a_n784_42308# 0.084978f
C886 a_2274_45254# a_n2661_43370# 0.019962f
C887 a_13249_42308# a_9313_44734# 0.031106f
C888 a_10193_42453# a_n2293_43922# 0.024214f
C889 a_5111_44636# a_n2293_42834# 0.110286f
C890 a_768_44030# a_2324_44458# 0.047942f
C891 a_n2661_46098# a_n1076_46494# 0.037593f
C892 a_n743_46660# a_4704_46090# 0.011859f
C893 a_11901_46660# a_12359_47026# 0.034619f
C894 a_n746_45260# a_n1099_45572# 0.015931f
C895 a_2107_46812# a_167_45260# 0.012514f
C896 VDAC_P C9_P_btm 0.441881p
C897 a_13635_43156# a_14543_43071# 0.013803f
C898 a_20567_45036# VDD 0.237324f
C899 a_14401_32519# a_14097_32519# 0.051264f
C900 a_10807_43548# a_5742_30871# 0.020937f
C901 a_n2956_37592# a_n4318_39768# 0.029002f
C902 a_10193_42453# a_n97_42460# 0.304653f
C903 a_5343_44458# a_5883_43914# 0.042199f
C904 a_n443_42852# a_8791_43396# 0.053902f
C905 a_n2810_45028# a_n3674_39768# 0.023163f
C906 a_18479_45785# a_11341_43940# 0.019493f
C907 a_9290_44172# a_10922_42852# 0.028552f
C908 a_6298_44484# a_8103_44636# 0.016067f
C909 a_n2956_39304# a_n4318_38680# 0.023405f
C910 a_n2956_38680# a_n3674_39304# 0.023431f
C911 a_n2956_39768# a_n4318_37592# 0.02357f
C912 a_n2312_38680# a_n3674_38680# 0.023204f
C913 a_12891_46348# a_8696_44636# 0.028033f
C914 a_n443_46116# a_2382_45260# 0.027844f
C915 a_n2661_46634# a_11682_45822# 0.010865f
C916 a_8016_46348# a_8199_44636# 0.33718f
C917 a_17591_47464# a_2437_43646# 0.013209f
C918 a_2063_45854# a_6171_45002# 0.029207f
C919 a_n1435_47204# DATA[5] 0.031859f
C920 a_n2017_45002# a_15743_43084# 0.049212f
C921 a_18494_42460# a_19319_43548# 0.016978f
C922 a_14539_43914# a_15493_43396# 0.024653f
C923 a_20766_44850# a_20980_44850# 0.097745f
C924 a_20679_44626# a_3422_30871# 0.078371f
C925 a_20835_44721# a_21398_44850# 0.049827f
C926 a_16241_47178# VDD 0.208959f
C927 a_2324_44458# a_11652_45724# 0.034041f
C928 a_11453_44696# a_17767_44458# 0.010225f
C929 a_3483_46348# a_14033_45822# 0.030627f
C930 a_12741_44636# a_16147_45260# 0.023061f
C931 a_9672_43914# a_9801_43940# 0.062574f
C932 a_742_44458# a_2905_42968# 0.15065f
C933 a_11341_43940# a_14021_43940# 3.06514f
C934 a_16721_46634# VDD 0.186443f
C935 a_n863_45724# a_n913_45002# 0.565852f
C936 a_20205_31679# a_413_45260# 0.034773f
C937 a_12549_44172# a_20269_44172# 0.049822f
C938 a_n755_45592# a_n2661_45010# 0.01648f
C939 a_n2956_38216# a_n2956_37592# 0.103811f
C940 a_13661_43548# a_13483_43940# 0.057042f
C941 a_584_46384# a_n1557_42282# 0.032459f
C942 a_n443_46116# a_3524_46660# 0.049574f
C943 a_13507_46334# a_13747_46662# 0.049663f
C944 a_4883_46098# a_5807_45002# 1.76125f
C945 a_19511_42282# a_13258_32519# 0.072135f
C946 a_n4318_37592# a_n4334_37440# 0.083644f
C947 a_10807_43548# a_10922_42852# 0.010566f
C948 en_comp a_22485_38105# 0.535686f
C949 a_n2810_45028# a_n4315_30879# 0.02588f
C950 a_9313_44734# a_22223_42860# 0.012144f
C951 a_3503_45724# VDD 0.129733f
C952 a_n97_42460# a_16137_43396# 0.134668f
C953 a_10227_46804# a_13460_43230# 0.243111f
C954 a_2382_45260# a_3537_45260# 0.250657f
C955 a_5937_45572# a_6756_44260# 0.010335f
C956 a_3483_46348# a_15682_43940# 0.261013f
C957 a_n237_47217# a_526_44458# 0.198088f
C958 a_12861_44030# a_12594_46348# 0.43362f
C959 a_7715_46873# a_7832_46660# 0.157972f
C960 a_n2109_47186# a_5066_45546# 0.02651f
C961 a_10428_46928# a_10554_47026# 0.181217f
C962 a_9863_46634# a_6755_46942# 0.014818f
C963 a_10467_46802# a_10623_46897# 0.107482f
C964 a_10150_46912# a_10249_46116# 0.066949f
C965 a_n4209_37414# a_n3565_37414# 6.90997f
C966 a_14180_45002# VDD 0.151315f
C967 a_4185_45028# a_13678_32519# 0.037732f
C968 a_11827_44484# a_11691_44458# 0.881979f
C969 a_3232_43370# a_n2661_43922# 0.197944f
C970 a_4791_45118# a_4921_42308# 0.172224f
C971 a_12465_44636# a_13249_42308# 0.541909f
C972 a_15227_44166# a_19335_46494# 0.024137f
C973 a_19466_46812# a_18985_46122# 0.033782f
C974 a_13887_32519# a_22400_42852# 0.098245f
C975 a_n4318_39304# a_n4064_40160# 0.062069f
C976 a_20679_44626# VDD 0.439119f
C977 a_18479_45785# a_10341_43396# 0.038969f
C978 a_n1059_45260# a_3626_43646# 0.025708f
C979 a_n2017_45002# a_3539_42460# 0.042001f
C980 a_4223_44672# a_3905_42865# 0.019153f
C981 a_11415_45002# a_10193_42453# 0.024787f
C982 a_18479_47436# a_11827_44484# 0.035345f
C983 a_n2497_47436# a_n356_44636# 0.019387f
C984 a_18597_46090# a_21101_45002# 0.033595f
C985 a_6765_43638# VDD 0.218204f
C986 a_18184_42460# a_13467_32519# 0.022572f
C987 a_10057_43914# a_10341_43396# 0.055207f
C988 a_n2293_43922# a_3080_42308# 0.084673f
C989 a_5891_43370# a_6293_42852# 0.107308f
C990 a_n755_45592# a_1576_42282# 0.025747f
C991 a_7927_46660# VDD 0.187888f
C992 a_n863_45724# a_1755_42282# 0.050501f
C993 a_16375_45002# a_16147_45260# 1.01554f
C994 a_526_44458# a_n2017_45002# 0.028467f
C995 a_2324_44458# a_7276_45260# 0.049304f
C996 a_n2312_40392# a_n3674_39768# 0.025146f
C997 a_n2312_39304# a_n4318_39768# 0.02345f
C998 a_2711_45572# a_13249_42308# 0.043493f
C999 a_3090_45724# a_5883_43914# 0.132458f
C1000 a_12861_44030# a_12465_44636# 0.242761f
C1001 a_11599_46634# a_13507_46334# 0.259318f
C1002 a_13575_42558# a_14113_42308# 0.11418f
C1003 a_n3674_37592# a_n4064_39616# 0.019733f
C1004 a_11967_42832# a_17333_42852# 0.14149f
C1005 a_n97_42460# a_3080_42308# 0.353977f
C1006 a_5111_44636# a_5379_42460# 0.118194f
C1007 a_15493_43396# a_17324_43396# 0.047612f
C1008 a_14021_43940# a_10341_43396# 1.5617f
C1009 a_n863_45724# a_n2661_44458# 0.091002f
C1010 a_15861_45028# a_6171_45002# 0.09425f
C1011 a_16327_47482# a_20556_43646# 0.014087f
C1012 a_4646_46812# a_n97_42460# 0.016161f
C1013 a_n2293_46634# a_7287_43370# 0.016986f
C1014 a_19692_46634# a_11341_43940# 0.06f
C1015 a_n881_46662# a_3090_45724# 0.107805f
C1016 a_584_46384# a_472_46348# 0.31609f
C1017 a_n2661_46634# a_10428_46928# 0.052586f
C1018 a_n237_47217# a_2521_46116# 0.039248f
C1019 a_n1151_42308# a_n1991_46122# 0.027139f
C1020 a_12465_44636# a_14180_46812# 0.026945f
C1021 a_4958_30871# EN_VIN_BSTR_N 0.021638f
C1022 a_n4209_39304# a_n4209_37414# 0.029637f
C1023 a_n3420_37984# a_n2946_37984# 0.238664f
C1024 a_n3690_38304# a_n4064_37984# 0.085872f
C1025 a_n3565_38216# a_n2302_37984# 0.067194f
C1026 a_22485_38105# a_22537_40625# 0.0722f
C1027 a_11551_42558# VDD 0.192086f
C1028 a_20528_45572# VDD 0.08228f
C1029 a_n356_44636# a_15764_42576# 0.012586f
C1030 a_5147_45002# a_4223_44672# 0.047867f
C1031 a_3537_45260# a_5343_44458# 0.378482f
C1032 a_n2312_39304# a_n2956_38216# 0.060648f
C1033 a_12861_44030# a_2711_45572# 0.104124f
C1034 a_2063_45854# a_8746_45002# 0.058531f
C1035 a_n443_46116# a_4880_45572# 0.048165f
C1036 a_n1925_46634# a_5066_45546# 0.195997f
C1037 EN_VIN_BSTR_N VCM 0.927954f
C1038 a_19998_34978# VIN_N 0.37444f
C1039 C3_N_btm C8_N_btm 0.134581f
C1040 C2_N_btm C9_N_btm 0.141891f
C1041 C1_N_btm C10_N_btm 0.31753f
C1042 C5_N_btm C6_N_btm 22.305399f
C1043 C4_N_btm C7_N_btm 0.145303f
C1044 a_13887_32519# a_22223_42860# 0.013362f
C1045 a_3080_42308# a_3823_42558# 0.016209f
C1046 a_n97_42460# a_7227_42308# 0.032716f
C1047 a_n755_45592# a_5649_42852# 0.02386f
C1048 a_n2293_42834# a_3905_42865# 0.039227f
C1049 a_8975_43940# a_n2661_43922# 0.11532f
C1050 a_2711_45572# a_19700_43370# 0.016505f
C1051 a_18479_45785# a_n97_42460# 0.072469f
C1052 a_20193_45348# a_19279_43940# 0.021458f
C1053 a_9482_43914# a_11750_44172# 0.020902f
C1054 a_n2312_40392# a_n4315_30879# 0.389397f
C1055 a_20820_30879# a_20205_31679# 0.087297f
C1056 a_8349_46414# a_8034_45724# 0.05863f
C1057 a_10227_46804# a_1307_43914# 0.081555f
C1058 a_n2472_43914# a_n3674_39768# 0.162742f
C1059 a_1414_42308# a_2998_44172# 0.447595f
C1060 a_n1059_45260# a_8037_42858# 0.048776f
C1061 a_19594_46812# VDD 0.349555f
C1062 a_2127_44172# a_2675_43914# 0.090298f
C1063 a_2479_44172# a_895_43940# 0.318312f
C1064 a_8049_45260# a_10210_45822# 0.01041f
C1065 a_13259_45724# a_10193_42453# 0.284945f
C1066 a_16327_47482# a_20980_44850# 0.012339f
C1067 a_10341_42308# VDD 0.931019f
C1068 a_n1741_47186# a_11599_46634# 0.164599f
C1069 a_4007_47204# a_4700_47436# 0.010942f
C1070 a_3785_47178# a_n443_46116# 0.040847f
C1071 a_8333_44056# a_8147_43396# 0.011009f
C1072 a_5164_46348# VDD 0.717083f
C1073 a_10193_42453# a_18057_42282# 0.099046f
C1074 a_1823_45246# a_3363_44484# 0.046566f
C1075 a_17339_46660# a_18579_44172# 0.016577f
C1076 a_11823_42460# a_n913_45002# 0.281323f
C1077 a_n2840_46634# a_n2956_39768# 0.156182f
C1078 a_n1613_43370# a_3524_46660# 0.28004f
C1079 a_n443_46116# a_3090_45724# 0.011392f
C1080 a_13747_46662# a_n743_46660# 0.042998f
C1081 a_10227_46804# a_10467_46802# 0.678578f
C1082 a_n2840_42282# VDD 0.294987f
C1083 a_2437_43646# a_11827_44484# 0.013953f
C1084 a_3232_43370# a_5837_45028# 0.01175f
C1085 a_19692_46634# a_10341_43396# 0.022785f
C1086 a_10193_42453# a_n2661_43922# 0.025533f
C1087 a_12549_44172# a_2324_44458# 0.506903f
C1088 a_n2661_46098# a_n901_46420# 0.054328f
C1089 a_15368_46634# a_15559_46634# 0.022471f
C1090 a_n743_46660# a_4419_46090# 0.032595f
C1091 a_11901_46660# a_12156_46660# 0.06121f
C1092 a_n971_45724# a_n1099_45572# 0.508925f
C1093 VDAC_Ni VDD 0.288547f
C1094 VDAC_P C10_P_btm 0.883474p
C1095 a_22629_38406# a_22629_37990# 0.32625f
C1096 a_13635_43156# a_13460_43230# 0.234322f
C1097 a_13113_42826# a_5534_30871# 0.024339f
C1098 a_18494_42460# VDD 0.73193f
C1099 a_10807_43548# a_11323_42473# 0.109765f
C1100 a_n443_42852# a_8147_43396# 0.060401f
C1101 a_n2810_45028# a_n4318_39768# 0.027945f
C1102 a_9290_44172# a_10991_42826# 0.045863f
C1103 a_13259_45724# a_16137_43396# 0.038525f
C1104 a_n2956_39304# a_n3674_39304# 0.029162f
C1105 a_n2442_46660# a_n4318_38216# 0.023718f
C1106 a_n443_46116# a_2274_45254# 0.041907f
C1107 a_8016_46348# a_8349_46414# 0.232167f
C1108 a_22959_46660# a_22959_46124# 0.026152f
C1109 a_3483_46348# a_10903_43370# 0.404121f
C1110 a_16327_47482# a_3357_43084# 0.114502f
C1111 a_2063_45854# a_3232_43370# 0.056568f
C1112 a_4361_42308# a_10723_42308# 0.010334f
C1113 a_16137_43396# a_18057_42282# 0.01884f
C1114 a_3499_42826# VDD 0.333472f
C1115 a_18184_42460# a_19319_43548# 0.032261f
C1116 a_n2661_42834# a_5663_43940# 0.01057f
C1117 a_20679_44626# a_21398_44850# 0.086708f
C1118 a_20835_44721# a_20980_44850# 0.057222f
C1119 a_15673_47210# VDD 0.569224f
C1120 a_n1435_47204# DATA[4] 0.033859f
C1121 a_9313_45822# CLK 0.027301f
C1122 a_12594_46348# a_13904_45546# 0.077346f
C1123 a_526_44458# a_4099_45572# 0.063912f
C1124 a_3090_45724# a_3537_45260# 0.198803f
C1125 a_n1613_43370# a_5343_44458# 0.03714f
C1126 a_11415_45002# a_18479_45785# 0.047896f
C1127 a_n1736_42282# a_n4318_37592# 0.153911f
C1128 a_1414_42308# a_1568_43370# 0.01352f
C1129 a_1467_44172# a_1756_43548# 0.100052f
C1130 a_16388_46812# VDD 0.797417f
C1131 a_n913_45002# a_20922_43172# 0.010679f
C1132 a_n863_45724# a_n1059_45260# 0.162875f
C1133 a_12549_44172# a_19862_44208# 0.262561f
C1134 a_n357_42282# a_n2661_45010# 0.017732f
C1135 a_n2956_38216# a_n2810_45028# 5.73989f
C1136 a_n2293_45546# a_n745_45366# 0.038459f
C1137 a_n443_46116# a_3699_46634# 0.036317f
C1138 a_13507_46334# a_13661_43548# 0.038602f
C1139 a_19787_47423# a_19594_46812# 0.108653f
C1140 a_11599_46634# a_n743_46660# 0.248412f
C1141 a_9313_45822# a_2107_46812# 0.298046f
C1142 a_133_42852# VDD 0.184203f
C1143 a_19511_42282# a_19647_42308# 0.038787f
C1144 a_n4318_37592# a_n4209_37414# 0.105251f
C1145 a_10807_43548# a_10991_42826# 0.01427f
C1146 a_9313_44734# a_22165_42308# 0.028818f
C1147 a_3316_45546# VDD 0.428912f
C1148 a_7499_43078# a_4223_44672# 0.02232f
C1149 a_10227_46804# a_13635_43156# 0.320228f
C1150 a_5937_45572# a_n2661_42282# 0.060993f
C1151 a_3483_46348# a_14955_43940# 0.242667f
C1152 a_2382_45260# a_3429_45260# 0.011518f
C1153 a_2680_45002# a_3065_45002# 0.13328f
C1154 a_n746_45260# a_526_44458# 0.096099f
C1155 a_n237_47217# a_2981_46116# 0.024703f
C1156 a_13507_46334# a_4185_45028# 0.479559f
C1157 a_10428_46928# a_10623_46897# 0.21686f
C1158 a_9863_46634# a_10249_46116# 0.027588f
C1159 a_8492_46660# a_6755_46942# 0.024647f
C1160 a_7411_46660# a_7832_46660# 0.086708f
C1161 a_10150_46912# a_10554_47026# 0.051162f
C1162 a_10227_46804# a_8016_46348# 0.093061f
C1163 a_11599_46634# a_11189_46129# 0.0158f
C1164 a_4883_46098# a_3483_46348# 0.813604f
C1165 a_n4209_37414# a_n4334_37440# 0.253282f
C1166 a_n2302_39866# VDD 0.361509f
C1167 a_n4315_30879# VIN_P 0.187f
C1168 a_743_42282# a_12089_42308# 0.016016f
C1169 a_13777_45326# VDD 0.145151f
C1170 a_3422_30871# a_5742_30871# 0.025558f
C1171 a_n357_42282# a_21381_43940# 0.060125f
C1172 a_3232_43370# a_n2661_42834# 0.127534f
C1173 a_11453_44696# a_11823_42460# 0.072491f
C1174 a_15227_44166# a_19553_46090# 0.047784f
C1175 a_19466_46812# a_18819_46122# 0.02948f
C1176 a_20640_44752# VDD 0.246486f
C1177 a_n357_42282# a_18249_42858# 0.047936f
C1178 a_n913_45002# a_2982_43646# 0.498826f
C1179 a_n699_43396# a_2998_44172# 0.127437f
C1180 a_n967_45348# a_n1557_42282# 0.092498f
C1181 a_n2017_45002# a_3626_43646# 0.023645f
C1182 a_10903_43370# a_n357_42282# 0.028411f
C1183 a_n2293_46098# a_4880_45572# 0.013174f
C1184 a_2063_45854# a_8975_43940# 0.149528f
C1185 a_20202_43084# a_10193_42453# 0.296862f
C1186 a_n2293_46634# a_14537_43396# 0.036569f
C1187 a_2324_44458# a_n2661_45546# 0.019247f
C1188 a_18597_46090# a_21005_45260# 0.034207f
C1189 a_6197_43396# VDD 0.408793f
C1190 a_n755_45592# a_1067_42314# 0.047422f
C1191 a_8145_46902# VDD 0.199702f
C1192 a_n863_45724# a_1606_42308# 0.20593f
C1193 a_5891_43370# a_6031_43396# 0.01824f
C1194 a_12861_44030# a_15682_43940# 0.016729f
C1195 a_4646_46812# a_n2661_43922# 0.06073f
C1196 a_9290_44172# a_9482_43914# 0.135239f
C1197 a_8016_46348# a_1307_43914# 0.035949f
C1198 a_10903_43370# a_11963_45334# 0.209081f
C1199 a_2324_44458# a_5205_44484# 0.523531f
C1200 a_n2312_40392# a_n4318_39768# 0.025298f
C1201 a_2711_45572# a_13904_45546# 0.021385f
C1202 a_16327_47482# a_18597_46090# 1.28053f
C1203 a_17591_47464# a_10227_46804# 0.292864f
C1204 a_13717_47436# a_12465_44636# 0.049141f
C1205 a_13575_42558# a_13657_42558# 0.171361f
C1206 a_n3674_38680# a_n3420_39072# 0.172947f
C1207 a_5934_30871# a_4958_30871# 0.018095f
C1208 a_11967_42832# a_18083_42858# 0.472348f
C1209 a_15493_43940# a_15781_43660# 0.049304f
C1210 a_n97_42460# a_4699_43561# 0.025323f
C1211 a_15493_43396# a_17499_43370# 0.038093f
C1212 a_5066_45546# VDD 1.34058f
C1213 a_5111_44636# a_5267_42460# 0.047489f
C1214 a_n913_45002# a_8325_42308# 0.233489f
C1215 a_15227_44166# a_15493_43940# 0.091653f
C1216 a_8696_44636# a_6171_45002# 0.070776f
C1217 a_7499_43078# a_n2293_42834# 0.352878f
C1218 a_n2293_46634# a_6547_43396# 0.010751f
C1219 a_16327_47482# a_743_42282# 0.026382f
C1220 a_12891_46348# a_11735_46660# 0.034334f
C1221 a_n1613_43370# a_3090_45724# 0.039515f
C1222 a_584_46384# a_376_46348# 0.232754f
C1223 a_n2661_46634# a_10150_46912# 0.010702f
C1224 a_n237_47217# a_167_45260# 0.280171f
C1225 a_n1151_42308# a_n1853_46287# 0.024093f
C1226 a_4958_30871# a_10890_34112# 0.021413f
C1227 a_5934_30871# VCM 0.121361f
C1228 a_n3565_38216# a_n4064_37984# 0.342209f
C1229 a_5742_30871# VDD 0.556723f
C1230 a_22485_38105# a_22589_40599# 0.132855f
C1231 a_15743_43084# a_22591_43396# 0.016556f
C1232 a_21188_45572# VDD 0.288663f
C1233 a_19479_31679# C1_N_btm 0.043983f
C1234 a_n4318_40392# a_n4064_40160# 0.077948f
C1235 a_8696_44636# a_14673_44172# 0.017655f
C1236 a_13259_45724# a_14021_43940# 0.028871f
C1237 a_3537_45260# a_4743_44484# 0.01411f
C1238 a_n443_42852# a_n2661_42282# 0.133617f
C1239 a_15227_44166# a_12741_44636# 0.250453f
C1240 a_19692_46634# a_11415_45002# 0.033537f
C1241 a_n2312_40392# a_n2956_38216# 0.053778f
C1242 a_n2661_46098# a_n1736_46482# 0.024986f
C1243 a_3090_45724# a_n2293_46098# 0.642755f
C1244 a_2063_45854# a_10193_42453# 0.114552f
C1245 EN_VIN_BSTR_N VREF_GND 0.857366f
C1246 C2_N_btm C8_N_btm 0.138777f
C1247 C1_N_btm C9_N_btm 0.132506f
C1248 C0_N_btm C10_N_btm 0.365593f
C1249 C4_N_btm C6_N_btm 0.143514f
C1250 C3_N_btm C7_N_btm 0.134911f
C1251 a_22223_43396# a_22223_42860# 0.026152f
C1252 a_3080_42308# a_3318_42354# 0.036372f
C1253 a_n97_42460# a_6761_42308# 0.012266f
C1254 a_2982_43646# a_1755_42282# 0.051666f
C1255 a_n357_42282# a_5649_42852# 0.011202f
C1256 a_11823_42460# a_9145_43396# 0.146085f
C1257 a_18184_42460# a_3422_30871# 0.649102f
C1258 a_10057_43914# a_n2661_43922# 0.034016f
C1259 a_8975_43940# a_n2661_42834# 0.083892f
C1260 a_n1151_42308# a_n2661_43370# 0.027798f
C1261 a_8016_46348# a_8034_45724# 0.254614f
C1262 a_5534_30871# a_13070_42354# 0.025818f
C1263 a_1414_42308# a_2889_44172# 0.128883f
C1264 a_13747_46662# START 0.062289f
C1265 a_n2840_43914# a_n3674_39768# 0.022122f
C1266 a_19321_45002# VDD 1.01574f
C1267 a_2127_44172# a_895_43940# 0.132679f
C1268 a_1823_45246# a_n913_45002# 0.041568f
C1269 a_18597_46090# a_20835_44721# 0.012854f
C1270 a_n443_46116# a_1414_42308# 0.18376f
C1271 a_18479_47436# a_19279_43940# 0.017993f
C1272 a_10922_42852# VDD 0.216186f
C1273 a_n971_45724# a_n1435_47204# 2.23698f
C1274 a_3785_47178# a_4791_45118# 0.010875f
C1275 a_n1151_42308# a_4915_47217# 0.1374f
C1276 a_n784_42308# a_5742_30871# 0.550812f
C1277 a_n356_44636# a_5342_30871# 0.133551f
C1278 a_5068_46348# VDD 0.085085f
C1279 a_n2017_45002# a_18707_42852# 0.026353f
C1280 a_7227_45028# a_6171_45002# 0.029883f
C1281 a_11823_42460# a_n1059_45260# 0.100641f
C1282 a_n1613_43370# a_3699_46634# 0.344308f
C1283 a_4915_47217# a_14084_46812# 0.038663f
C1284 a_4791_45118# a_3090_45724# 0.206257f
C1285 a_16327_47482# a_6755_46942# 0.067305f
C1286 a_10227_46804# a_10428_46928# 0.060058f
C1287 a_n4064_39616# a_n4064_39072# 0.062881f
C1288 a_n4064_40160# a_n4209_38502# 0.05515f
C1289 a_n4315_30879# a_n3565_38502# 0.085594f
C1290 a_21513_45002# a_11827_44484# 0.010541f
C1291 a_16019_45002# a_1307_43914# 0.01609f
C1292 a_5691_45260# a_5837_45028# 0.171361f
C1293 a_327_44734# a_n2661_43370# 0.035472f
C1294 a_10193_42453# a_n2661_42834# 0.034215f
C1295 a_12891_46348# a_2324_44458# 0.026746f
C1296 a_n2661_46098# a_n1641_46494# 0.035694f
C1297 a_n743_46660# a_4185_45028# 0.036891f
C1298 a_11813_46116# a_12156_46660# 0.157972f
C1299 a_16327_47482# a_8049_45260# 0.605463f
C1300 a_7754_38636# VDD 0.036155f
C1301 CAL_P a_22629_37990# 0.205295f
C1302 a_22629_38406# a_22725_38406# 0.090011f
C1303 a_12545_42858# a_5534_30871# 0.17182f
C1304 a_18184_42460# VDD 2.05053f
C1305 a_n357_42282# a_8685_43396# 0.319118f
C1306 a_9290_44172# a_10796_42968# 0.050429f
C1307 a_n2956_39768# a_n3674_38216# 0.023755f
C1308 a_15227_44166# a_16375_45002# 0.117865f
C1309 a_16763_47508# a_2437_43646# 0.014946f
C1310 a_22959_46660# a_10809_44734# 0.015306f
C1311 a_584_46384# a_3232_43370# 0.277433f
C1312 a_4361_42308# a_10533_42308# 0.017218f
C1313 a_16922_45042# a_20974_43370# 0.077191f
C1314 a_20640_44752# a_21398_44850# 0.056391f
C1315 a_11459_47204# DATA[5] 0.370451f
C1316 a_15811_47375# VDD 0.979053f
C1317 a_n1435_47204# DATA[3] 0.02843f
C1318 a_12594_46348# a_13527_45546# 0.100424f
C1319 a_6755_46942# a_14537_43396# 0.120241f
C1320 a_17715_44484# a_10193_42453# 0.074403f
C1321 a_8199_44636# a_10907_45822# 0.081841f
C1322 a_2324_44458# a_11322_45546# 0.068998f
C1323 a_10903_43370# a_13249_42308# 0.211356f
C1324 a_n1925_42282# a_2711_45572# 0.019937f
C1325 a_n3674_38216# a_n4318_37592# 2.7294f
C1326 a_9028_43914# a_9420_43940# 0.016359f
C1327 a_n3674_39768# a_n4318_39304# 2.75695f
C1328 a_n356_44636# a_743_42282# 0.063042f
C1329 a_13059_46348# VDD 0.955445f
C1330 a_1467_44172# a_1568_43370# 0.055004f
C1331 a_742_44458# a_1847_42826# 0.372436f
C1332 a_9313_44734# a_15743_43084# 1.48048f
C1333 a_13259_45724# a_21613_42308# 0.077442f
C1334 a_13904_45546# a_14033_45822# 0.062574f
C1335 a_8746_45002# a_8696_44636# 0.058163f
C1336 a_10193_42453# a_15861_45028# 0.432483f
C1337 a_n863_45724# a_n2017_45002# 0.111825f
C1338 a_12861_44030# a_21381_43940# 0.019154f
C1339 a_1823_45246# a_n2661_44458# 0.036985f
C1340 a_12549_44172# a_19478_44306# 0.010691f
C1341 a_n2293_45546# a_n913_45002# 0.043147f
C1342 a_2063_45854# a_4646_46812# 0.093604f
C1343 a_n443_46116# a_2959_46660# 0.036727f
C1344 a_13507_46334# a_5807_45002# 1.64614f
C1345 a_19787_47423# a_19321_45002# 0.029499f
C1346 a_19386_47436# a_19594_46812# 0.069651f
C1347 a_18479_47436# a_20916_46384# 0.014237f
C1348 a_10807_43548# a_10796_42968# 0.030352f
C1349 a_8791_43396# a_9396_43370# 0.011032f
C1350 a_9313_44734# a_21671_42860# 0.012466f
C1351 a_3218_45724# VDD 0.133843f
C1352 a_3483_46348# a_13483_43940# 0.194464f
C1353 a_10227_46804# a_12895_43230# 0.152365f
C1354 a_20202_43084# a_14021_43940# 0.020234f
C1355 a_2382_45260# a_3065_45002# 0.632538f
C1356 a_n971_45724# a_526_44458# 0.21769f
C1357 a_n1151_42308# a_10809_44734# 0.334692f
C1358 a_19594_46812# a_19551_46910# 0.07027f
C1359 a_8667_46634# a_6755_46942# 0.011524f
C1360 a_10428_46928# a_10467_46802# 0.820079f
C1361 a_12861_44030# a_10903_43370# 0.378457f
C1362 a_n4064_39616# VDD 1.68728f
C1363 a_n2661_42282# COMP_P 0.02767f
C1364 a_13556_45296# VDD 0.569056f
C1365 a_626_44172# a_n356_44636# 0.249281f
C1366 a_4185_45028# a_4361_42308# 0.042181f
C1367 a_3232_43370# a_11649_44734# 0.011508f
C1368 a_15227_44166# a_18985_46122# 0.287996f
C1369 a_n2438_43548# a_n755_45592# 0.213107f
C1370 a_13678_32519# a_14097_32519# 0.04945f
C1371 a_20362_44736# VDD 0.275577f
C1372 a_5111_44636# a_n97_42460# 0.211832f
C1373 a_n357_42282# a_17333_42852# 0.05273f
C1374 a_n1059_45260# a_2982_43646# 0.020128f
C1375 a_4223_44672# a_2998_44172# 0.035464f
C1376 a_n2661_44458# a_n3674_39768# 0.037999f
C1377 a_14537_43396# a_15037_43940# 0.018234f
C1378 a_16327_47482# a_20193_45348# 0.359904f
C1379 a_19335_46494# a_19443_46116# 0.057222f
C1380 a_2063_45854# a_10057_43914# 0.06633f
C1381 a_10227_46804# a_11827_44484# 0.065169f
C1382 a_n443_46116# a_n699_43396# 0.042248f
C1383 a_4791_45118# a_4743_44484# 0.165321f
C1384 a_13291_42460# a_14635_42282# 0.111986f
C1385 a_6293_42852# VDD 0.401011f
C1386 a_n2293_42282# a_n1794_35082# 0.18361f
C1387 a_n755_45592# a_n1794_35082# 0.044103f
C1388 a_7577_46660# VDD 0.249866f
C1389 a_17339_46660# a_11827_44484# 0.031147f
C1390 a_3877_44458# a_n2661_43922# 0.021496f
C1391 a_4646_46812# a_n2661_42834# 0.030297f
C1392 a_2324_44458# a_6431_45366# 0.046214f
C1393 a_22959_46124# a_413_45260# 0.020082f
C1394 a_16588_47582# a_10227_46804# 0.039575f
C1395 a_n1741_47186# a_5807_45002# 0.029376f
C1396 a_2063_45854# a_9804_47204# 0.249806f
C1397 a_12861_44030# a_4883_46098# 0.076083f
C1398 a_n1151_42308# a_n881_46662# 1.41446f
C1399 a_n1794_35082# a_n3565_39590# 0.035115f
C1400 a_n3674_37592# a_n3420_39616# 0.019754f
C1401 a_14021_43940# a_14955_43396# 0.01294f
C1402 a_11967_42832# a_17701_42308# 0.030406f
C1403 a_15493_43940# a_15681_43442# 0.03571f
C1404 a_15493_43396# a_16759_43396# 0.029803f
C1405 a_n2017_45002# a_8685_42308# 0.016058f
C1406 en_comp a_5934_30871# 0.028707f
C1407 a_8696_44636# a_3232_43370# 0.169534f
C1408 a_n2293_46634# a_6765_43638# 0.011639f
C1409 a_n237_47217# a_2202_46116# 0.049087f
C1410 a_n1151_42308# a_n2157_46122# 0.027101f
C1411 a_4915_47217# a_12741_44636# 0.031734f
C1412 a_n743_46660# a_5257_43370# 0.036418f
C1413 a_n1925_46634# a_7715_46873# 0.01948f
C1414 a_n2661_46634# a_9863_46634# 0.010932f
C1415 a_n746_45260# a_167_45260# 0.234425f
C1416 a_n4334_38304# a_n4064_37984# 0.410244f
C1417 a_n3690_38304# a_n3420_37984# 0.414894f
C1418 a_n3565_38216# a_n2946_37984# 0.411006f
C1419 a_n4209_38216# a_n2302_37984# 0.407312f
C1420 a_2684_37794# a_2113_38308# 0.468006f
C1421 a_n4315_30879# VDAC_P 0.011363f
C1422 a_11323_42473# VDD 0.205172f
C1423 a_22485_38105# CAL_N 0.072058f
C1424 a_3422_30871# a_20753_42852# 0.048434f
C1425 a_n4318_40392# a_n4334_40480# 0.089305f
C1426 a_15743_43084# a_13887_32519# 0.075021f
C1427 a_21363_45546# VDD 0.36538f
C1428 a_1307_43914# a_11827_44484# 0.025083f
C1429 a_n1059_45260# a_14539_43914# 0.029964f
C1430 a_n2293_42834# a_n2661_43370# 0.038946f
C1431 a_3537_45260# a_n699_43396# 0.025655f
C1432 a_n2312_39304# a_n2661_45546# 0.022905f
C1433 a_12891_46348# a_12839_46116# 0.038804f
C1434 a_19692_46634# a_20202_43084# 0.172738f
C1435 a_19466_46812# a_11415_45002# 0.037852f
C1436 a_n2661_46098# a_n2956_38680# 0.123968f
C1437 C0_P_btm VDD 1.02806f
C1438 a_18194_34908# VIN_N 0.068773f
C1439 C1_N_btm C8_N_btm 0.129306f
C1440 C0_N_btm C9_N_btm 0.146135f
C1441 C0_dummy_N_btm C10_N_btm 0.749362f
C1442 C4_N_btm C5_N_btm 18.6196f
C1443 C3_N_btm C6_N_btm 0.133742f
C1444 C2_N_btm C7_N_btm 0.138288f
C1445 a_3080_42308# a_2903_42308# 0.154008f
C1446 a_2982_43646# a_1606_42308# 0.021878f
C1447 a_15095_43370# a_15597_42852# 0.071983f
C1448 a_13249_42308# a_8685_43396# 0.03355f
C1449 a_11827_44484# a_18579_44172# 0.045146f
C1450 a_10057_43914# a_n2661_42834# 0.053564f
C1451 a_2711_45572# a_15743_43084# 0.075024f
C1452 a_9482_43914# a_10949_43914# 0.025292f
C1453 a_7920_46348# a_8034_45724# 0.032141f
C1454 a_11415_45002# a_20205_31679# 0.070403f
C1455 a_20916_46384# a_2437_43646# 0.010579f
C1456 a_7499_43940# VDD 0.193884f
C1457 a_5534_30871# a_12563_42308# 0.179331f
C1458 a_1414_42308# a_2675_43914# 0.305556f
C1459 a_n2840_43914# a_n4318_39768# 0.170372f
C1460 a_n1059_45260# a_7871_42858# 0.032582f
C1461 a_7640_43914# a_7499_43940# 0.049504f
C1462 a_453_43940# a_895_43940# 0.420851f
C1463 a_2127_44172# a_2479_44172# 0.168988f
C1464 a_20202_43084# a_21613_42308# 0.07574f
C1465 a_13661_43548# START 0.012406f
C1466 a_21076_30879# a_13258_32519# 0.059077f
C1467 a_1823_45246# a_n1059_45260# 0.021319f
C1468 a_18597_46090# a_20679_44626# 0.025074f
C1469 a_18189_46348# a_18175_45572# 0.018402f
C1470 a_1138_42852# a_n913_45002# 0.032304f
C1471 a_n443_46116# a_1467_44172# 0.031058f
C1472 a_n23_45546# a_n443_42852# 0.039956f
C1473 a_n237_47217# a_9313_45822# 0.063143f
C1474 a_3815_47204# a_4007_47204# 0.224415f
C1475 a_n1151_42308# a_n443_46116# 0.099874f
C1476 a_3785_47178# a_4700_47436# 0.090466f
C1477 a_10991_42826# VDD 0.201891f
C1478 a_5379_42460# a_5932_42308# 0.761308f
C1479 a_n2661_42282# a_6452_43396# 0.011968f
C1480 a_10193_42453# a_17303_42282# 0.028322f
C1481 a_n2956_38216# a_n3565_38502# 0.072968f
C1482 a_4704_46090# VDD 0.225404f
C1483 a_11967_42832# a_4361_42308# 0.012085f
C1484 a_13661_43548# a_18533_43940# 0.046643f
C1485 a_11823_42460# a_n2017_45002# 0.098619f
C1486 a_n1613_43370# a_2959_46660# 0.187029f
C1487 a_4915_47217# a_13607_46688# 0.082884f
C1488 a_9313_45822# a_8270_45546# 0.0271f
C1489 a_5807_45002# a_n743_46660# 0.669712f
C1490 a_10227_46804# a_10150_46912# 0.236747f
C1491 a_20753_42852# VDD 0.193909f
C1492 a_n784_42308# C0_P_btm 0.281635f
C1493 a_n97_42460# a_791_42968# 0.039538f
C1494 en_comp a_7754_40130# 0.011333f
C1495 a_21513_45002# a_21359_45002# 0.289039f
C1496 a_413_45260# a_n2661_43370# 1.31746f
C1497 a_8199_44636# a_9801_43940# 0.048015f
C1498 a_n2661_46098# a_n1423_46090# 0.021984f
C1499 a_n743_46660# a_3699_46348# 0.010053f
C1500 a_11735_46660# a_12156_46660# 0.086708f
C1501 a_14976_45028# a_15368_46634# 0.097092f
C1502 a_n746_45260# a_n863_45724# 0.664707f
C1503 a_n971_45724# a_n452_45724# 0.03667f
C1504 a_12089_42308# a_5534_30871# 0.012295f
C1505 a_13113_42826# a_13460_43230# 0.051162f
C1506 a_19778_44110# VDD 0.469922f
C1507 a_3357_43084# a_3499_42826# 0.134316f
C1508 a_4223_44672# a_5883_43914# 0.967973f
C1509 a_413_45260# a_2998_44172# 0.161528f
C1510 a_n443_42852# a_7287_43370# 0.010578f
C1511 a_9290_44172# a_10835_43094# 0.172486f
C1512 a_5343_44458# a_6298_44484# 0.128602f
C1513 a_n2442_46660# a_n3674_38680# 0.023617f
C1514 a_18597_46090# a_20528_45572# 0.03478f
C1515 a_7920_46348# a_8016_46348# 0.318386f
C1516 a_12741_44636# a_10809_44734# 0.088683f
C1517 a_743_42282# a_11551_42558# 0.014689f
C1518 a_17767_44458# a_17973_43940# 0.012863f
C1519 a_5111_44636# a_9885_43646# 0.010527f
C1520 a_n2661_42834# a_5013_44260# 0.021017f
C1521 a_20640_44752# a_20980_44850# 0.027606f
C1522 a_n2293_42834# a_1568_43370# 0.037512f
C1523 a_9313_45822# DATA[5] 0.055804f
C1524 a_n1435_47204# DATA[2] 0.028258f
C1525 a_15507_47210# VDD 0.441662f
C1526 SMPL_ON_N a_21753_35474# 0.39912f
C1527 a_526_44458# a_5837_42852# 0.057897f
C1528 a_12594_46348# a_13163_45724# 0.053634f
C1529 a_2324_44458# a_10490_45724# 0.015189f
C1530 a_5937_45572# a_9241_45822# 0.010703f
C1531 a_8199_44636# a_10210_45822# 0.012124f
C1532 a_10903_43370# a_13904_45546# 0.081466f
C1533 a_526_44458# a_2711_45572# 0.392618f
C1534 a_11415_45002# a_16147_45260# 0.058206f
C1535 a_3090_45724# a_3065_45002# 0.475346f
C1536 a_n2104_42282# a_n4318_37592# 0.033328f
C1537 a_n4318_39768# a_n4318_39304# 0.042825f
C1538 a_9028_43914# a_9165_43940# 0.126609f
C1539 a_15227_46910# VDD 0.229766f
C1540 a_3905_42865# a_n97_42460# 0.071125f
C1541 a_n1761_44111# a_n1557_42282# 0.018977f
C1542 a_n2293_46634# a_3499_42826# 0.022726f
C1543 a_10193_42453# a_8696_44636# 0.225102f
C1544 a_n2810_45572# a_n2956_37592# 0.048284f
C1545 a_584_46384# a_3080_42308# 0.010326f
C1546 a_12549_44172# a_15493_43396# 0.079226f
C1547 a_1138_42852# a_n2661_44458# 0.026505f
C1548 a_n2293_45546# a_n1059_45260# 0.076047f
C1549 a_2063_45854# a_3877_44458# 0.024649f
C1550 a_n443_46116# a_3177_46902# 0.019328f
C1551 a_19386_47436# a_19321_45002# 0.086877f
C1552 a_10807_43548# a_10835_43094# 0.02952f
C1553 a_14401_32519# a_15743_43084# 0.017308f
C1554 a_9313_44734# a_21195_42852# 0.02195f
C1555 a_2957_45546# VDD 0.192471f
C1556 a_10227_46804# a_13113_42826# 0.159547f
C1557 a_4883_46098# a_9127_43156# 0.011077f
C1558 a_2324_44458# a_6453_43914# 0.010794f
C1559 a_2382_45260# a_2680_45002# 0.023953f
C1560 a_10150_46912# a_10467_46802# 0.102355f
C1561 a_7927_46660# a_6755_46942# 0.036549f
C1562 a_n2946_39866# VDD 0.393552f
C1563 a_n2661_42282# a_n4318_37592# 0.03806f
C1564 a_743_42282# a_10341_42308# 0.020229f
C1565 a_9482_43914# VDD 1.75061f
C1566 a_11827_44484# a_22223_45036# 0.179208f
C1567 a_n2956_38216# a_n4318_39304# 0.023138f
C1568 a_4185_45028# a_13467_32519# 0.033397f
C1569 a_5111_44636# a_n2661_43922# 0.061031f
C1570 a_13249_42308# a_13483_43940# 0.193724f
C1571 a_n2293_42834# a_5883_43914# 0.015714f
C1572 a_20567_45036# a_20193_45348# 0.037561f
C1573 a_15227_44166# a_18819_46122# 0.288885f
C1574 a_n743_46660# a_n755_45592# 0.020454f
C1575 a_n2438_43548# a_n357_42282# 0.026249f
C1576 a_n2293_46634# a_3316_45546# 0.067277f
C1577 a_13678_32519# a_22400_42852# 0.03513f
C1578 a_20159_44458# VDD 0.345429f
C1579 a_5147_45002# a_n97_42460# 0.085495f
C1580 a_n357_42282# a_18083_42858# 0.026806f
C1581 a_n2017_45002# a_2982_43646# 0.023101f
C1582 a_n699_43396# a_2675_43914# 0.015641f
C1583 a_n4318_40392# a_n3674_39768# 0.026429f
C1584 a_16327_47482# a_11691_44458# 0.536141f
C1585 a_19553_46090# a_19443_46116# 0.097745f
C1586 a_18479_47436# a_21005_45260# 0.015257f
C1587 a_4791_45118# a_n699_43396# 0.024838f
C1588 a_6031_43396# VDD 0.47547f
C1589 a_18494_42460# a_743_42282# 0.476713f
C1590 a_n357_42282# a_n1794_35082# 0.086672f
C1591 a_7715_46873# VDD 0.414019f
C1592 a_n755_45592# a_564_42282# 0.036154f
C1593 a_2324_44458# a_6171_45002# 2.73828f
C1594 a_10809_44734# a_413_45260# 0.333257f
C1595 a_3090_45724# a_6298_44484# 0.013998f
C1596 a_5066_45546# a_3357_43084# 0.033559f
C1597 a_13259_45724# a_16147_45260# 0.033344f
C1598 a_16763_47508# a_10227_46804# 0.070681f
C1599 a_16327_47482# a_18479_47436# 0.723416f
C1600 a_n1151_42308# a_n1613_43370# 1.19311f
C1601 a_3160_47472# a_n881_46662# 0.070909f
C1602 a_2063_45854# a_8128_46384# 0.032153f
C1603 a_13070_42354# a_13333_42558# 0.011552f
C1604 a_6123_31319# a_4958_30871# 0.021709f
C1605 COMP_P a_1169_39587# 0.388738f
C1606 a_15493_43396# a_16977_43638# 0.018523f
C1607 a_n97_42460# a_4093_43548# 0.028602f
C1608 a_3065_45002# a_3905_42558# 0.044632f
C1609 a_11967_42832# a_17595_43084# 0.0964f
C1610 a_2324_44458# a_14673_44172# 0.015622f
C1611 a_16327_47482# a_4190_30871# 0.335014f
C1612 a_15227_44166# a_11341_43940# 0.04747f
C1613 a_9290_44172# a_11967_42832# 0.0995f
C1614 a_3090_45724# a_10555_44260# 0.041801f
C1615 a_n2293_46634# a_6197_43396# 0.05355f
C1616 a_21188_45572# a_3357_43084# 0.057919f
C1617 a_n237_47217# a_1823_45246# 0.370766f
C1618 a_n1151_42308# a_n2293_46098# 0.040266f
C1619 a_4883_46098# a_14035_46660# 0.019262f
C1620 a_n1925_46634# a_7411_46660# 0.047823f
C1621 a_18597_46090# a_16388_46812# 0.011997f
C1622 a_4958_30871# EN_VIN_BSTR_P 0.021638f
C1623 a_n4209_38216# a_n4064_37984# 0.19304f
C1624 a_n3565_38216# a_n3420_37984# 0.238595f
C1625 a_n4064_39616# a_n4064_37440# 0.050913f
C1626 a_6123_31319# VCM 0.144585f
C1627 a_10723_42308# VDD 0.223902f
C1628 a_8685_43396# a_9127_43156# 0.01312f
C1629 a_n4318_40392# a_n4315_30879# 0.151169f
C1630 a_20623_45572# VDD 0.200978f
C1631 a_n356_44636# a_14113_42308# 0.019853f
C1632 a_3537_45260# a_4223_44672# 0.1907f
C1633 a_n2017_45002# a_14539_43914# 0.01532f
C1634 a_7229_43940# a_n2661_44458# 0.028622f
C1635 a_14537_43396# a_11691_44458# 0.092307f
C1636 a_n2312_39304# a_n2810_45572# 0.044713f
C1637 C1_P_btm VDD 0.264503f
C1638 EN_VIN_BSTR_P VCM 0.929382f
C1639 EN_VIN_BSTR_N VIN_N 1.41696f
C1640 C3_N_btm C5_N_btm 0.135528f
C1641 C0_N_btm C8_N_btm 0.146541f
C1642 C0_dummy_N_btm C9_N_btm 0.111645f
C1643 C2_N_btm C6_N_btm 0.137206f
C1644 C1_N_btm C7_N_btm 0.128479f
C1645 a_5649_42852# a_22165_42308# 0.077779f
C1646 a_n1809_44850# VDD 0.132538f
C1647 a_16922_45042# a_20512_43084# 0.055985f
C1648 a_20193_45348# a_20679_44626# 0.017743f
C1649 a_n755_45592# a_4361_42308# 0.035265f
C1650 a_1307_43914# a_n2661_42282# 0.042336f
C1651 a_7499_43078# a_10341_43396# 0.061281f
C1652 a_9482_43914# a_10729_43914# 0.047853f
C1653 a_11813_46116# a_10193_42453# 0.02832f
C1654 a_19321_45002# a_3357_43084# 0.030763f
C1655 a_3483_46348# a_10586_45546# 0.099824f
C1656 a_n881_46662# a_413_45260# 0.026808f
C1657 a_6671_43940# VDD 0.227011f
C1658 a_5342_30871# a_5742_30871# 0.031909f
C1659 a_1414_42308# a_895_43940# 0.208524f
C1660 a_13747_46662# VDD 3.70214f
C1661 a_20202_43084# a_21887_42336# 0.082645f
C1662 a_1823_45246# a_n2017_45002# 0.024027f
C1663 a_18597_46090# a_20640_44752# 0.027095f
C1664 a_5066_45546# a_9159_45572# 0.040307f
C1665 a_18189_46348# a_16147_45260# 0.129202f
C1666 a_n356_45724# a_n443_42852# 0.056063f
C1667 a_2063_45854# a_6151_47436# 0.448977f
C1668 a_n1151_42308# a_4791_45118# 1.16458f
C1669 a_3785_47178# a_4007_47204# 0.106797f
C1670 a_3160_47472# a_n443_46116# 0.018382f
C1671 a_10796_42968# VDD 0.270235f
C1672 a_4933_42558# a_4921_42308# 0.012385f
C1673 a_5267_42460# a_5932_42308# 0.026805f
C1674 a_5379_42460# a_6171_42473# 0.110293f
C1675 a_4419_46090# VDD 0.664887f
C1676 a_n356_44636# a_5534_30871# 0.054103f
C1677 a_20512_43084# a_15743_43084# 0.761578f
C1678 a_10193_42453# a_4958_30871# 0.108497f
C1679 a_13661_43548# a_19319_43548# 0.189089f
C1680 a_n443_42852# a_14537_43396# 0.03432f
C1681 a_17478_45572# a_16147_45260# 0.050291f
C1682 a_n1613_43370# a_n1809_43762# 0.012235f
C1683 a_n1613_43370# a_3177_46902# 0.209276f
C1684 a_10227_46804# a_9863_46634# 0.278164f
C1685 a_768_44030# a_2107_46812# 0.087742f
C1686 a_n2946_39866# a_n2946_39072# 0.052227f
C1687 a_n4064_39616# a_n3420_39072# 0.05019f
C1688 a_n3420_39616# a_n4064_39072# 6.32746f
C1689 a_1666_39587# a_1273_38525# 0.277775f
C1690 a_n4315_30879# a_n4209_38502# 0.082287f
C1691 a_n784_42308# C1_P_btm 0.027772f
C1692 a_10341_43396# a_15781_43660# 0.011941f
C1693 a_n97_42460# a_685_42968# 0.034735f
C1694 a_5111_44636# a_5837_45028# 0.019542f
C1695 a_4927_45028# a_5093_45028# 0.143754f
C1696 a_15595_45028# a_16019_45002# 0.017418f
C1697 a_3537_45260# a_n2293_42834# 0.195818f
C1698 a_9482_43914# a_1423_45028# 0.014596f
C1699 a_15227_44166# a_10341_43396# 0.068268f
C1700 a_8746_45002# a_10617_44484# 0.01623f
C1701 a_n743_46660# a_3483_46348# 0.050648f
C1702 a_n2661_46098# a_n1991_46122# 0.025798f
C1703 a_3090_45724# a_15368_46634# 0.440843f
C1704 a_n971_45724# a_n863_45724# 0.199707f
C1705 a_12379_42858# a_5534_30871# 0.128429f
C1706 a_12545_42858# a_13460_43230# 0.118423f
C1707 a_18911_45144# VDD 0.218047f
C1708 a_2711_45572# a_3626_43646# 0.072582f
C1709 a_413_45260# a_2889_44172# 0.127135f
C1710 a_7499_43078# a_n97_42460# 0.212833f
C1711 a_9290_44172# a_10518_42984# 0.04331f
C1712 a_5343_44458# a_5518_44484# 0.054464f
C1713 a_n2956_39768# a_n4318_38216# 0.023554f
C1714 a_n971_45724# a_8191_45002# 0.015833f
C1715 a_16327_47482# a_2437_43646# 0.046662f
C1716 a_4646_46812# a_7227_45028# 0.305597f
C1717 a_20820_30879# a_10809_44734# 0.234047f
C1718 a_n443_46116# a_413_45260# 0.369976f
C1719 a_743_42282# a_5742_30871# 0.02341f
C1720 a_9313_45822# DATA[4] 0.0373f
C1721 a_11599_46634# VDD 5.64965f
C1722 a_n1059_45260# a_17499_43370# 0.385066f
C1723 a_n1435_47204# DATA[1] 0.037154f
C1724 SMPL_ON_N a_19998_34978# 0.01194f
C1725 a_19279_43940# a_18579_44172# 0.372064f
C1726 a_526_44458# a_5193_42852# 0.058324f
C1727 a_2324_44458# a_8746_45002# 0.34917f
C1728 a_5937_45572# a_8697_45822# 0.019555f
C1729 a_10903_43370# a_13527_45546# 0.035694f
C1730 a_12594_46348# a_12791_45546# 0.026771f
C1731 a_3483_46348# a_11136_45572# 0.020129f
C1732 a_768_44030# a_n2661_44458# 0.028401f
C1733 a_n1613_43370# a_4223_44672# 0.022154f
C1734 a_n4318_38216# a_n4318_37592# 0.139499f
C1735 a_n356_44636# a_4190_30871# 0.04771f
C1736 a_n2017_45002# a_19987_42826# 0.142839f
C1737 a_n863_45724# a_n2293_45010# 0.090522f
C1738 a_n2293_46098# a_4223_44672# 0.422068f
C1739 a_12549_44172# a_19328_44172# 0.012953f
C1740 a_n2810_45572# a_n2810_45028# 0.063288f
C1741 a_n443_46116# a_2609_46660# 0.349838f
C1742 a_11453_44696# a_768_44030# 0.031665f
C1743 a_10227_46804# a_20916_46384# 0.013668f
C1744 a_n2109_47186# a_5257_43370# 0.153164f
C1745 a_18597_46090# a_19321_45002# 0.024487f
C1746 a_18479_47436# a_20843_47204# 0.021416f
C1747 a_17303_42282# a_21613_42308# 0.061584f
C1748 a_6547_43396# a_6655_43762# 0.057222f
C1749 a_1848_45724# VDD 0.100884f
C1750 a_21381_43940# a_15743_43084# 0.02274f
C1751 a_2324_44458# a_5663_43940# 0.010841f
C1752 a_10227_46804# a_12545_42858# 0.03565f
C1753 a_15227_44166# a_n97_42460# 0.044664f
C1754 a_13661_43548# a_19095_43396# 0.048302f
C1755 a_12549_44172# a_20749_43396# 0.018798f
C1756 a_n443_42852# a_n356_44636# 0.262144f
C1757 a_n755_45592# a_5891_43370# 0.062112f
C1758 a_2274_45254# a_2680_45002# 0.076507f
C1759 a_10150_46912# a_10428_46928# 0.118759f
C1760 a_9863_46634# a_10467_46802# 0.043587f
C1761 a_8145_46902# a_6755_46942# 0.02566f
C1762 a_n1151_42308# a_6945_45028# 0.024325f
C1763 a_n2293_46634# a_13059_46348# 0.207934f
C1764 a_12549_44172# a_18280_46660# 0.03199f
C1765 a_n3420_39616# VDD 0.569005f
C1766 a_n4064_38528# EN_VIN_BSTR_P 0.032872f
C1767 a_n13_43084# a_133_43172# 0.013377f
C1768 a_18783_43370# a_18817_42826# 0.012757f
C1769 a_13348_45260# VDD 0.083657f
C1770 a_3232_43370# a_10617_44484# 0.020516f
C1771 a_375_42282# a_n356_44636# 0.015238f
C1772 a_5111_44636# a_n2661_42834# 0.04935f
C1773 a_5147_45002# a_n2661_43922# 0.029995f
C1774 a_18494_42460# a_20193_45348# 0.116597f
C1775 a_13507_46334# a_22400_42852# 0.235269f
C1776 a_11453_44696# a_11652_45724# 0.01055f
C1777 a_12816_46660# a_10809_44734# 0.011603f
C1778 a_n743_46660# a_n357_42282# 0.03365f
C1779 a_19615_44636# VDD 0.203841f
C1780 a_3080_42308# a_4958_30871# 0.01856f
C1781 a_n357_42282# a_17701_42308# 0.026888f
C1782 a_n2442_46660# a_n2302_39866# 0.161638f
C1783 a_n4318_40392# a_n4318_39768# 2.73673f
C1784 a_18597_46090# a_18184_42460# 0.020766f
C1785 a_n1613_43370# a_n2293_42834# 0.123758f
C1786 a_18985_46122# a_19443_46116# 0.027606f
C1787 a_1823_45246# a_4099_45572# 0.047087f
C1788 a_5066_45546# a_8049_45260# 0.076918f
C1789 a_4791_45118# a_4223_44672# 0.399086f
C1790 a_3080_42308# VCM 0.148824f
C1791 a_n2293_42282# a_n3674_37592# 0.08084f
C1792 a_18184_42460# a_743_42282# 0.126294f
C1793 a_7411_46660# VDD 0.41059f
C1794 a_n357_42282# a_564_42282# 0.026735f
C1795 a_n863_45724# a_961_42354# 0.038222f
C1796 a_n755_45592# a_n3674_37592# 0.063692f
C1797 a_12861_44030# a_12429_44172# 0.108591f
C1798 a_2324_44458# a_3232_43370# 0.410727f
C1799 a_526_44458# a_n2661_45010# 0.703081f
C1800 a_8049_45260# a_21188_45572# 0.015577f
C1801 a_13747_46662# a_21398_44850# 0.011329f
C1802 a_16763_47508# a_17591_47464# 0.010417f
C1803 a_16023_47582# a_10227_46804# 0.036076f
C1804 a_12861_44030# a_13507_46334# 0.315418f
C1805 a_3160_47472# a_n1613_43370# 0.043254f
C1806 a_2905_45572# a_n881_46662# 0.050468f
C1807 a_13070_42354# a_13249_42558# 0.010303f
C1808 a_n1794_35082# a_n4209_39590# 0.177877f
C1809 a_9803_42558# a_10149_42308# 0.013377f
C1810 a_15493_43396# a_16409_43396# 0.566182f
C1811 a_n97_42460# a_1756_43548# 0.052563f
C1812 en_comp a_6123_31319# 0.028754f
C1813 a_11967_42832# a_16795_42852# 0.061673f
C1814 a_n2293_46634# a_6293_42852# 0.014742f
C1815 a_4185_45028# a_3422_30871# 0.176529f
C1816 a_n2956_38216# a_n4318_40392# 0.027558f
C1817 a_21363_45546# a_3357_43084# 0.061421f
C1818 a_16327_47482# a_765_45546# 0.043622f
C1819 a_2959_46660# a_3067_47026# 0.057222f
C1820 a_n1925_46634# a_5257_43370# 0.01497f
C1821 a_11599_46634# a_20107_46660# 0.266678f
C1822 a_4958_30871# a_n1057_35014# 0.017626f
C1823 a_n3565_38216# a_n3690_38304# 0.247167f
C1824 a_n4209_38216# a_n2946_37984# 0.022779f
C1825 a_10533_42308# VDD 0.216201f
C1826 a_15743_43084# a_5649_42852# 0.024346f
C1827 a_20512_43084# a_20256_43172# 0.047194f
C1828 a_20841_45814# VDD 0.209907f
C1829 a_n2293_43922# a_5932_42308# 0.178011f
C1830 a_3065_45002# a_n699_43396# 0.020711f
C1831 a_13507_46334# a_22223_42860# 0.049534f
C1832 a_n2312_40392# a_n2810_45572# 0.052551f
C1833 a_15227_44166# a_11415_45002# 0.047556f
C1834 a_16388_46812# a_18285_46348# 0.028532f
C1835 a_19321_45002# a_8049_45260# 0.030309f
C1836 C2_P_btm VDD 0.268945f
C1837 EN_VIN_BSTR_P VREF_GND 0.857366f
C1838 a_10890_34112# VIN_N 1.547f
C1839 C2_N_btm C5_N_btm 0.13795f
C1840 C3_N_btm C4_N_btm 9.61674f
C1841 C1_N_btm C6_N_btm 0.127656f
C1842 C0_dummy_N_btm C8_N_btm 0.234177f
C1843 C0_N_btm C7_N_btm 0.140846f
C1844 a_13678_32519# a_22165_42308# 0.018986f
C1845 a_n2012_44484# VDD 0.077632f
C1846 a_20193_45348# a_20640_44752# 0.017592f
C1847 a_n357_42282# a_4361_42308# 0.069224f
C1848 a_8975_43940# a_10617_44484# 0.025058f
C1849 a_9482_43914# a_10405_44172# 0.01085f
C1850 a_n1613_43370# a_413_45260# 0.046335f
C1851 a_4791_45118# a_n2293_42834# 0.046352f
C1852 a_20075_46420# a_20708_46348# 0.017547f
C1853 a_8953_45546# a_5066_45546# 0.191859f
C1854 a_5829_43940# VDD 0.156797f
C1855 a_13661_43548# VDD 3.93017f
C1856 a_742_44458# a_1756_43548# 0.152145f
C1857 a_1467_44172# a_895_43940# 0.017277f
C1858 a_1414_42308# a_2479_44172# 0.110442f
C1859 a_9290_44172# a_9885_42558# 0.021204f
C1860 a_20202_43084# a_21335_42336# 0.227943f
C1861 a_n699_43396# a_458_43396# 0.064001f
C1862 a_n755_45592# a_8292_43218# 0.010247f
C1863 a_n2293_46098# a_413_45260# 0.034414f
C1864 a_11453_44696# a_17517_44484# 0.014468f
C1865 a_17715_44484# a_16147_45260# 0.020415f
C1866 a_18479_47436# a_20679_44626# 0.018117f
C1867 a_10835_43094# VDD 0.43308f
C1868 a_n1151_42308# a_4700_47436# 0.01362f
C1869 a_2905_45572# a_n443_46116# 0.14923f
C1870 a_3785_47178# a_3815_47204# 0.270823f
C1871 a_n1605_47204# a_n1435_47204# 0.110832f
C1872 a_5891_43370# a_10083_42826# 0.016347f
C1873 a_n2956_38216# a_n4209_38502# 0.023653f
C1874 a_4185_45028# VDD 1.65665f
C1875 a_20447_31679# a_14097_32519# 0.05131f
C1876 a_6511_45714# a_6171_45002# 0.012882f
C1877 a_15861_45028# a_16147_45260# 0.146279f
C1878 a_17478_45572# a_17786_45822# 0.017351f
C1879 a_21588_30879# a_22612_30879# 7.53611f
C1880 a_n1613_43370# a_2609_46660# 0.631348f
C1881 a_4915_47217# a_12991_46634# 0.068619f
C1882 a_5807_45002# a_n1925_46634# 0.933976f
C1883 a_5111_44636# a_5093_45028# 0.021262f
C1884 a_4927_45028# a_5009_45028# 0.096132f
C1885 a_11823_42460# a_9313_44734# 0.0934f
C1886 a_7499_43078# a_n2661_43922# 0.087751f
C1887 a_14537_43396# a_16751_45260# 0.011362f
C1888 a_768_44030# a_13925_46122# 0.02161f
C1889 a_4883_46098# a_526_44458# 0.010154f
C1890 a_n743_46660# a_3147_46376# 0.016933f
C1891 a_n2661_46098# a_n1853_46287# 0.019613f
C1892 a_n971_45724# a_n1079_45724# 0.150623f
C1893 a_n746_45260# a_n2293_45546# 0.404324f
C1894 a_3090_45724# a_14976_45028# 0.730613f
C1895 a_6755_46942# a_13059_46348# 0.239671f
C1896 a_n4064_37440# C1_P_btm 0.031032f
C1897 a_22537_39537# a_22629_37990# 0.490939f
C1898 a_13113_42826# a_12895_43230# 0.209641f
C1899 a_12545_42858# a_13635_43156# 0.041762f
C1900 a_18587_45118# VDD 0.085535f
C1901 a_526_44458# a_5649_42852# 0.058712f
C1902 a_413_45260# a_2675_43914# 0.048283f
C1903 a_9290_44172# a_10083_42826# 0.136441f
C1904 a_13059_46348# a_8049_45260# 0.068978f
C1905 a_16327_47482# a_21513_45002# 0.013118f
C1906 a_3483_46348# a_9290_44172# 0.207611f
C1907 a_12741_44636# a_6945_45028# 0.021699f
C1908 a_15227_44166# a_13259_45724# 0.916975f
C1909 a_22591_46660# a_10809_44734# 0.013929f
C1910 a_1847_42826# a_2713_42308# 0.015903f
C1911 a_18817_42826# a_18707_42852# 0.097745f
C1912 a_n2661_42834# a_3905_42865# 0.018962f
C1913 a_11967_42832# a_3422_30871# 0.139082f
C1914 a_14311_47204# RST_Z 0.184572f
C1915 a_14955_47212# VDD 0.301751f
C1916 a_n1435_47204# DATA[0] 0.053257f
C1917 a_526_44458# a_4649_42852# 0.028795f
C1918 a_2324_44458# a_10193_42453# 0.041338f
C1919 a_8199_44636# a_8697_45822# 0.067739f
C1920 a_19321_45002# a_20193_45348# 0.489018f
C1921 a_10903_43370# a_13163_45724# 0.06577f
C1922 a_12594_46348# a_11823_42460# 0.081079f
C1923 a_6755_46942# a_13556_45296# 0.103107f
C1924 a_n2104_42282# a_n3674_38216# 0.155459f
C1925 a_n2472_42282# a_n4318_37592# 0.030006f
C1926 a_13259_45724# a_7174_31319# 0.033027f
C1927 a_n2017_45002# a_19164_43230# 0.048221f
C1928 a_12549_44172# a_18451_43940# 0.013387f
C1929 a_11823_42460# a_15037_45618# 0.099829f
C1930 a_584_46384# a_4235_43370# 0.016368f
C1931 a_n443_46116# a_2443_46660# 0.041057f
C1932 a_11453_44696# a_12549_44172# 0.066205f
C1933 a_n971_45724# a_6540_46812# 0.31827f
C1934 a_12861_44030# a_n743_46660# 0.100542f
C1935 a_19386_47436# a_13747_46662# 0.145228f
C1936 a_18479_47436# a_19594_46812# 0.108004f
C1937 a_6765_43638# a_6655_43762# 0.097745f
C1938 a_6547_43396# a_6452_43396# 0.049827f
C1939 a_20692_30879# VCM 0.035438f
C1940 a_997_45618# VDD 0.12359f
C1941 a_9313_44734# a_20922_43172# 0.011702f
C1942 a_n357_42282# a_5891_43370# 0.304889f
C1943 a_2274_45254# a_2382_45260# 0.130215f
C1944 a_7577_46660# a_6755_46942# 0.035922f
C1945 a_9863_46634# a_10428_46928# 0.042509f
C1946 a_12549_44172# a_17639_46660# 0.129285f
C1947 a_7754_38470# a_8530_39574# 0.143675f
C1948 a_7754_40130# CAL_N 0.050321f
C1949 a_n3690_39616# VDD 0.358567f
C1950 a_n2661_42282# a_n3674_38216# 0.051505f
C1951 a_13159_45002# VDD 0.321035f
C1952 a_21381_43940# a_21195_42852# 0.238789f
C1953 a_11967_42832# a_15803_42450# 0.258862f
C1954 a_526_44458# a_8685_43396# 0.04962f
C1955 a_10193_42453# a_19862_44208# 0.099944f
C1956 w_1575_34786# a_5742_30871# 0.776103f
C1957 a_5147_45002# a_n2661_42834# 0.060392f
C1958 a_4791_45118# a_5379_42460# 0.197725f
C1959 a_18184_42460# a_20193_45348# 0.074414f
C1960 a_n743_46660# a_310_45028# 0.143623f
C1961 a_15227_44166# a_18189_46348# 0.066472f
C1962 a_12465_44636# a_11823_42460# 0.127538f
C1963 a_11967_42832# VDD 2.67441f
C1964 a_13467_32519# a_14097_32519# 0.048755f
C1965 en_comp a_3080_42308# 1.2852f
C1966 a_n699_43396# a_2479_44172# 0.063139f
C1967 a_n2442_46660# a_n4064_39616# 0.224005f
C1968 a_9290_44172# a_n357_42282# 0.138435f
C1969 a_n443_46116# a_949_44458# 0.045448f
C1970 a_9313_44734# a_2982_43646# 0.027994f
C1971 a_18494_42460# a_4190_30871# 0.242908f
C1972 a_5257_43370# VDD 0.922495f
C1973 a_n863_45724# a_1184_42692# 0.563857f
C1974 a_n357_42282# a_n3674_37592# 0.327427f
C1975 a_4185_45028# a_1423_45028# 0.016283f
C1976 a_2711_45572# a_11823_42460# 0.065343f
C1977 a_2324_44458# a_5691_45260# 0.013607f
C1978 a_3090_45724# a_5343_44458# 0.023693f
C1979 a_8049_45260# a_21363_45546# 0.013686f
C1980 a_11415_45002# a_n2661_43370# 0.092334f
C1981 a_16763_47508# a_16588_47582# 0.233657f
C1982 a_16327_47482# a_10227_46804# 0.630403f
C1983 a_2905_45572# a_n1613_43370# 0.044171f
C1984 a_15493_43396# a_16547_43609# 0.022221f
C1985 a_n97_42460# a_1568_43370# 0.074153f
C1986 a_20974_43370# a_2982_43646# 0.051776f
C1987 a_11967_42832# a_16414_43172# 0.058563f
C1988 a_1337_46116# VDD 0.20087f
C1989 a_n913_45002# a_8515_42308# 0.01424f
C1990 a_n2661_45546# a_n2661_44458# 0.032856f
C1991 a_n2293_46634# a_6031_43396# 0.037881f
C1992 a_20623_45572# a_3357_43084# 0.041244f
C1993 a_n971_45724# a_1823_45246# 0.514159f
C1994 a_2905_45572# a_n2293_46098# 0.028964f
C1995 a_768_44030# a_8270_45546# 0.03575f
C1996 a_4915_47217# a_11415_45002# 0.134061f
C1997 a_13507_46334# a_14035_46660# 0.027121f
C1998 a_16327_47482# a_17339_46660# 0.058779f
C1999 a_3177_46902# a_3067_47026# 0.097745f
C2000 a_3699_46634# a_3524_46660# 0.233657f
C2001 a_2959_46660# a_2864_46660# 0.049827f
C2002 a_n2109_47186# a_3483_46348# 0.03221f
C2003 a_n4209_38216# a_n3420_37984# 0.067687f
C2004 a_n4064_39616# a_n3420_37440# 0.056826f
C2005 a_n3420_39616# a_n4064_37440# 0.047863f
C2006 a_15743_43084# a_13678_32519# 0.020598f
C2007 a_20273_45572# VDD 0.571099f
C2008 a_5205_44484# a_n2661_44458# 0.072981f
C2009 a_n357_42282# a_10807_43548# 0.031251f
C2010 a_n443_42852# a_3499_42826# 0.023367f
C2011 a_13507_46334# a_22165_42308# 0.126777f
C2012 a_2063_45854# a_7499_43078# 0.478913f
C2013 a_9313_45822# a_2711_45572# 0.016843f
C2014 a_4646_46812# a_2324_44458# 0.023652f
C2015 a_15227_44166# a_20202_43084# 0.086371f
C2016 C3_P_btm VDD 0.26836f
C2017 C2_N_btm C4_N_btm 7.72909f
C2018 C1_N_btm C5_N_btm 0.127408f
C2019 C0_N_btm C6_N_btm 0.139059f
C2020 C0_dummy_N_btm C7_N_btm 0.119061f
C2021 a_18989_43940# VDD 0.342796f
C2022 a_13678_32519# a_21671_42860# 0.014189f
C2023 a_20193_45348# a_20362_44736# 0.013057f
C2024 a_11827_44484# a_19279_43940# 0.078733f
C2025 a_10057_43914# a_10617_44484# 0.033364f
C2026 a_14539_43914# a_9313_44734# 0.016028f
C2027 a_9482_43914# a_9672_43914# 0.122568f
C2028 a_4883_46098# a_8953_45002# 0.013985f
C2029 a_20075_46420# a_19900_46494# 0.233657f
C2030 a_5937_45572# a_5066_45546# 0.419426f
C2031 a_10227_46804# a_14537_43396# 0.094463f
C2032 a_5745_43940# VDD 0.144352f
C2033 a_5534_30871# a_5742_30871# 0.069311f
C2034 a_5807_45002# VDD 1.75047f
C2035 a_742_44458# a_1568_43370# 0.525694f
C2036 a_1115_44172# a_895_43940# 0.029554f
C2037 a_1414_42308# a_2127_44172# 0.091064f
C2038 a_n1925_42282# a_n1794_35082# 0.049072f
C2039 a_20820_30879# a_13258_32519# 0.056725f
C2040 a_n699_43396# a_n229_43646# 0.043893f
C2041 a_18479_47436# a_20640_44752# 0.018112f
C2042 a_16327_47482# a_18579_44172# 0.043297f
C2043 a_10518_42984# VDD 0.273357f
C2044 SMPL_ON_P a_n1435_47204# 0.082028f
C2045 a_n237_47217# a_9067_47204# 0.0235f
C2046 a_n1151_42308# a_4007_47204# 0.015013f
C2047 a_3381_47502# a_3815_47204# 0.021997f
C2048 a_5267_42460# a_5755_42308# 0.055455f
C2049 a_5891_43370# a_8952_43230# 0.016573f
C2050 a_3699_46348# VDD 0.208984f
C2051 a_n2810_45572# a_n3565_38502# 0.409424f
C2052 a_8696_44636# a_16147_45260# 0.284694f
C2053 a_n1613_43370# a_2443_46660# 0.917984f
C2054 a_n881_46662# a_n2661_46098# 0.096736f
C2055 a_n3420_39616# a_n3420_39072# 0.115485f
C2056 a_n4064_39616# a_n3565_39304# 0.028003f
C2057 a_14097_32519# RST_Z 0.051182f
C2058 a_n3565_39590# a_n4064_39072# 0.033734f
C2059 a_15143_45578# VDD 0.12071f
C2060 a_3626_43646# a_5649_42852# 0.032897f
C2061 a_7499_43078# a_n2661_42834# 0.089963f
C2062 a_15415_45028# a_15595_45028# 0.185422f
C2063 a_14537_43396# a_1307_43914# 0.0516f
C2064 a_n467_45028# a_n2661_43370# 0.016799f
C2065 a_3065_45002# a_n2293_42834# 0.021132f
C2066 a_768_44030# a_13759_46122# 0.024686f
C2067 a_4915_47217# a_13259_45724# 0.04489f
C2068 a_n743_46660# a_2804_46116# 0.012952f
C2069 a_n971_45724# a_n2293_45546# 0.097168f
C2070 a_15009_46634# a_14976_45028# 0.071873f
C2071 a_n2661_46098# a_n2157_46122# 0.227082f
C2072 a_n3420_37440# C0_P_btm 0.033333f
C2073 a_7754_38968# VDD 0.041093f
C2074 a_12545_42858# a_12895_43230# 0.215953f
C2075 a_12379_42858# a_13460_43230# 0.102325f
C2076 a_18315_45260# VDD 0.12623f
C2077 a_n2661_43370# a_n2661_43922# 0.13591f
C2078 a_n2956_39768# a_n3674_38680# 0.023454f
C2079 w_1575_34786# a_n4064_39616# 0.03159f
C2080 a_18597_46090# a_20623_45572# 0.046479f
C2081 a_n881_46662# a_16020_45572# 0.013745f
C2082 a_11415_45002# a_10809_44734# 0.140489f
C2083 a_4190_30871# a_5742_30871# 0.029789f
C2084 a_18249_42858# a_18707_42852# 0.027606f
C2085 a_11967_42832# a_21398_44850# 0.01381f
C2086 a_n2661_42834# a_3600_43914# 0.012088f
C2087 a_13487_47204# RST_Z 0.07884f
C2088 a_13717_47436# SINGLE_ENDED 0.032092f
C2089 a_14311_47204# VDD 0.241476f
C2090 a_2324_44458# a_10180_45724# 0.064932f
C2091 a_9290_44172# a_13249_42308# 0.033421f
C2092 a_19321_45002# a_11691_44458# 0.064467f
C2093 a_12594_46348# a_12427_45724# 0.040872f
C2094 a_6755_46942# a_9482_43914# 0.01168f
C2095 a_5257_43370# a_1423_45028# 0.020778f
C2096 a_12465_44636# a_14539_43914# 0.054102f
C2097 a_12005_46116# a_11823_42460# 0.010777f
C2098 a_10903_43370# a_12791_45546# 0.042213f
C2099 a_17364_32525# EN_VIN_BSTR_N 1.00237f
C2100 a_16867_43762# VDD 0.132317f
C2101 a_n4318_38216# a_n3674_38216# 2.91597f
C2102 a_n3674_38680# a_n4318_37592# 0.084223f
C2103 a_n2956_38680# a_n2302_38778# 0.038021f
C2104 a_n2017_45002# a_19339_43156# 0.028127f
C2105 a_19862_44208# a_14021_43940# 0.021104f
C2106 a_n863_45724# a_n2661_45010# 0.345234f
C2107 a_n443_46116# a_n97_42460# 0.131756f
C2108 a_12549_44172# a_18326_43940# 0.013334f
C2109 a_11823_42460# a_14033_45822# 0.093809f
C2110 a_9049_44484# a_8696_44636# 0.043734f
C2111 a_n2293_45546# a_n2293_45010# 0.257189f
C2112 a_11453_44696# a_12891_46348# 0.029995f
C2113 a_10227_46804# a_20843_47204# 0.02328f
C2114 a_n443_46116# a_n2661_46098# 0.198865f
C2115 a_18597_46090# a_13747_46662# 0.391702f
C2116 a_18479_47436# a_19321_45002# 0.262984f
C2117 a_19332_42282# a_19647_42308# 0.084365f
C2118 a_n2293_42282# VDD 0.464485f
C2119 a_6197_43396# a_6655_43762# 0.027317f
C2120 a_20193_45348# a_20753_42852# 0.04748f
C2121 a_20205_31679# VCM 0.035399f
C2122 a_20692_30879# VREF_GND 0.010456f
C2123 a_n755_45592# VDD 2.41485f
C2124 a_10227_46804# a_12379_42858# 0.298444f
C2125 a_13059_46348# a_13565_43940# 0.011241f
C2126 a_413_45260# a_3065_45002# 0.027891f
C2127 a_2711_45572# a_14539_43914# 0.199754f
C2128 a_n1613_43370# a_n1076_43230# 0.224215f
C2129 a_7715_46873# a_6755_46942# 0.089466f
C2130 a_9863_46634# a_10150_46912# 0.233657f
C2131 a_7411_46660# a_6969_46634# 0.033891f
C2132 a_13747_46662# a_19123_46287# 0.191545f
C2133 a_n881_46662# a_11415_45002# 0.017774f
C2134 a_12861_44030# a_9290_44172# 0.09212f
C2135 a_7754_40130# a_11206_38545# 0.736866f
C2136 a_n3565_39590# VDD 1.32666f
C2137 a_n3420_38528# EN_VIN_BSTR_P 0.031989f
C2138 a_13017_45260# VDD 0.263701f
C2139 a_21381_43940# a_21356_42826# 0.196864f
C2140 a_11967_42832# a_15764_42576# 0.012941f
C2141 a_n2810_45572# a_n4318_39304# 0.023142f
C2142 a_1307_43914# a_n356_44636# 0.013327f
C2143 a_4791_45118# a_5267_42460# 0.138738f
C2144 a_19778_44110# a_20193_45348# 0.020562f
C2145 a_n743_46660# a_n1099_45572# 0.108295f
C2146 a_15227_44166# a_17715_44484# 0.385336f
C2147 a_12251_46660# a_10809_44734# 0.023146f
C2148 a_19006_44850# VDD 0.077608f
C2149 a_19237_31679# EN_VIN_BSTR_N 0.095737f
C2150 a_13467_32519# a_22400_42852# 0.029863f
C2151 a_7227_42852# a_7309_42852# 0.171361f
C2152 a_n357_42282# a_16795_42852# 0.180926f
C2153 a_n913_45002# a_n1557_42282# 0.015193f
C2154 a_3537_45260# a_n97_42460# 0.74108f
C2155 a_n2661_42834# a_12189_44484# 0.010003f
C2156 a_n2312_38680# a_n3565_39590# 0.031736f
C2157 a_n2442_46660# a_n2946_39866# 0.024649f
C2158 a_n443_46116# a_742_44458# 0.018829f
C2159 a_15227_44166# a_15861_45028# 0.208121f
C2160 a_1823_45246# a_2711_45572# 0.262616f
C2161 a_n2293_42282# a_n784_42308# 0.055588f
C2162 a_n755_45592# a_n784_42308# 0.711298f
C2163 a_18184_42460# a_4190_30871# 0.630738f
C2164 a_n863_45724# a_1576_42282# 0.05148f
C2165 a_2711_45572# a_12427_45724# 0.014959f
C2166 a_3090_45724# a_4743_44484# 0.05313f
C2167 a_8049_45260# a_20623_45572# 0.01128f
C2168 a_13059_46348# a_11691_44458# 0.015799f
C2169 a_11599_46634# a_18597_46090# 0.191253f
C2170 a_16241_47178# a_10227_46804# 0.022072f
C2171 a_16327_47482# a_17591_47464# 0.339529f
C2172 a_11967_42832# a_15567_42826# 0.067391f
C2173 a_15493_43396# a_16243_43396# 0.041358f
C2174 a_n97_42460# a_1049_43396# 0.195034f
C2175 a_17973_43940# a_17499_43370# 0.018568f
C2176 a_n913_45002# a_5934_30871# 0.126791f
C2177 a_10809_44734# a_n2661_43922# 0.073946f
C2178 a_19692_46634# a_19862_44208# 0.027038f
C2179 a_13507_46334# a_15743_43084# 0.158635f
C2180 a_2711_45572# a_14309_45028# 0.028068f
C2181 a_20841_45814# a_3357_43084# 0.047766f
C2182 a_2609_46660# a_3067_47026# 0.027317f
C2183 a_13747_46662# a_6755_46942# 0.316914f
C2184 a_15673_47210# a_765_45546# 0.028544f
C2185 a_11599_46634# a_19123_46287# 0.024241f
C2186 a_6123_31319# VIN_N 0.01057f
C2187 a_5742_30871# C7_N_btm 0.04157f
C2188 a_2112_39137# VDAC_Pi 0.01062f
C2189 a_n4209_38216# a_n3690_38304# 0.045342f
C2190 a_9885_42558# VDD 0.18767f
C2191 a_20107_45572# VDD 0.458237f
C2192 a_3422_30871# a_14097_32519# 0.031284f
C2193 a_13556_45296# a_11691_44458# 0.399095f
C2194 a_2382_45260# a_n699_43396# 0.075387f
C2195 a_16388_46812# a_765_45546# 0.164902f
C2196 a_6151_47436# a_6598_45938# 0.173467f
C2197 a_7927_46660# a_8349_46414# 0.01072f
C2198 a_n881_46662# a_13259_45724# 0.507296f
C2199 a_3877_44458# a_2324_44458# 0.153319f
C2200 a_13747_46662# a_8049_45260# 0.208778f
C2201 a_n743_46660# a_n1925_42282# 0.010043f
C2202 a_n2438_43548# a_526_44458# 0.107408f
C2203 C4_P_btm VDD 0.265463f
C2204 C1_N_btm C4_N_btm 0.128167f
C2205 C0_N_btm C5_N_btm 0.138093f
C2206 C2_N_btm C3_N_btm 5.99608f
C2207 C0_dummy_N_btm C6_N_btm 0.1194f
C2208 a_18374_44850# VDD 0.203584f
C2209 a_5883_43914# a_n2661_43922# 0.028328f
C2210 a_10440_44484# a_10617_44484# 0.134298f
C2211 a_9482_43914# a_9028_43914# 0.092045f
C2212 a_n2293_42834# a_2479_44172# 0.021799f
C2213 a_2063_45854# a_n2661_43370# 0.039988f
C2214 a_13059_46348# a_n443_42852# 0.09278f
C2215 a_8199_44636# a_5066_45546# 0.178583f
C2216 a_1414_42308# a_453_43940# 0.248504f
C2217 a_644_44056# a_895_43940# 0.106452f
C2218 a_16131_47204# VDD 0.142103f
C2219 a_20202_43084# a_20712_42282# 0.028679f
C2220 a_11309_47204# CLK 0.01087f
C2221 a_380_45546# a_603_45572# 0.011458f
C2222 a_4185_45028# a_3357_43084# 0.027077f
C2223 a_2063_45854# a_4915_47217# 0.055521f
C2224 a_n237_47217# a_6575_47204# 0.0275f
C2225 a_n1151_42308# a_3815_47204# 0.01223f
C2226 a_n1741_47186# a_n1435_47204# 0.047534f
C2227 a_10083_42826# VDD 0.461256f
C2228 COMP_P a_5742_30871# 0.109332f
C2229 a_5267_42460# a_5421_42558# 0.010303f
C2230 a_3483_46348# VDD 2.29096f
C2231 a_19963_31679# a_14097_32519# 0.051059f
C2232 a_5891_43370# a_9127_43156# 0.457718f
C2233 a_n1059_45260# a_16877_42852# 0.058551f
C2234 a_n1613_43370# a_n97_42460# 0.011527f
C2235 a_n755_45592# a_1423_45028# 0.032517f
C2236 a_11599_46634# a_6755_46942# 0.321942f
C2237 a_13661_43548# a_n2293_46634# 0.055067f
C2238 a_n881_46662# a_1799_45572# 0.028083f
C2239 a_n1613_43370# a_n2661_46098# 1.40554f
C2240 a_1606_42308# EN_VIN_BSTR_N 0.035204f
C2241 a_n3420_39616# a_n3690_39392# 0.018295f
C2242 a_22400_42852# RST_Z 0.059672f
C2243 a_5934_30871# VDAC_P 0.029185f
C2244 a_14097_32519# VDD 0.285619f
C2245 a_10490_45724# CLK 0.029352f
C2246 a_14495_45572# VDD 0.238674f
C2247 a_9049_44484# a_9159_44484# 0.031707f
C2248 a_15227_44166# a_15095_43370# 0.022423f
C2249 a_3090_45724# a_12281_43396# 0.027472f
C2250 a_n357_42282# a_3422_30871# 0.122733f
C2251 a_n2293_46098# a_n97_42460# 0.333817f
C2252 a_n2293_46634# a_4185_45028# 0.027799f
C2253 a_n2497_47436# a_n755_45592# 0.45034f
C2254 a_n237_47217# a_n2661_45546# 0.038356f
C2255 a_11599_46634# a_8049_45260# 0.14064f
C2256 a_n743_46660# a_2698_46116# 0.013101f
C2257 a_15009_46634# a_3090_45724# 0.154981f
C2258 a_n2661_46098# a_n2293_46098# 0.063852f
C2259 a_22527_39145# a_22737_36887# 0.011525f
C2260 a_22537_39537# a_22629_38406# 0.198762f
C2261 a_12545_42858# a_13113_42826# 0.178024f
C2262 a_12379_42858# a_13635_43156# 0.043475f
C2263 a_17719_45144# VDD 0.1297f
C2264 a_n1925_42282# a_4361_42308# 0.08654f
C2265 a_n2661_43370# a_n2661_42834# 0.306215f
C2266 a_n443_42852# a_6293_42852# 0.033407f
C2267 a_4185_45028# a_5342_30871# 0.067871f
C2268 a_18597_46090# a_20841_45814# 0.024341f
C2269 a_n881_46662# a_17478_45572# 0.11503f
C2270 a_4646_46812# a_6511_45714# 0.421269f
C2271 a_20202_43084# a_10809_44734# 0.014133f
C2272 a_11415_45002# a_22223_46124# 0.011454f
C2273 a_743_42282# a_10533_42308# 0.016446f
C2274 a_4361_42308# a_9803_42558# 0.011987f
C2275 a_14539_43914# a_15682_43940# 0.161926f
C2276 a_n2661_42834# a_2998_44172# 0.790177f
C2277 a_13487_47204# VDD 0.273369f
C2278 a_9067_47204# DATA[4] 0.354356f
C2279 a_13717_47436# START 0.034426f
C2280 a_12861_44030# RST_Z 0.290405f
C2281 a_19321_45002# a_19113_45348# 0.147788f
C2282 a_13747_46662# a_20193_45348# 0.049365f
C2283 a_12594_46348# a_11962_45724# 0.177228f
C2284 a_n443_46116# a_n2661_43922# 0.044169f
C2285 a_10903_43370# a_11823_42460# 1.16382f
C2286 a_12005_46116# a_12427_45724# 0.01091f
C2287 a_16664_43396# VDD 0.077608f
C2288 a_n2840_42282# a_n4318_37592# 0.037154f
C2289 a_n2472_42282# a_n3674_38216# 0.040147f
C2290 a_n2956_38680# a_n4064_38528# 0.058755f
C2291 a_14513_46634# VDD 0.223375f
C2292 a_11341_43940# a_11173_44260# 0.049235f
C2293 a_n2017_45002# a_18599_43230# 0.029677f
C2294 a_20512_43084# a_2982_43646# 0.029475f
C2295 a_4791_45118# a_n97_42460# 0.02536f
C2296 a_12861_44030# a_19319_43548# 0.024237f
C2297 a_7499_43078# a_8696_44636# 0.155392f
C2298 a_10210_45822# a_10907_45822# 0.013775f
C2299 a_10227_46804# a_19594_46812# 0.01518f
C2300 a_n443_46116# a_1799_45572# 0.081828f
C2301 a_18597_46090# a_13661_43548# 0.266647f
C2302 a_18780_47178# a_13747_46662# 0.028845f
C2303 a_19332_42282# a_19511_42282# 0.174683f
C2304 a_22959_42860# VDD 0.30747f
C2305 a_17303_42282# a_7174_31319# 0.027048f
C2306 a_6197_43396# a_6452_43396# 0.06121f
C2307 a_n357_42282# VDD 1.90108f
C2308 a_20692_30879# VREF 0.098117f
C2309 a_13661_43548# a_743_42282# 0.132115f
C2310 a_413_45260# a_2680_45002# 0.01804f
C2311 a_2711_45572# a_16112_44458# 0.183744f
C2312 a_n1613_43370# a_n901_43156# 0.281398f
C2313 a_2063_45854# a_10809_44734# 0.169005f
C2314 a_7411_46660# a_6755_46942# 0.265786f
C2315 a_13661_43548# a_19123_46287# 0.073049f
C2316 a_3754_38470# a_8530_39574# 0.059662f
C2317 a_7754_40130# VDAC_P 0.334598f
C2318 VDAC_Pi a_6886_37412# 0.259481f
C2319 a_n4334_39616# VDD 0.385881f
C2320 a_6171_45002# CLK 0.032376f
C2321 a_11963_45334# VDD 0.229584f
C2322 a_n2661_42282# a_n4318_38216# 0.023731f
C2323 a_3232_43370# a_3363_44484# 0.103472f
C2324 a_3537_45260# a_n2661_43922# 0.058875f
C2325 a_21101_45002# a_21359_45002# 0.22264f
C2326 a_4185_45028# a_743_42282# 0.031243f
C2327 a_10193_42453# a_15493_43396# 0.024143f
C2328 a_19778_44110# a_11691_44458# 0.013164f
C2329 a_n743_46660# a_380_45546# 0.010247f
C2330 a_12469_46902# a_10809_44734# 0.014309f
C2331 a_18588_44850# VDD 0.132317f
C2332 a_8387_43230# a_8483_43230# 0.013793f
C2333 a_n1059_45260# a_n1557_42282# 0.031252f
C2334 a_n2956_39768# a_n2302_39866# 0.037924f
C2335 a_2107_46812# a_6171_45002# 0.023061f
C2336 a_5257_43370# a_3357_43084# 0.894879f
C2337 a_18479_47436# a_19778_44110# 0.038618f
C2338 a_15227_44166# a_8696_44636# 0.203885f
C2339 a_16327_47482# a_11827_44484# 0.107078f
C2340 a_3080_42308# VIN_N 0.025929f
C2341 a_n755_45592# a_196_42282# 0.090568f
C2342 a_n863_45724# a_1067_42314# 0.289393f
C2343 a_2324_44458# a_5111_44636# 0.090721f
C2344 a_3483_46348# a_1423_45028# 0.110369f
C2345 a_9290_44172# a_10951_45334# 0.136064f
C2346 a_2711_45572# a_11962_45724# 0.054424f
C2347 a_3090_45724# a_n699_43396# 0.058797f
C2348 a_n1613_43370# a_n984_44318# 0.245331f
C2349 a_9313_45822# a_4883_46098# 0.026043f
C2350 a_16327_47482# a_16588_47582# 0.276601f
C2351 a_15673_47210# a_10227_46804# 0.02634f
C2352 a_n443_46116# a_2747_46873# 0.047485f
C2353 a_2063_45854# a_n881_46662# 0.612456f
C2354 a_n971_45724# a_768_44030# 0.069358f
C2355 a_11967_42832# a_5342_30871# 0.077151f
C2356 a_15493_43396# a_16137_43396# 0.023247f
C2357 a_n97_42460# a_1209_43370# 0.027601f
C2358 a_104_43370# a_458_43396# 0.07022f
C2359 a_21381_43940# a_2982_43646# 0.236232f
C2360 a_17737_43940# a_17499_43370# 0.013048f
C2361 a_n1059_45260# a_5934_30871# 0.010576f
C2362 a_n913_45002# a_7963_42308# 0.044607f
C2363 a_10809_44734# a_n2661_42834# 0.14417f
C2364 a_n2810_45572# a_n4318_40392# 0.02461f
C2365 a_20273_45572# a_3357_43084# 0.358383f
C2366 a_15903_45785# a_6171_45002# 0.011492f
C2367 a_2107_46812# a_4955_46873# 0.031068f
C2368 a_2609_46660# a_2864_46660# 0.055869f
C2369 a_3177_46902# a_3524_46660# 0.051162f
C2370 a_n2661_46634# a_7577_46660# 0.047111f
C2371 a_13661_43548# a_6755_46942# 0.088986f
C2372 a_n2293_46634# a_5257_43370# 0.061974f
C2373 a_15811_47375# a_765_45546# 0.035109f
C2374 a_11599_46634# a_18285_46348# 0.030958f
C2375 a_n3565_39590# a_n4064_37440# 0.031724f
C2376 a_6123_31319# VIN_P 0.01057f
C2377 a_5742_30871# C6_N_btm 0.170624f
C2378 a_n4209_38216# a_n3565_38216# 6.80743f
C2379 a_n4064_39616# a_n3565_37414# 0.028438f
C2380 a_n3420_39616# a_n3420_37440# 0.053603f
C2381 a_15743_43084# a_4361_42308# 0.020459f
C2382 a_3422_30871# a_22400_42852# 0.023064f
C2383 a_14537_43396# a_11827_44484# 0.076354f
C2384 a_9482_43914# a_11691_44458# 0.616964f
C2385 a_5937_45572# a_6031_43396# 0.010894f
C2386 a_16388_46812# a_17339_46660# 0.24887f
C2387 a_6151_47436# a_6667_45809# 0.1609f
C2388 a_12891_46348# a_12638_46436# 0.13727f
C2389 a_n743_46660# a_526_44458# 0.020498f
C2390 a_13661_43548# a_8049_45260# 0.032643f
C2391 EN_VIN_BSTR_P VIN_P 1.41696f
C2392 C5_P_btm VDD 0.267489f
C2393 C0_N_btm C4_N_btm 0.138331f
C2394 C0_dummy_N_btm C5_N_btm 0.11375f
C2395 C1_N_btm C3_N_btm 8.06688f
C2396 a_18443_44721# VDD 0.193515f
C2397 a_4361_42308# a_21671_42860# 0.012186f
C2398 a_5883_43914# a_n2661_42834# 0.106812f
C2399 a_1307_43914# a_3499_42826# 0.532672f
C2400 a_11823_42460# a_8685_43396# 0.057344f
C2401 a_768_44030# a_n2293_45010# 0.03517f
C2402 a_584_46384# a_n2661_43370# 0.034714f
C2403 a_5807_45002# a_3357_43084# 0.071743f
C2404 a_11453_44696# a_6171_45002# 1.39146f
C2405 a_19553_46090# a_19900_46494# 0.051162f
C2406 a_4185_45028# a_8049_45260# 0.014062f
C2407 a_1467_44172# a_453_43940# 0.05905f
C2408 a_9290_44172# a_9803_42558# 0.094028f
C2409 a_n1925_42282# a_n3674_37592# 0.072052f
C2410 a_12861_44030# a_3422_30871# 0.018986f
C2411 a_768_44030# a_9313_44734# 0.044729f
C2412 a_380_45546# a_509_45572# 0.010132f
C2413 a_584_46384# a_2998_44172# 0.181241f
C2414 a_4185_45028# a_19479_31679# 0.03554f
C2415 a_1848_45724# a_1609_45822# 0.042695f
C2416 a_n1613_43370# a_n2661_43922# 0.113996f
C2417 a_18597_46090# a_11967_42832# 0.021692f
C2418 a_n237_47217# a_7903_47542# 0.086772f
C2419 a_n1151_42308# a_3785_47178# 0.029415f
C2420 a_2063_45854# a_n443_46116# 0.177177f
C2421 a_8952_43230# VDD 0.273404f
C2422 a_5379_42460# a_4921_42308# 0.033756f
C2423 a_5267_42460# a_5337_42558# 0.011552f
C2424 a_1606_42308# a_5934_30871# 0.095492f
C2425 a_3147_46376# VDD 0.341038f
C2426 a_11967_42832# a_743_42282# 0.043946f
C2427 a_5891_43370# a_8387_43230# 0.010767f
C2428 a_n1059_45260# a_16245_42852# 0.130348f
C2429 a_n2810_45572# a_n4209_38502# 0.066112f
C2430 a_13507_46334# a_3626_43646# 0.04477f
C2431 a_n2293_46098# a_n2661_43922# 0.026124f
C2432 a_n3420_39616# a_n3565_39304# 0.035199f
C2433 a_1169_39587# a_1666_39587# 0.105143f
C2434 a_n3690_39616# a_n3690_39392# 0.052468f
C2435 a_n3565_39590# a_n3420_39072# 0.033891f
C2436 a_n4209_39590# a_n4064_39072# 0.03458f
C2437 a_n4064_39616# a_n4209_39304# 0.029393f
C2438 a_22400_42852# VDD 0.888056f
C2439 a_3539_42460# a_4361_42308# 0.027414f
C2440 a_2982_43646# a_5649_42852# 0.205161f
C2441 a_20512_43084# a_19987_42826# 0.11919f
C2442 a_8746_45002# CLK 0.018523f
C2443 a_13249_42308# VDD 0.653917f
C2444 a_4558_45348# a_5009_45028# 0.013349f
C2445 a_5937_45572# a_6671_43940# 0.06027f
C2446 a_2382_45260# a_n2293_42834# 0.026697f
C2447 a_n881_46662# a_17715_44484# 0.014166f
C2448 a_n2497_47436# a_n357_42282# 0.046314f
C2449 a_n746_45260# a_n2661_45546# 0.022378f
C2450 a_12549_44172# a_13351_46090# 0.014836f
C2451 a_n743_46660# a_2521_46116# 0.013075f
C2452 a_n2438_43548# a_167_45260# 0.050543f
C2453 a_1799_45572# a_n2293_46098# 0.014011f
C2454 a_n2661_46098# a_n2472_46090# 0.094589f
C2455 a_n3565_37414# C0_P_btm 0.040442f
C2456 a_22581_37893# a_22629_37990# 0.333805f
C2457 a_22527_39145# a_22737_37285# 0.012249f
C2458 a_22537_39537# CAL_P 0.024815f
C2459 VDAC_N EN_VIN_BSTR_N 0.341739f
C2460 a_12379_42858# a_12895_43230# 0.109156f
C2461 a_17613_45144# VDD 0.094022f
C2462 a_4223_44672# a_5343_44458# 0.229803f
C2463 a_526_44458# a_4361_42308# 0.072573f
C2464 a_413_45260# a_2127_44172# 0.104737f
C2465 a_n443_42852# a_6031_43396# 0.020526f
C2466 a_n699_43396# a_4743_44484# 0.235328f
C2467 a_18479_45785# a_15493_43396# 0.235084f
C2468 w_1575_34786# a_n3420_39616# 0.039343f
C2469 a_18597_46090# a_20273_45572# 0.048762f
C2470 a_15507_47210# a_2437_43646# 0.027848f
C2471 a_n881_46662# a_15861_45028# 0.153795f
C2472 a_4646_46812# a_6472_45840# 0.129446f
C2473 a_22365_46825# a_10809_44734# 0.010841f
C2474 a_2107_46812# a_8746_45002# 0.020783f
C2475 a_n1441_43940# VDD 0.142719f
C2476 a_12861_44030# VDD 3.56689f
C2477 a_6575_47204# DATA[4] 0.15718f
C2478 a_17517_44484# a_22591_44484# 0.196232f
C2479 a_14539_43914# a_14955_43940# 0.064683f
C2480 a_13717_47436# RST_Z 4.51263f
C2481 a_n1059_45260# a_16547_43609# 0.024317f
C2482 a_626_44172# a_648_43396# 0.04847f
C2483 a_20766_44850# a_19279_43940# 0.021466f
C2484 a_16375_45002# a_18051_46116# 0.038793f
C2485 a_2324_44458# a_9049_44484# 0.102942f
C2486 a_4791_45118# a_n2661_43922# 0.034957f
C2487 a_n443_46116# a_n2661_42834# 0.075503f
C2488 a_10903_43370# a_12427_45724# 0.083943f
C2489 a_14209_32519# EN_VIN_BSTR_N 0.032872f
C2490 a_19700_43370# VDD 0.28578f
C2491 a_n3674_38680# a_n3674_38216# 0.059687f
C2492 a_15493_43396# a_14021_43940# 0.139192f
C2493 a_n2956_38680# a_n2946_38778# 0.14863f
C2494 a_14180_46812# VDD 0.755623f
C2495 a_13259_45724# a_13258_32519# 0.037974f
C2496 a_3357_43084# a_n2293_42282# 0.146926f
C2497 a_12549_44172# a_17973_43940# 0.015874f
C2498 a_4185_45028# a_20193_45348# 0.015456f
C2499 a_584_46384# a_1568_43370# 0.057089f
C2500 a_n2293_45546# a_n2661_45010# 0.014846f
C2501 a_6755_46942# a_11967_42832# 0.030705f
C2502 a_18780_47178# a_13661_43548# 0.153988f
C2503 a_18479_47436# a_13747_46662# 0.083389f
C2504 a_10227_46804# a_19321_45002# 0.111029f
C2505 a_12465_44636# a_768_44030# 0.120859f
C2506 a_2747_46873# a_n1613_43370# 0.03071f
C2507 a_22223_42860# VDD 0.250812f
C2508 a_4958_30871# a_7174_31319# 0.107892f
C2509 a_7287_43370# a_7112_43396# 0.234322f
C2510 a_6293_42852# a_6452_43396# 0.157972f
C2511 a_19319_43548# a_19268_43646# 0.17076f
C2512 a_20205_31679# VREF 0.056031f
C2513 a_310_45028# VDD 0.360949f
C2514 a_9313_44734# a_19339_43156# 0.01152f
C2515 a_20692_30879# VIN_N 0.038535f
C2516 a_8746_45002# a_n2661_44458# 0.017636f
C2517 a_10227_46804# a_10922_42852# 0.159426f
C2518 a_13661_43548# a_20301_43646# 0.072262f
C2519 a_413_45260# a_2382_45260# 0.048205f
C2520 a_8696_44636# a_n2661_43370# 0.674122f
C2521 a_n1613_43370# a_n1641_43230# 0.152896f
C2522 a_13661_43548# a_18285_46348# 0.049064f
C2523 VDAC_Pi a_5700_37509# 2.20213f
C2524 a_7174_31319# VCM 0.076834f
C2525 a_7754_39964# a_6886_37412# 0.035115f
C2526 a_7754_40130# a_8912_37509# 1.81084f
C2527 a_n4209_39590# VDD 2.07895f
C2528 a_n2661_42282# a_n2472_42282# 0.028691f
C2529 a_n1641_43230# a_n1533_42852# 0.057222f
C2530 a_18525_43370# a_18083_42858# 0.016073f
C2531 a_11787_45002# VDD 0.153399f
C2532 a_3537_45260# a_n2661_42834# 0.097192f
C2533 a_11823_42460# a_13483_43940# 0.029429f
C2534 a_n2293_42834# a_5343_44458# 0.165923f
C2535 a_18911_45144# a_11691_44458# 0.013593f
C2536 a_4915_47217# a_8696_44636# 0.02426f
C2537 a_768_44030# a_2711_45572# 0.529995f
C2538 a_22959_46660# a_21076_30879# 0.165603f
C2539 a_11901_46660# a_10809_44734# 0.048084f
C2540 a_n2293_46634# a_n755_45592# 0.094759f
C2541 a_n2438_43548# a_n863_45724# 0.07341f
C2542 a_n743_46660# a_n452_45724# 0.070244f
C2543 a_18817_42826# a_19164_43230# 0.051162f
C2544 a_5755_42852# a_5837_42852# 0.171361f
C2545 a_8387_43230# a_8292_43218# 0.049827f
C2546 a_17730_32519# EN_VIN_BSTR_N 0.073198f
C2547 a_n2017_45002# a_n1557_42282# 0.090464f
C2548 a_n2956_39768# a_n4064_39616# 0.058734f
C2549 a_n913_45002# a_4905_42826# 0.101072f
C2550 a_n2312_38680# a_n4209_39590# 0.020921f
C2551 a_1823_45246# a_4649_42852# 0.042816f
C2552 a_742_44458# a_895_43940# 0.025021f
C2553 a_3065_45002# a_n97_42460# 0.019675f
C2554 a_n699_43396# a_1414_42308# 0.104607f
C2555 a_5066_45546# a_8034_45724# 0.242476f
C2556 a_2107_46812# a_3232_43370# 0.026265f
C2557 a_19335_46494# a_19431_46494# 0.013793f
C2558 a_3080_42308# VIN_P 0.025929f
C2559 a_10057_43914# a_10695_43548# 0.148476f
C2560 a_n357_42282# a_196_42282# 0.033292f
C2561 a_n755_45592# a_n473_42460# 0.061354f
C2562 a_9290_44172# a_10775_45002# 0.215292f
C2563 a_2324_44458# a_5147_45002# 0.056065f
C2564 a_2711_45572# a_11652_45724# 0.013232f
C2565 a_8049_45260# a_20273_45572# 0.040989f
C2566 a_3090_45724# a_4223_44672# 0.269823f
C2567 a_n2956_38680# a_n2956_37592# 0.047258f
C2568 a_n1613_43370# a_n809_44244# 0.291484f
C2569 a_8199_44636# a_9482_43914# 0.276776f
C2570 a_16241_47178# a_16588_47582# 0.051162f
C2571 a_15811_47375# a_10227_46804# 0.019973f
C2572 a_2063_45854# a_n1613_43370# 0.04116f
C2573 a_584_46384# a_n881_46662# 0.286501f
C2574 a_16327_47482# a_16763_47508# 0.338544f
C2575 a_n4318_37592# a_n4064_39616# 0.021014f
C2576 a_5932_42308# a_4958_30871# 0.01835f
C2577 a_n97_42460# a_458_43396# 0.013064f
C2578 a_11967_42832# a_15279_43071# 0.027468f
C2579 a_3065_45002# a_3823_42558# 0.198186f
C2580 a_n913_45002# a_6123_31319# 0.21316f
C2581 a_21363_45546# a_21513_45002# 0.06363f
C2582 a_16327_47482# a_16823_43084# 0.535969f
C2583 a_7227_45028# a_n2661_43370# 0.026158f
C2584 a_3090_45724# a_15493_43940# 0.255251f
C2585 a_526_44458# a_5891_43370# 1.12739f
C2586 a_20107_45572# a_3357_43084# 0.308463f
C2587 a_2063_45854# a_n2293_46098# 0.994164f
C2588 a_10227_46804# a_13059_46348# 0.656528f
C2589 a_2609_46660# a_3524_46660# 0.118759f
C2590 a_2443_46660# a_2864_46660# 0.090164f
C2591 a_5807_45002# a_6755_46942# 1.47519f
C2592 a_5932_42308# VCM 0.146001f
C2593 a_5742_30871# C5_N_btm 0.089375f
C2594 a_n4209_38216# a_n4334_38304# 0.253307f
C2595 a_15743_43084# a_13467_32519# 0.02051f
C2596 a_19268_43646# a_19095_43396# 0.032587f
C2597 a_5891_43370# a_9223_42460# 0.13879f
C2598 a_3232_43370# a_n2661_44458# 0.468391f
C2599 a_6151_47436# a_6511_45714# 0.3215f
C2600 a_2063_45854# a_7230_45938# 0.016263f
C2601 a_3090_45724# a_12741_44636# 0.093609f
C2602 a_5807_45002# a_8049_45260# 1.37423f
C2603 a_n1057_35014# VIN_P 1.547f
C2604 C6_P_btm VDD 0.210613f
C2605 C0_dummy_N_btm C4_N_btm 0.113156f
C2606 C1_N_btm C2_N_btm 5.24136f
C2607 C0_N_btm C3_N_btm 0.409238f
C2608 a_18287_44626# VDD 0.389383f
C2609 a_4361_42308# a_21195_42852# 0.020952f
C2610 a_13467_32519# a_21671_42860# 0.015185f
C2611 a_743_42282# a_n2293_42282# 0.058933f
C2612 a_21101_45002# a_20766_44850# 0.01337f
C2613 a_11827_44484# a_20679_44626# 0.030022f
C2614 a_18184_42460# a_18579_44172# 0.161593f
C2615 a_20193_45348# a_11967_42832# 0.01602f
C2616 a_18114_32519# a_17517_44484# 0.055077f
C2617 a_n755_45592# a_743_42282# 0.160592f
C2618 a_10227_46804# a_13556_45296# 0.013693f
C2619 a_11453_44696# a_3232_43370# 0.132496f
C2620 a_18985_46122# a_19900_46494# 0.118759f
C2621 a_9290_44172# a_526_44458# 0.200352f
C2622 a_8016_46348# a_5066_45546# 0.054471f
C2623 a_17538_32519# EN_VIN_BSTR_N 0.068222f
C2624 a_2711_45572# a_19339_43156# 0.020184f
C2625 a_11309_47204# DATA[5] 0.080873f
C2626 a_1115_44172# a_453_43940# 0.150214f
C2627 a_1467_44172# a_1414_42308# 0.335735f
C2628 a_20202_43084# a_13258_32519# 0.685083f
C2629 a_13059_46348# a_1307_43914# 0.04241f
C2630 a_3483_46348# a_3357_43084# 0.030022f
C2631 a_2107_46812# a_8975_43940# 0.075583f
C2632 a_n755_45592# a_2277_45546# 0.065177f
C2633 a_10809_44734# a_8696_44636# 0.117876f
C2634 a_1138_42852# a_n2661_45010# 0.017849f
C2635 a_n1613_43370# a_n2661_42834# 0.112184f
C2636 a_3090_45724# a_n2293_42834# 0.023056f
C2637 a_16327_47482# a_19279_43940# 0.446333f
C2638 a_9127_43156# VDD 0.468721f
C2639 a_n2109_47186# a_n1435_47204# 0.041807f
C2640 a_n1741_47186# a_11459_47204# 0.015445f
C2641 a_n237_47217# a_7227_47204# 0.013654f
C2642 a_2063_45854# a_4791_45118# 0.039758f
C2643 a_n1151_42308# a_3381_47502# 0.051194f
C2644 a_n971_45724# a_6575_47204# 0.01923f
C2645 a_584_46384# a_n443_46116# 0.496286f
C2646 a_1755_42282# a_6123_31319# 0.033073f
C2647 a_5267_42460# a_4921_42308# 0.04229f
C2648 a_14539_43914# a_17333_42852# 0.072085f
C2649 a_2804_46116# VDD 0.159351f
C2650 a_10193_42453# a_n913_45002# 0.562004f
C2651 a_n2293_46098# a_n2661_42834# 0.029385f
C2652 a_13661_43548# a_13565_43940# 0.017205f
C2653 a_12549_44172# a_20974_43370# 0.061866f
C2654 a_n1613_43370# a_n1352_43396# 0.244933f
C2655 a_n755_45592# a_626_44172# 0.100613f
C2656 a_n3420_39616# a_n4334_39392# 0.014828f
C2657 a_3626_43646# a_4361_42308# 5.20633f
C2658 a_12293_43646# a_12281_43396# 0.01129f
C2659 a_10193_42453# CLK 0.023289f
C2660 a_13904_45546# VDD 0.135068f
C2661 a_n967_45348# a_n2661_43370# 0.016831f
C2662 a_n2293_46634# a_3483_46348# 0.157275f
C2663 a_n971_45724# a_n2661_45546# 0.083094f
C2664 a_12891_46348# a_13351_46090# 0.019821f
C2665 a_12549_44172# a_12594_46348# 0.031894f
C2666 a_n743_46660# a_167_45260# 0.045398f
C2667 a_383_46660# a_805_46414# 0.01072f
C2668 a_n2312_39304# a_n2956_38680# 0.048558f
C2669 a_n2661_46098# a_n2840_46090# 0.170439f
C2670 VDAC_P EN_VIN_BSTR_P 0.340512f
C2671 VDAC_N a_10890_34112# 0.067549f
C2672 a_n97_42460# a_14635_42282# 0.077798f
C2673 a_12089_42308# a_12545_42858# 0.261463f
C2674 a_12379_42858# a_13113_42826# 0.06628f
C2675 a_17023_45118# VDD 0.086861f
C2676 a_4223_44672# a_4743_44484# 0.043867f
C2677 a_4185_45028# a_5534_30871# 0.05188f
C2678 a_n2661_44458# a_8975_43940# 0.075732f
C2679 a_584_46384# a_3537_45260# 0.108506f
C2680 a_18597_46090# a_20107_45572# 0.069963f
C2681 a_n881_46662# a_8696_44636# 0.178516f
C2682 a_18479_47436# a_20841_45814# 0.011134f
C2683 a_12741_44636# a_20075_46420# 0.027561f
C2684 a_3090_45724# a_16375_45002# 0.026416f
C2685 a_22365_46825# a_22223_46124# 0.011912f
C2686 a_3483_46348# a_9625_46129# 0.038063f
C2687 a_20202_43084# a_6945_45028# 0.02248f
C2688 a_11453_44696# a_18341_45572# 0.026938f
C2689 a_1847_42826# a_2351_42308# 0.120686f
C2690 a_5342_30871# a_14097_32519# 0.028503f
C2691 a_n356_44636# a_n2661_42282# 2.54767f
C2692 a_13717_47436# VDD 0.314317f
C2693 a_6575_47204# DATA[3] 0.055018f
C2694 a_n2661_42834# a_2675_43914# 0.024352f
C2695 a_n1435_47204# RST_Z 0.179508f
C2696 a_n1059_45260# a_16243_43396# 0.012252f
C2697 a_526_44458# a_8292_43218# 0.02177f
C2698 a_17517_44484# a_22485_44484# 0.110643f
C2699 a_20835_44721# a_19279_43940# 0.036128f
C2700 a_13661_43548# a_11691_44458# 0.263889f
C2701 a_n1613_43370# a_n1352_44484# 0.232498f
C2702 a_2324_44458# a_7499_43078# 0.018394f
C2703 a_8270_45546# a_6171_45002# 0.027058f
C2704 a_3090_45724# a_413_45260# 0.135828f
C2705 a_4791_45118# a_n2661_42834# 0.024946f
C2706 a_11453_44696# a_8975_43940# 0.027482f
C2707 a_12465_44636# a_13720_44458# 0.019702f
C2708 a_10903_43370# a_11962_45724# 0.357882f
C2709 a_19268_43646# VDD 0.237793f
C2710 a_n2472_42282# a_n4318_38216# 0.157105f
C2711 a_n2840_42282# a_n3674_38216# 0.03703f
C2712 a_2479_44172# a_n97_42460# 0.196935f
C2713 a_n2956_38680# a_n3420_38528# 0.233147f
C2714 a_14035_46660# VDD 0.363878f
C2715 a_n2472_45546# a_n2472_45002# 0.026152f
C2716 a_584_46384# a_1049_43396# 0.148494f
C2717 a_n357_42282# a_3357_43084# 0.010127f
C2718 a_18479_47436# a_13661_43548# 0.024025f
C2719 a_2905_45572# a_3524_46660# 0.011982f
C2720 a_n237_47217# a_4955_46873# 0.032268f
C2721 a_12465_44636# a_12549_44172# 0.093222f
C2722 a_11599_46634# a_n2661_46634# 0.067552f
C2723 a_22165_42308# VDD 0.336187f
C2724 a_6031_43396# a_6452_43396# 0.086708f
C2725 en_comp a_7174_31319# 5.65156f
C2726 a_19319_43548# a_15743_43084# 0.035611f
C2727 a_n1099_45572# VDD 0.89411f
C2728 a_20205_31679# VIN_N 0.028376f
C2729 a_3483_46348# a_9672_43914# 0.125466f
C2730 a_10227_46804# a_10991_42826# 0.152133f
C2731 a_13661_43548# a_4190_30871# 0.147163f
C2732 a_n1613_43370# a_n1423_42826# 0.15981f
C2733 a_2063_45854# a_6945_45028# 0.074119f
C2734 VDAC_Pi a_5088_37509# 0.391059f
C2735 a_7754_40130# VDAC_N 0.434929f
C2736 a_n4064_39072# C7_P_btm 0.072179f
C2737 a_7754_39964# a_5700_37509# 0.095724f
C2738 a_n1423_42826# a_n1533_42852# 0.097745f
C2739 a_10951_45334# VDD 0.226705f
C2740 a_11823_42460# a_12429_44172# 0.018664f
C2741 a_21005_45260# a_21101_45002# 0.419086f
C2742 a_18494_42460# a_11827_44484# 0.031498f
C2743 a_3065_45002# a_n2661_43922# 0.023551f
C2744 a_10193_42453# a_18451_43940# 0.20167f
C2745 a_4185_45028# a_4190_30871# 0.16524f
C2746 a_18911_45144# a_19113_45348# 0.054737f
C2747 a_5147_45002# a_5708_44484# 0.055267f
C2748 a_13661_43548# a_n443_42852# 0.045364f
C2749 a_11453_44696# a_10193_42453# 0.071253f
C2750 a_12549_44172# a_2711_45572# 2.05236f
C2751 a_15227_44166# a_2324_44458# 0.190521f
C2752 a_n2293_46634# a_n357_42282# 0.034749f
C2753 a_18249_42858# a_19164_43230# 0.118759f
C2754 a_n357_42282# a_5342_30871# 0.039779f
C2755 a_n913_45002# a_3080_42308# 0.044741f
C2756 a_n1059_45260# a_4905_42826# 0.027099f
C2757 a_742_44458# a_2479_44172# 0.019563f
C2758 a_n699_43396# a_1467_44172# 0.030347f
C2759 a_n2956_39768# a_n2946_39866# 0.14868f
C2760 a_n2442_46660# a_n3565_39590# 0.134948f
C2761 a_4185_45028# a_n443_42852# 0.027973f
C2762 a_19335_46494# a_19240_46482# 0.049827f
C2763 a_n1151_42308# a_n699_43396# 0.022019f
C2764 a_n357_42282# a_n473_42460# 0.179066f
C2765 a_n2956_38680# a_n2810_45028# 0.043221f
C2766 a_8049_45260# a_20107_45572# 0.024509f
C2767 a_n2956_39304# a_n2956_37592# 0.044994f
C2768 a_n1613_43370# a_n1549_44318# 0.16289f
C2769 a_2711_45572# a_11525_45546# 0.0154f
C2770 a_15673_47210# a_16588_47582# 0.125324f
C2771 a_584_46384# a_n1613_43370# 0.085833f
C2772 a_15507_47210# a_10227_46804# 0.23187f
C2773 a_16327_47482# a_16023_47582# 0.159305f
C2774 a_n97_42460# a_n229_43646# 0.046961f
C2775 a_11967_42832# a_5534_30871# 0.017079f
C2776 a_15682_43940# a_16759_43396# 0.013707f
C2777 a_n1925_42282# VDD 0.728256f
C2778 a_3065_45002# a_3318_42354# 0.146272f
C2779 en_comp a_5932_42308# 0.23313f
C2780 a_n913_45002# a_7227_42308# 0.052824f
C2781 a_n2661_46634# a_7411_46660# 0.023716f
C2782 a_584_46384# a_n2293_46098# 0.039917f
C2783 a_11599_46634# a_765_45546# 0.332797f
C2784 a_2107_46812# a_4646_46812# 0.03082f
C2785 a_3177_46902# a_2959_46660# 0.209641f
C2786 a_2609_46660# a_3699_46634# 0.042415f
C2787 a_2443_46660# a_3524_46660# 0.102325f
C2788 a_5807_45002# a_10249_46116# 0.041839f
C2789 a_n3565_39590# a_n3420_37440# 0.035128f
C2790 a_n4209_39590# a_n4064_37440# 0.033425f
C2791 a_5742_30871# C4_N_btm 0.03103f
C2792 a_n2302_38778# a_n2302_37984# 0.052227f
C2793 a_n4064_39616# a_n4209_37414# 0.028043f
C2794 a_n3420_39616# a_n3565_37414# 0.028169f
C2795 a_9803_42558# VDD 0.253745f
C2796 a_15743_43084# a_19095_43396# 0.012939f
C2797 a_9290_44172# a_3626_43646# 0.014922f
C2798 a_6151_47436# a_6472_45840# 0.045851f
C2799 a_2063_45854# a_6812_45938# 0.026385f
C2800 a_18597_46090# a_n357_42282# 0.250702f
C2801 a_5257_43370# a_5937_45572# 0.262028f
C2802 a_6755_46942# a_3483_46348# 0.014154f
C2803 a_n1696_34930# VIN_P 0.068773f
C2804 C7_P_btm VDD 0.121904f
C2805 C0_dummy_N_btm C3_N_btm 0.087354f
C2806 C0_N_btm C2_N_btm 0.827449f
C2807 a_18248_44752# VDD 0.251171f
C2808 a_3080_42308# a_1755_42282# 0.047244f
C2809 a_4361_42308# a_21356_42826# 0.017293f
C2810 a_13467_32519# a_21195_42852# 0.034759f
C2811 a_6298_44484# a_n2661_43922# 0.048814f
C2812 a_n2293_42834# a_1414_42308# 0.02233f
C2813 a_10193_42453# a_9145_43396# 0.02642f
C2814 a_19778_44110# a_18579_44172# 0.268475f
C2815 a_11827_44484# a_20640_44752# 0.016882f
C2816 a_11691_44458# a_11967_42832# 0.041904f
C2817 a_5883_43914# a_9159_44484# 0.049132f
C2818 a_n357_42282# a_743_42282# 0.067793f
C2819 a_7920_46348# a_5066_45546# 0.04093f
C2820 a_3483_46348# a_8049_45260# 0.012066f
C2821 a_768_44030# a_n2661_45010# 0.015059f
C2822 a_10227_46804# a_9482_43914# 0.032461f
C2823 a_8270_45546# a_8746_45002# 0.017581f
C2824 a_18985_46122# a_20075_46420# 0.042415f
C2825 a_18819_46122# a_19900_46494# 0.102355f
C2826 a_19553_46090# a_19335_46494# 0.209641f
C2827 a_13747_46662# a_21513_45002# 0.02166f
C2828 a_3737_43940# VDD 0.18423f
C2829 a_12089_42308# a_12563_42308# 0.03299f
C2830 a_n1925_42282# a_n784_42308# 0.235613f
C2831 a_644_44056# a_453_43940# 0.077973f
C2832 a_n913_45002# a_2075_43172# 0.175893f
C2833 a_1115_44172# a_1414_42308# 0.134389f
C2834 a_8953_45546# a_9885_42558# 0.024699f
C2835 a_n2661_45546# a_2711_45572# 0.359276f
C2836 a_18479_47436# a_11967_42832# 0.017885f
C2837 SMPL_ON_P a_n3674_39768# 0.03705f
C2838 a_4646_46812# a_n2661_44458# 0.05901f
C2839 a_997_45618# a_n443_42852# 0.093108f
C2840 a_n755_45592# a_1609_45822# 0.12055f
C2841 a_21076_30879# a_413_45260# 0.141502f
C2842 a_n356_45724# a_n23_45546# 0.360492f
C2843 a_16327_47482# a_20766_44850# 0.17113f
C2844 a_8387_43230# VDD 0.200672f
C2845 a_n1741_47186# a_9313_45822# 0.102019f
C2846 a_3160_47472# a_3381_47502# 0.099936f
C2847 a_2905_45572# a_3785_47178# 0.013619f
C2848 a_1606_42308# a_6123_31319# 1.43958f
C2849 a_5891_43370# a_8037_42858# 0.12253f
C2850 a_3422_30871# a_15743_43084# 0.022574f
C2851 a_2698_46116# VDD 0.195879f
C2852 a_19479_31679# a_14097_32519# 0.05096f
C2853 a_n1059_45260# a_15597_42852# 0.056846f
C2854 a_10193_42453# a_n1059_45260# 0.440111f
C2855 a_n1613_43370# a_n1177_43370# 0.325171f
C2856 a_13507_46334# a_2982_43646# 0.063751f
C2857 a_n357_42282# a_626_44172# 0.551369f
C2858 a_n1151_42308# a_14084_46812# 0.063788f
C2859 a_9804_47204# a_2107_46812# 0.033493f
C2860 a_1606_42308# EN_VIN_BSTR_P 0.035204f
C2861 a_n1794_35082# a_21753_35474# 0.018844f
C2862 a_n3565_39590# a_n3565_39304# 0.046203f
C2863 a_n4209_39590# a_n3420_39072# 0.034738f
C2864 a_n3420_39616# a_n4209_39304# 0.05141f
C2865 a_10180_45724# CLK 0.095799f
C2866 a_3422_30871# a_21671_42860# 0.199876f
C2867 a_13527_45546# VDD 0.1902f
C2868 en_comp a_n2661_43370# 0.164814f
C2869 a_14537_43396# a_14797_45144# 0.082443f
C2870 a_9482_43914# a_1307_43914# 0.010221f
C2871 a_8696_44636# a_8701_44490# 0.095858f
C2872 a_12891_46348# a_12594_46348# 0.088156f
C2873 a_n2312_40392# a_n2956_38680# 0.052782f
C2874 a_n2312_39304# a_n2956_39304# 6.38528f
C2875 a_6755_46942# a_14513_46634# 0.036712f
C2876 a_5807_45002# a_5937_45572# 0.038681f
C2877 a_n743_46660# a_2202_46116# 0.012092f
C2878 a_768_44030# a_10903_43370# 0.082359f
C2879 a_22581_37893# a_22629_38406# 0.236891f
C2880 a_7754_39300# VDD 0.048307f
C2881 a_22589_40055# a_22725_37990# 0.016815f
C2882 a_22537_40625# a_22737_36887# 0.011861f
C2883 a_22527_39145# a_22629_37990# 0.172129f
C2884 VDAC_P a_n1057_35014# 0.057328f
C2885 a_12379_42858# a_12545_42858# 0.810394f
C2886 a_n97_42460# a_13291_42460# 0.419357f
C2887 a_18114_32519# EN_VIN_BSTR_N 0.149623f
C2888 a_16922_45042# VDD 1.54713f
C2889 a_4223_44672# a_n699_43396# 0.217586f
C2890 SMPL_ON_P a_n4315_30879# 3.7658f
C2891 a_11691_44458# a_18989_43940# 0.066207f
C2892 a_413_45260# a_1414_42308# 0.12534f
C2893 a_n881_46662# a_16680_45572# 0.051767f
C2894 a_18479_47436# a_20273_45572# 0.028755f
C2895 a_15368_46634# a_13259_45724# 0.0178f
C2896 a_3483_46348# a_8953_45546# 0.133493f
C2897 a_n2293_46634# a_13249_42308# 0.027384f
C2898 a_5257_43370# a_n443_42852# 0.016836f
C2899 a_4361_42308# a_8685_42308# 0.014949f
C2900 a_n2661_42834# a_895_43940# 0.095907f
C2901 a_9482_43914# a_9396_43370# 0.011522f
C2902 a_n1059_45260# a_16137_43396# 0.438785f
C2903 a_17517_44484# a_20512_43084# 0.027951f
C2904 a_20835_44721# a_20766_44850# 0.209641f
C2905 a_20679_44626# a_19279_43940# 0.279785f
C2906 a_n1435_47204# VDD 0.267875f
C2907 a_7903_47542# DATA[3] 0.01066f
C2908 a_5807_45002# a_11691_44458# 0.117249f
C2909 a_n1613_43370# a_n1177_44458# 0.332209f
C2910 a_8270_45546# a_3232_43370# 0.020859f
C2911 a_12465_44636# a_13076_44458# 0.01224f
C2912 a_10903_43370# a_11652_45724# 0.010404f
C2913 a_19321_45002# a_11827_44484# 0.037739f
C2914 a_13887_32519# EN_VIN_BSTR_N 0.031797f
C2915 a_15743_43084# VDD 0.572249f
C2916 a_n3674_38680# a_n4318_38216# 2.82961f
C2917 a_15493_43940# a_22959_43948# 0.182001f
C2918 a_n2956_38680# a_n3690_38528# 0.015398f
C2919 a_13885_46660# VDD 0.499249f
C2920 a_n971_45724# a_n1557_42282# 0.06901f
C2921 a_12549_44172# a_15682_43940# 0.058263f
C2922 a_n1925_42282# a_1423_45028# 0.021671f
C2923 a_584_46384# a_1209_43370# 0.02923f
C2924 a_2324_44458# a_n2661_43370# 0.082794f
C2925 a_n2956_38216# a_n2840_45002# 0.01122f
C2926 a_4883_46098# a_768_44030# 0.045313f
C2927 a_10227_46804# a_13747_46662# 0.16398f
C2928 a_18143_47464# a_13661_43548# 0.011802f
C2929 a_9313_45822# a_n743_46660# 0.029372f
C2930 a_12465_44636# a_12891_46348# 0.033919f
C2931 a_6545_47178# a_2107_46812# 0.028617f
C2932 a_17303_42282# a_13258_32519# 0.064259f
C2933 a_21671_42860# VDD 0.229963f
C2934 a_380_45546# VDD 0.154763f
C2935 a_6765_43638# a_7112_43396# 0.051162f
C2936 a_n913_45002# a_21613_42308# 0.259761f
C2937 a_10227_46804# a_10796_42968# 0.024053f
C2938 a_n1613_43370# a_n1991_42858# 0.029351f
C2939 a_8667_46634# a_8492_46660# 0.233657f
C2940 a_4915_47217# a_2324_44458# 0.022906f
C2941 a_13747_46662# a_17339_46660# 0.015626f
C2942 VDAC_Pi a_4338_37500# 1.92369f
C2943 a_n3420_39072# C6_P_btm 0.054459f
C2944 a_7754_39964# a_5088_37509# 0.392826f
C2945 a_n1991_42858# a_n1533_42852# 0.034619f
C2946 a_n3674_39304# a_n4318_38680# 2.92578f
C2947 a_5649_42852# a_5755_42852# 0.089078f
C2948 a_n2661_42282# a_n2840_42282# 0.173771f
C2949 a_10775_45002# VDD 0.148349f
C2950 a_18184_42460# a_11827_44484# 0.027981f
C2951 a_3065_45002# a_n2661_42834# 0.022516f
C2952 a_10193_42453# a_18326_43940# 0.130866f
C2953 a_n2293_46634# a_310_45028# 0.020873f
C2954 a_n881_46662# a_6598_45938# 0.031336f
C2955 a_4791_45118# a_8696_44636# 0.097007f
C2956 a_n2438_43548# a_n2293_45546# 0.051617f
C2957 a_12891_46348# a_2711_45572# 0.027614f
C2958 a_12741_44636# a_22959_46660# 0.17409f
C2959 a_20820_30879# a_21076_30879# 8.6867f
C2960 a_11735_46660# a_10809_44734# 0.030929f
C2961 a_18817_42826# a_18599_43230# 0.209641f
C2962 a_18249_42858# a_19339_43156# 0.042415f
C2963 a_8037_42858# a_8292_43218# 0.064178f
C2964 a_5111_42852# a_5193_42852# 0.171361f
C2965 a_n1059_45260# a_3080_42308# 0.025424f
C2966 a_n2017_45002# a_4905_42826# 0.042734f
C2967 a_13249_42308# a_743_42282# 0.010211f
C2968 a_2382_45260# a_n97_42460# 0.02063f
C2969 a_11823_42460# a_4361_42308# 0.056415f
C2970 a_n2956_39768# a_n3420_39616# 0.233256f
C2971 a_n2661_46634# a_13159_45002# 0.062031f
C2972 a_17957_46116# a_18051_46116# 0.062574f
C2973 a_8953_45546# a_n357_42282# 0.054106f
C2974 a_2959_46660# a_413_45260# 0.011261f
C2975 a_3539_42460# VDD 0.363092f
C2976 a_10057_43914# a_9145_43396# 0.121499f
C2977 a_13059_46348# a_11827_44484# 0.495367f
C2978 a_8270_45546# a_8975_43940# 0.207334f
C2979 a_n2956_39304# a_n2810_45028# 0.042912f
C2980 a_7227_45028# a_7230_45938# 0.170618f
C2981 a_n1613_43370# a_n1331_43914# 0.16678f
C2982 a_8016_46348# a_9482_43914# 0.293982f
C2983 a_2711_45572# a_11322_45546# 0.056109f
C2984 a_15673_47210# a_16763_47508# 0.042509f
C2985 a_16241_47178# a_16023_47582# 0.209641f
C2986 a_11599_46634# a_10227_46804# 0.60865f
C2987 a_12861_44030# a_18597_46090# 0.045766f
C2988 a_n3674_37592# a_n4064_40160# 0.022617f
C2989 a_n4318_37592# a_n3420_39616# 0.020563f
C2990 a_n1794_35082# a_n4315_30879# 0.133824f
C2991 a_n3674_38216# a_n4064_39616# 0.020042f
C2992 a_n447_43370# a_n229_43646# 0.08213f
C2993 a_11967_42832# a_14543_43071# 0.022161f
C2994 a_14021_43940# a_9145_43396# 0.032057f
C2995 a_526_44458# VDD 2.35177f
C2996 a_2382_45260# a_3823_42558# 0.058499f
C2997 a_n913_45002# a_6761_42308# 0.350952f
C2998 a_10809_44734# a_10617_44484# 0.014699f
C2999 a_3090_45724# a_11341_43940# 0.041393f
C3000 a_11453_44696# a_19692_46634# 0.05834f
C3001 a_11599_46634# a_17339_46660# 0.131185f
C3002 a_2107_46812# a_3877_44458# 0.070722f
C3003 a_n746_45260# a_376_46348# 0.010981f
C3004 a_2443_46660# a_3699_46634# 0.043475f
C3005 a_2609_46660# a_2959_46660# 0.216095f
C3006 a_9223_42460# VDD 0.205797f
C3007 a_5742_30871# C3_N_btm 0.030866f
C3008 a_18783_43370# a_19095_43396# 0.038241f
C3009 a_5891_43370# a_8685_42308# 0.048111f
C3010 a_413_45260# a_n699_43396# 0.100762f
C3011 a_13556_45296# a_11827_44484# 0.05613f
C3012 a_14976_45028# a_11415_45002# 0.039578f
C3013 a_4791_45118# a_7227_45028# 0.288276f
C3014 a_6151_47436# a_6194_45824# 0.227219f
C3015 a_n1550_35448# VIN_P 0.37444f
C3016 C8_P_btm VDD 0.19922f
C3017 C0_dummy_N_btm C2_N_btm 7.14548f
C3018 C0_N_btm C1_N_btm 11.2332f
C3019 a_17970_44736# VDD 0.27753f
C3020 a_3080_42308# a_1606_42308# 4.87174f
C3021 a_10440_44484# CLK 0.013272f
C3022 a_20692_30879# a_17364_32525# 0.054134f
C3023 a_5518_44484# a_n2661_43922# 0.011667f
C3024 a_n356_44636# a_n23_44458# 0.220577f
C3025 a_18494_42460# a_19279_43940# 0.137363f
C3026 a_21359_45002# a_20640_44752# 0.013689f
C3027 a_6419_46155# a_5066_45546# 0.038923f
C3028 a_n1151_42308# a_n2293_42834# 0.051075f
C3029 a_765_45546# a_997_45618# 0.026457f
C3030 a_18819_46122# a_20075_46420# 0.043567f
C3031 a_18985_46122# a_19335_46494# 0.210876f
C3032 a_2324_44458# a_10809_44734# 0.026995f
C3033 a_n1613_43370# a_n967_45348# 0.213625f
C3034 a_14401_32519# EN_VIN_BSTR_N 0.814839f
C3035 a_175_44278# a_453_43940# 0.112594f
C3036 a_n913_45002# a_1847_42826# 0.294312f
C3037 a_1115_44172# a_1467_44172# 0.115277f
C3038 a_526_44458# a_n784_42308# 0.011818f
C3039 a_13259_45724# a_13291_42460# 0.089962f
C3040 a_20202_43084# a_19511_42282# 0.082529f
C3041 SMPL_ON_P a_n4318_39768# 0.039185f
C3042 a_22959_46660# a_413_45260# 0.018266f
C3043 a_584_46384# a_895_43940# 0.025246f
C3044 a_3877_44458# a_n2661_44458# 0.035165f
C3045 a_n755_45592# a_n443_42852# 0.469263f
C3046 a_16327_47482# a_20835_44721# 0.157393f
C3047 a_8605_42826# VDD 0.204898f
C3048 a_5342_30871# C6_P_btm 0.012f
C3049 a_n2497_47436# a_n1435_47204# 0.010029f
C3050 a_2905_45572# a_3381_47502# 0.208262f
C3051 a_3160_47472# a_n1151_42308# 0.357683f
C3052 a_14539_43914# a_17701_42308# 0.039977f
C3053 a_5891_43370# a_7765_42852# 0.168516f
C3054 a_n2661_42282# a_6197_43396# 0.033187f
C3055 a_2521_46116# VDD 0.163553f
C3056 a_10193_42453# a_n2017_45002# 0.081859f
C3057 a_12549_44172# a_21381_43940# 0.099617f
C3058 a_n1613_43370# a_n1917_43396# 0.153085f
C3059 a_n863_45724# a_2304_45348# 0.091195f
C3060 a_n755_45592# a_375_42282# 0.366231f
C3061 a_11599_46634# a_10467_46802# 0.261176f
C3062 a_5807_45002# a_n2661_46634# 0.087532f
C3063 a_2747_46873# a_2864_46660# 0.174836f
C3064 a_8128_46384# a_2107_46812# 0.028382f
C3065 a_12861_44030# a_6755_46942# 0.376009f
C3066 a_4958_30871# a_n4064_37984# 0.030919f
C3067 a_n1794_35082# a_19998_34978# 0.020261f
C3068 a_3422_30871# a_21195_42852# 0.289298f
C3069 a_2982_43646# a_4361_42308# 0.545077f
C3070 a_13163_45724# VDD 0.322298f
C3071 a_14358_43442# a_14621_43646# 0.011552f
C3072 a_n2956_37592# a_n2661_43370# 0.044152f
C3073 a_20692_30879# a_19237_31679# 0.051625f
C3074 a_14180_45002# a_14797_45144# 0.070624f
C3075 a_3090_45724# a_10341_43396# 0.07129f
C3076 a_5691_45260# a_5837_45348# 0.013377f
C3077 a_2711_45572# a_16241_44734# 0.03035f
C3078 a_12861_44030# a_8049_45260# 0.109405f
C3079 a_n2438_43548# a_1138_42852# 0.646257f
C3080 a_n881_46662# a_2324_44458# 0.085939f
C3081 a_n2312_40392# a_n2956_39304# 0.052343f
C3082 SMPL_ON_P a_n2956_38216# 0.0385f
C3083 a_12549_44172# a_10903_43370# 0.792848f
C3084 a_n743_46660# a_1823_45246# 0.04372f
C3085 a_6755_46942# a_14180_46812# 0.063843f
C3086 a_13607_46688# a_14084_46812# 0.014875f
C3087 a_22581_37893# CAL_P 0.026818f
C3088 a_n4209_37414# C1_P_btm 0.043983f
C3089 a_22589_40055# a_22629_37990# 0.234448f
C3090 a_n4064_37984# VCM 0.011087f
C3091 a_12379_42858# a_12089_42308# 0.16885f
C3092 a_8953_45546# a_8952_43230# 0.01883f
C3093 a_11691_44458# a_18374_44850# 0.02267f
C3094 a_2779_44458# a_n699_43396# 0.025176f
C3095 a_n971_45724# a_6171_45002# 0.030962f
C3096 a_n1151_42308# a_413_45260# 0.135643f
C3097 a_n881_46662# a_16855_45546# 0.052296f
C3098 a_584_46384# a_3065_45002# 0.085314f
C3099 a_13717_47436# a_3357_43084# 0.024679f
C3100 a_18479_47436# a_20107_45572# 0.025968f
C3101 a_16327_47482# a_20731_45938# 0.012637f
C3102 a_5204_45822# a_5497_46414# 0.099282f
C3103 a_765_45546# a_1337_46116# 0.011452f
C3104 a_3483_46348# a_5937_45572# 0.767636f
C3105 a_14976_45028# a_13259_45724# 0.018965f
C3106 a_11453_44696# a_18175_45572# 0.036949f
C3107 a_5534_30871# a_14097_32519# 0.041746f
C3108 a_4361_42308# a_8325_42308# 0.020707f
C3109 a_19615_44636# a_18579_44172# 0.158449f
C3110 a_5111_44636# a_9803_43646# 0.118936f
C3111 a_n2661_42834# a_2479_44172# 0.027713f
C3112 a_n2017_45002# a_16137_43396# 0.63011f
C3113 a_20640_44752# a_19279_43940# 0.22152f
C3114 a_20679_44626# a_20766_44850# 0.052825f
C3115 a_13381_47204# VDD 0.130765f
C3116 a_7227_47204# DATA[3] 0.357377f
C3117 a_6151_47436# CLK 0.036587f
C3118 a_10903_43370# a_11525_45546# 0.040993f
C3119 a_n1613_43370# a_n1917_44484# 0.153277f
C3120 a_6945_45028# a_7227_45028# 0.016808f
C3121 a_9290_44172# a_11823_42460# 0.864145f
C3122 a_12465_44636# a_12883_44458# 0.017889f
C3123 a_n2840_42282# a_n4318_38216# 0.015074f
C3124 a_18783_43370# VDD 0.289099f
C3125 a_n2956_38680# a_n3565_38502# 0.302523f
C3126 a_9313_44734# a_16547_43609# 0.010576f
C3127 a_12549_44172# a_14955_43940# 0.010132f
C3128 a_n755_45592# a_2437_43646# 0.017992f
C3129 a_3483_46348# a_11691_44458# 0.039125f
C3130 a_4185_45028# a_22959_45036# 0.17601f
C3131 a_3090_45724# a_n2293_43922# 0.02667f
C3132 a_n2661_45546# a_n2661_45010# 0.014492f
C3133 a_526_44458# a_1423_45028# 0.133656f
C3134 a_584_46384# a_458_43396# 0.196763f
C3135 a_4883_46098# a_12549_44172# 0.021771f
C3136 a_n237_47217# a_4646_46812# 0.020773f
C3137 a_10227_46804# a_13661_43548# 0.072131f
C3138 a_6151_47436# a_2107_46812# 0.019997f
C3139 a_4958_30871# a_13258_32519# 0.033151f
C3140 a_21195_42852# VDD 0.285496f
C3141 a_14021_43940# a_22959_43396# 0.191956f
C3142 a_6197_43396# a_7112_43396# 0.118423f
C3143 a_20193_45348# a_22400_42852# 0.05078f
C3144 a_n452_45724# VDD 0.112977f
C3145 a_n913_45002# a_21887_42336# 0.060677f
C3146 a_n1613_43370# a_n1853_43023# 0.423772f
C3147 a_413_45260# a_327_44734# 0.195096f
C3148 a_10227_46804# a_10835_43094# 0.295543f
C3149 a_13661_43548# a_19177_43646# 0.015951f
C3150 a_n913_45002# a_5111_44636# 0.070773f
C3151 a_n2497_47436# a_526_44458# 0.06857f
C3152 a_n443_46116# a_2324_44458# 0.055032f
C3153 a_5807_45002# a_765_45546# 0.103324f
C3154 a_13661_43548# a_17339_46660# 0.599051f
C3155 a_n2302_40160# VDD 0.428934f
C3156 a_7754_38636# a_7754_38470# 0.296258f
C3157 VDAC_Pi a_3726_37500# 1.17174f
C3158 a_7174_31319# VIN_N 0.022822f
C3159 a_13258_32519# VCM 0.033198f
C3160 a_7754_39964# a_4338_37500# 0.021449f
C3161 a_7754_40130# a_5700_37509# 0.037095f
C3162 a_15743_43084# a_15567_42826# 0.215954f
C3163 a_8953_45002# VDD 1.24336f
C3164 a_5649_42852# a_5111_42852# 0.110096f
C3165 a_1823_45246# a_4361_42308# 0.11884f
C3166 a_20567_45036# a_21005_45260# 0.015494f
C3167 a_19778_44110# a_11827_44484# 0.029054f
C3168 a_n2293_42834# a_4223_44672# 0.015649f
C3169 a_2382_45260# a_n2661_43922# 0.026472f
C3170 a_10193_42453# a_18079_43940# 0.076581f
C3171 a_n2438_43548# a_n2956_38216# 0.020852f
C3172 a_20820_30879# a_22959_46660# 0.01739f
C3173 a_18249_42858# a_18599_43230# 0.210876f
C3174 a_18083_42858# a_19164_43230# 0.101963f
C3175 a_4190_30871# a_14097_32519# 0.031855f
C3176 a_7765_42852# a_8292_43218# 0.157652f
C3177 a_n2017_45002# a_3080_42308# 0.034898f
C3178 a_n357_42282# a_5534_30871# 0.04831f
C3179 a_1307_43914# a_5829_43940# 0.016223f
C3180 a_n2956_39768# a_n3690_39616# 0.015398f
C3181 a_n2442_46660# a_n4209_39590# 0.095025f
C3182 a_n2661_46634# a_13017_45260# 0.123713f
C3183 a_18985_46122# a_19240_46482# 0.05936f
C3184 a_18189_46348# a_18051_46116# 0.045453f
C3185 a_12861_44030# a_20193_45348# 0.680394f
C3186 a_13661_43548# a_1307_43914# 0.396211f
C3187 a_3626_43646# VDD 0.340378f
C3188 a_n2293_42282# COMP_P 0.026882f
C3189 a_5275_47026# VDD 0.135766f
C3190 a_19321_45002# a_19279_43940# 0.019898f
C3191 a_13661_43548# a_18579_44172# 0.229269f
C3192 a_2711_45572# a_10490_45724# 0.036939f
C3193 a_2324_44458# a_3537_45260# 0.015845f
C3194 a_n1925_42282# a_3357_43084# 0.067793f
C3195 a_4185_45028# a_1307_43914# 0.025209f
C3196 a_n1613_43370# a_n1899_43946# 0.038349f
C3197 a_15673_47210# a_16023_47582# 0.228897f
C3198 a_15507_47210# a_16588_47582# 0.102325f
C3199 a_14955_47212# a_10227_46804# 0.175517f
C3200 a_16241_47178# a_16327_47482# 0.185907f
C3201 a_15493_43396# a_15781_43660# 0.047833f
C3202 a_11967_42832# a_13460_43230# 0.038517f
C3203 a_20193_45348# a_22223_42860# 0.017179f
C3204 a_2981_46116# VDD 0.111597f
C3205 a_2382_45260# a_3318_42354# 0.028613f
C3206 a_20623_45572# a_20719_45572# 0.013793f
C3207 a_15227_44166# a_15493_43396# 0.046514f
C3208 a_12861_44030# a_18285_46348# 0.247326f
C3209 a_2609_46660# a_3177_46902# 0.17072f
C3210 a_2443_46660# a_2959_46660# 0.110816f
C3211 a_8791_42308# VDD 0.226318f
C3212 a_n3565_39590# a_n3565_37414# 0.032079f
C3213 a_7174_31319# CAL_N 0.018266f
C3214 a_n4209_39590# a_n3420_37440# 0.038354f
C3215 a_5932_42308# VIN_N 0.023512f
C3216 a_5742_30871# C2_N_btm 0.030783f
C3217 a_n3420_39616# a_n4209_37414# 0.027966f
C3218 a_n4064_38528# a_n4064_37984# 0.057015f
C3219 a_5891_43370# a_8325_42308# 0.053347f
C3220 a_5111_44636# a_n2661_44458# 0.048314f
C3221 a_9482_43914# a_11827_44484# 0.031913f
C3222 a_n2956_38680# a_n4318_39304# 0.023179f
C3223 a_3090_45724# a_11415_45002# 0.16525f
C3224 a_6151_47436# a_5907_45546# 0.274247f
C3225 a_7715_46873# a_7920_46348# 0.080253f
C3226 SMPL_ON_N a_20692_30879# 0.029397f
C3227 a_n2293_46634# a_n1925_42282# 0.030317f
C3228 a_n2002_35448# VIN_P 0.029412f
C3229 C9_P_btm VDD 0.345685f
C3230 C0_dummy_N_btm C1_N_btm 1.24905f
C3231 a_17767_44458# VDD 0.348803f
C3232 a_10334_44484# CLK 0.012484f
C3233 a_21487_43396# a_21195_42852# 0.01192f
C3234 a_20205_31679# a_17364_32525# 0.053947f
C3235 a_5343_44458# a_n2661_43922# 0.094786f
C3236 a_n357_42282# a_4190_30871# 0.035963f
C3237 a_413_45260# a_15493_43940# 0.013529f
C3238 a_7499_43078# a_10695_43548# 0.124597f
C3239 a_18184_42460# a_19279_43940# 0.132218f
C3240 a_11827_44484# a_20159_44458# 0.012941f
C3241 a_6165_46155# a_5066_45546# 0.041118f
C3242 a_12741_44636# a_16375_45002# 0.042457f
C3243 a_18819_46122# a_19335_46494# 0.108964f
C3244 a_18985_46122# a_19553_46090# 0.16939f
C3245 a_12465_44636# a_6171_45002# 0.03098f
C3246 a_12089_42308# a_11551_42558# 0.109508f
C3247 a_13678_32519# a_22485_38105# 0.034444f
C3248 a_n699_43396# a_104_43370# 0.21575f
C3249 a_n913_45002# a_791_42968# 0.054288f
C3250 a_n1059_45260# a_1847_42826# 0.038913f
C3251 a_584_46384# a_2479_44172# 0.054912f
C3252 a_10227_46804# a_11967_42832# 0.461417f
C3253 a_n357_42282# a_n443_42852# 0.763015f
C3254 a_10586_45546# a_11962_45724# 0.137051f
C3255 a_16327_47482# a_20679_44626# 0.318301f
C3256 a_12465_44636# a_14673_44172# 0.101564f
C3257 a_n237_47217# a_6545_47178# 0.021104f
C3258 a_2905_45572# a_n1151_42308# 0.072935f
C3259 a_n971_45724# a_6851_47204# 0.028789f
C3260 a_8037_42858# VDD 0.344922f
C3261 a_3823_42558# a_3905_42558# 0.171361f
C3262 a_14539_43914# a_17595_43084# 0.141972f
C3263 a_167_45260# VDD 1.41955f
C3264 a_5891_43370# a_7871_42858# 0.051552f
C3265 a_n2661_42282# a_6293_42852# 0.16527f
C3266 a_17339_46660# a_11967_42832# 0.493072f
C3267 a_5907_45546# a_5111_44636# 0.01337f
C3268 a_n1613_43370# a_n1699_43638# 0.160308f
C3269 a_11415_45002# a_14815_43914# 0.070306f
C3270 a_2711_45572# a_6171_45002# 0.457554f
C3271 a_n357_42282# a_375_42282# 0.142311f
C3272 a_16115_45572# a_16211_45572# 0.013793f
C3273 a_n3565_39590# a_n4209_39304# 5.4667f
C3274 a_n4064_40160# a_n4064_39072# 0.0667f
C3275 a_n4334_39616# a_n4334_39392# 0.052468f
C3276 a_18707_42852# VDD 0.132317f
C3277 a_n4209_39590# a_n3565_39304# 0.032081f
C3278 a_10341_43396# a_12281_43396# 0.012652f
C3279 a_14358_43442# a_14537_43646# 0.010303f
C3280 a_12791_45546# VDD 0.205486f
C3281 a_3422_30871# a_21356_42826# 0.024863f
C3282 a_21363_45546# a_21359_45002# 0.01738f
C3283 a_20205_31679# a_19237_31679# 0.051574f
C3284 a_14180_45002# a_14537_43396# 0.143922f
C3285 a_2711_45572# a_14673_44172# 0.04263f
C3286 a_8953_45002# a_1423_45028# 0.011739f
C3287 a_6755_46942# a_14035_46660# 0.040006f
C3288 a_n743_46660# a_1138_42852# 0.056829f
C3289 a_n2438_43548# a_1176_45822# 0.073092f
C3290 a_n2661_46634# a_3483_46348# 0.051915f
C3291 a_n1613_43370# a_2324_44458# 0.027159f
C3292 a_12891_46348# a_10903_43370# 0.132903f
C3293 a_22527_39145# a_22629_38406# 0.123152f
C3294 a_22581_37893# a_22944_39857# 0.011943f
C3295 a_22589_40055# a_22725_38406# 0.010302f
C3296 a_22537_40625# a_22725_37990# 0.010408f
C3297 a_22589_40599# a_22737_37285# 0.010048f
C3298 a_n4064_37984# VREF_GND 0.047292f
C3299 a_22889_38993# a_22537_39537# 0.033924f
C3300 a_13249_42308# a_13565_43940# 0.048533f
C3301 a_11691_44458# a_18443_44721# 0.042634f
C3302 a_n1925_42282# a_743_42282# 0.052333f
C3303 a_1307_43914# a_11967_42832# 0.031135f
C3304 a_n971_45724# a_3232_43370# 0.058382f
C3305 a_3160_47472# a_413_45260# 0.208121f
C3306 a_2107_46812# a_9049_44484# 0.240008f
C3307 a_n881_46662# a_16115_45572# 0.033547f
C3308 a_n1435_47204# a_3357_43084# 1.08491f
C3309 a_16327_47482# a_20528_45572# 0.011969f
C3310 a_5164_46348# a_5497_46414# 0.203417f
C3311 a_n2293_46098# a_2324_44458# 0.018455f
C3312 a_3483_46348# a_8199_44636# 1.81719f
C3313 a_3090_45724# a_13259_45724# 0.261789f
C3314 a_13487_47204# a_2437_43646# 0.014506f
C3315 a_11453_44696# a_16147_45260# 0.026325f
C3316 a_1847_42826# a_1606_42308# 0.025123f
C3317 a_743_42282# a_9803_42558# 0.010183f
C3318 a_13249_42308# a_5534_30871# 0.215947f
C3319 a_11967_42832# a_18579_44172# 0.158329f
C3320 a_5111_44636# a_9145_43396# 0.057312f
C3321 a_n2661_42834# a_2127_44172# 0.019594f
C3322 a_20640_44752# a_20766_44850# 0.17072f
C3323 a_20362_44736# a_19279_43940# 0.039759f
C3324 a_20679_44626# a_20835_44721# 0.105995f
C3325 a_11459_47204# VDD 0.34771f
C3326 a_6851_47204# DATA[3] 0.146601f
C3327 a_12465_44636# a_12607_44458# 0.186652f
C3328 a_10903_43370# a_11322_45546# 0.313957f
C3329 a_n1613_43370# a_n1699_44726# 0.166123f
C3330 a_5257_43370# a_1307_43914# 0.020655f
C3331 a_13747_46662# a_11827_44484# 0.044822f
C3332 a_18525_43370# VDD 0.263553f
C3333 a_14955_43940# a_15301_44260# 0.013377f
C3334 a_1414_42308# a_n97_42460# 0.196768f
C3335 a_22223_43948# a_15493_43940# 0.051823f
C3336 a_n2293_43922# a_12281_43396# 0.147288f
C3337 a_3090_45724# a_n2661_43922# 0.044809f
C3338 a_11525_45546# a_11778_45572# 0.011913f
C3339 a_4883_46098# a_12891_46348# 0.085714f
C3340 a_n237_47217# a_3877_44458# 0.059355f
C3341 a_3160_47472# a_2609_46660# 0.018687f
C3342 a_2905_45572# a_3177_46902# 0.014554f
C3343 a_13507_46334# a_768_44030# 0.019457f
C3344 a_10227_46804# a_5807_45002# 0.262866f
C3345 a_18057_42282# a_18310_42308# 0.011913f
C3346 a_21356_42826# VDD 0.225688f
C3347 a_14021_43940# a_14209_32519# 0.042544f
C3348 a_6197_43396# a_7287_43370# 0.041762f
C3349 a_6765_43638# a_6547_43396# 0.209641f
C3350 a_n913_45002# a_21335_42336# 0.062808f
C3351 a_n863_45724# VDD 1.89058f
C3352 a_n1059_45260# a_5111_44636# 0.038143f
C3353 a_n1613_43370# a_n2157_42858# 0.303592f
C3354 a_13249_42308# a_11691_44458# 0.017891f
C3355 a_9049_44484# a_n2661_44458# 0.015549f
C3356 a_10227_46804# a_10518_42984# 0.225803f
C3357 a_19692_46634# a_21845_43940# 0.014352f
C3358 a_8145_46902# a_8492_46660# 0.051162f
C3359 a_4791_45118# a_2324_44458# 0.19212f
C3360 a_5807_45002# a_17339_46660# 0.02927f
C3361 a_n4064_40160# VDD 2.37407f
C3362 VDAC_Ni a_3754_38470# 0.911632f
C3363 a_n3565_39304# C6_P_btm 0.080378f
C3364 a_13258_32519# VREF_GND 0.033872f
C3365 a_7754_39964# a_3726_37500# 0.030605f
C3366 a_7754_40130# a_5088_37509# 0.036831f
C3367 a_7174_31319# VIN_P 0.022822f
C3368 a_n1641_43230# a_n1545_43230# 0.013793f
C3369 a_8191_45002# VDD 0.39677f
C3370 a_n3674_39768# a_n3674_37592# 0.024722f
C3371 a_10193_42453# a_17973_43940# 0.084505f
C3372 a_3232_43370# a_9313_44734# 0.11426f
C3373 a_2382_45260# a_n2661_42834# 0.055134f
C3374 a_n2661_43370# a_n2129_44697# 0.014856f
C3375 a_n881_46662# a_6511_45714# 0.149116f
C3376 a_20820_30879# a_12741_44636# 0.103478f
C3377 a_3090_45724# a_18189_46348# 0.029136f
C3378 a_10227_46804# a_15143_45578# 0.010124f
C3379 a_18083_42858# a_19339_43156# 0.042271f
C3380 a_7871_42858# a_8292_43218# 0.086377f
C3381 a_4520_42826# a_4649_42852# 0.062574f
C3382 a_18989_43940# a_18579_44172# 0.035827f
C3383 a_18443_44721# a_18753_44484# 0.013793f
C3384 a_742_44458# a_1414_42308# 0.052151f
C3385 a_n2956_39768# a_n3565_39590# 0.302561f
C3386 a_n2661_46634# a_11963_45334# 0.036874f
C3387 a_18597_46090# a_16922_45042# 0.028931f
C3388 a_18819_46122# a_19240_46482# 0.089677f
C3389 a_8199_44636# a_n357_42282# 0.023438f
C3390 a_12861_44030# a_11691_44458# 0.196929f
C3391 a_2609_46660# a_413_45260# 0.022446f
C3392 a_16327_47482# a_18494_42460# 0.083754f
C3393 a_3090_45724# a_17478_45572# 0.128299f
C3394 a_3540_43646# VDD 0.209044f
C3395 a_2982_43646# RST_Z 0.015013f
C3396 a_16922_45042# a_743_42282# 0.120316f
C3397 a_n863_45724# a_n784_42308# 0.358682f
C3398 a_5072_46660# VDD 0.081835f
C3399 a_167_45260# a_1423_45028# 0.123079f
C3400 a_2711_45572# a_8746_45002# 0.010166f
C3401 a_6598_45938# a_6812_45938# 0.097745f
C3402 a_6667_45809# a_7230_45938# 0.049827f
C3403 a_526_44458# a_3357_43084# 0.04478f
C3404 a_n1613_43370# a_n1761_44111# 0.148121f
C3405 a_n443_42852# a_13249_42308# 0.033352f
C3406 a_12861_44030# a_18479_47436# 0.065796f
C3407 a_15673_47210# a_16327_47482# 0.206019f
C3408 a_15507_47210# a_16763_47508# 0.043475f
C3409 a_n237_47217# a_8128_46384# 0.113499f
C3410 a_n4318_38216# a_n4064_39616# 0.024304f
C3411 a_n3674_38216# a_n3420_39616# 0.02009f
C3412 a_11551_42558# a_11633_42558# 0.171361f
C3413 a_20193_45348# a_22165_42308# 0.252856f
C3414 a_15493_43396# a_15681_43442# 0.029338f
C3415 a_11967_42832# a_13635_43156# 0.053949f
C3416 a_18597_46090# a_15743_43084# 0.023066f
C3417 a_16327_47482# a_16388_46812# 0.01513f
C3418 a_12861_44030# a_17829_46910# 0.058114f
C3419 a_11453_44696# a_19333_46634# 0.026664f
C3420 a_2443_46660# a_3177_46902# 0.053479f
C3421 a_8685_42308# VDD 0.286875f
C3422 a_5742_30871# C1_N_btm 0.026156f
C3423 a_5932_42308# VIN_P 0.023512f
C3424 a_15743_43084# a_743_42282# 0.029529f
C3425 a_19700_43370# a_4190_30871# 0.046581f
C3426 a_5147_45002# a_n2661_44458# 0.024256f
C3427 a_413_45260# a_2779_44458# 0.024142f
C3428 a_n2956_39304# a_n4318_39304# 0.023717f
C3429 a_12861_44030# a_n443_42852# 0.015171f
C3430 SMPL_ON_N a_20205_31679# 0.029367f
C3431 a_n2293_46634# a_526_44458# 0.579444f
C3432 C0_dummy_N_btm C0_N_btm 7.97415f
C3433 C10_P_btm VDD 2.40001f
C3434 a_16979_44734# VDD 0.256327f
C3435 a_20692_30879# a_14209_32519# 0.051612f
C3436 a_5343_44458# a_n2661_42834# 0.038788f
C3437 a_19778_44110# a_19279_43940# 0.020911f
C3438 a_8975_43940# a_9313_44734# 0.391938f
C3439 a_5497_46414# a_5066_45546# 0.05403f
C3440 a_765_45546# a_n357_42282# 0.209746f
C3441 a_18819_46122# a_19553_46090# 0.052547f
C3442 a_2324_44458# a_6945_45028# 0.183081f
C3443 a_2455_43940# VDD 0.144352f
C3444 a_n699_43396# a_n97_42460# 0.152094f
C3445 a_n1059_45260# a_791_42968# 0.122941f
C3446 a_n913_45002# a_685_42968# 0.015577f
C3447 a_n2017_45002# a_1847_42826# 0.017915f
C3448 a_644_44056# a_1115_44172# 0.013441f
C3449 a_9804_47204# DATA[4] 0.015379f
C3450 a_8953_45546# a_9803_42558# 0.031932f
C3451 a_310_45028# a_n443_42852# 0.376934f
C3452 a_13059_46348# a_14797_45144# 0.066603f
C3453 a_20820_30879# a_413_45260# 0.033659f
C3454 a_13507_46334# a_17517_44484# 0.018934f
C3455 a_n357_42282# a_509_45822# 0.039776f
C3456 a_10586_45546# a_11652_45724# 0.046802f
C3457 a_16327_47482# a_20640_44752# 0.044807f
C3458 a_2905_45572# a_3160_47472# 0.54473f
C3459 a_n971_45724# a_6491_46660# 0.011282f
C3460 a_2952_47436# a_n1151_42308# 0.068429f
C3461 a_n237_47217# a_6151_47436# 0.360224f
C3462 a_n1741_47186# a_9067_47204# 0.012401f
C3463 a_7765_42852# VDD 0.333322f
C3464 a_5342_30871# C8_P_btm 0.093874f
C3465 a_1755_42282# a_6481_42558# 0.012532f
C3466 a_5534_30871# C6_P_btm 0.01116f
C3467 a_14539_43914# a_16795_42852# 0.037061f
C3468 a_2202_46116# VDD 0.20904f
C3469 a_5891_43370# a_7227_42852# 0.129383f
C3470 a_n2661_42282# a_6031_43396# 0.036698f
C3471 a_310_45028# a_375_42282# 0.078376f
C3472 a_n2293_45546# a_2304_45348# 0.032829f
C3473 a_n2956_38680# a_n4318_40392# 0.024261f
C3474 a_7499_43078# a_n913_45002# 0.548687f
C3475 a_n1613_43370# a_n2267_43396# 0.04778f
C3476 a_n863_45724# a_1423_45028# 0.113534f
C3477 a_n1151_42308# a_12991_46634# 0.013856f
C3478 a_6151_47436# a_8270_45546# 0.142873f
C3479 a_768_44030# a_n743_46660# 0.028134f
C3480 a_n1613_43370# a_491_47026# 0.038998f
C3481 a_4958_30871# a_n3420_37984# 0.031033f
C3482 a_n1794_35082# a_18194_34908# 0.466071f
C3483 a_n2302_39866# a_n2216_39866# 0.011479f
C3484 a_3539_42460# a_743_42282# 0.054149f
C3485 a_11823_42460# VDD 4.44574f
C3486 a_n2956_37592# a_n4064_37984# 0.012393f
C3487 a_3422_30871# a_20922_43172# 0.045027f
C3488 a_4927_45028# a_5365_45348# 0.013015f
C3489 a_10193_42453# a_9313_44734# 0.078654f
C3490 a_20692_30879# a_17730_32519# 0.05146f
C3491 a_3090_45724# a_14955_43396# 0.07523f
C3492 a_6755_46942# a_13885_46660# 0.078788f
C3493 a_n2497_47436# a_n863_45724# 0.337007f
C3494 a_n743_46660# a_1176_45822# 0.08607f
C3495 a_7754_39632# RST_Z 0.030938f
C3496 a_22589_40055# a_22629_38406# 0.1922f
C3497 a_n3420_37984# VCM 0.014539f
C3498 a_22581_37893# a_22848_39857# 0.01318f
C3499 a_22613_38993# a_22537_39537# 0.049665f
C3500 a_22537_40625# a_22629_37990# 0.130478f
C3501 a_n1059_45260# a_3905_42865# 0.01898f
C3502 a_11691_44458# a_18287_44626# 0.032949f
C3503 a_742_44458# a_n699_43396# 0.047576f
C3504 a_526_44458# a_743_42282# 0.042759f
C3505 a_2905_45572# a_413_45260# 0.124898f
C3506 a_n881_46662# a_16333_45814# 0.04285f
C3507 a_584_46384# a_2382_45260# 0.185451f
C3508 a_16327_47482# a_21188_45572# 0.227468f
C3509 a_3877_44458# a_4099_45572# 0.01632f
C3510 a_5164_46348# a_5204_45822# 0.132894f
C3511 a_12861_44030# a_2437_43646# 0.022753f
C3512 a_5649_42852# a_5934_30871# 0.058776f
C3513 a_743_42282# a_9223_42460# 0.010592f
C3514 a_n1644_44306# VDD 0.082968f
C3515 a_n2661_43370# a_n2433_43396# 0.021188f
C3516 a_9313_45822# VDD 0.5747f
C3517 a_6151_47436# DATA[5] 0.19492f
C3518 a_6491_46660# DATA[3] 0.011549f
C3519 a_n2661_42834# a_453_43940# 0.04708f
C3520 a_20362_44736# a_20766_44850# 0.051162f
C3521 a_n2661_43922# a_1414_42308# 0.010195f
C3522 a_20640_44752# a_20835_44721# 0.20669f
C3523 a_20159_44458# a_19279_43940# 0.06519f
C3524 a_8270_45546# a_5111_44636# 0.035253f
C3525 a_n1613_43370# a_n2267_44484# 0.025052f
C3526 a_6945_45028# a_6667_45809# 0.015851f
C3527 a_10903_43370# a_10490_45724# 0.057318f
C3528 a_13747_46662# a_21359_45002# 0.060042f
C3529 a_13661_43548# a_11827_44484# 0.120515f
C3530 a_13678_32519# EN_VIN_BSTR_N 0.031831f
C3531 a_18429_43548# VDD 0.163446f
C3532 a_22400_42852# COMP_P 0.595635f
C3533 a_n2840_42282# a_n3674_38680# 0.154001f
C3534 a_1467_44172# a_n97_42460# 0.190191f
C3535 a_3422_30871# a_2982_43646# 0.140944f
C3536 a_11341_43940# a_15493_43940# 0.216602f
C3537 a_9313_44734# a_16137_43396# 0.044229f
C3538 a_n2956_38680# a_n4209_38502# 0.235751f
C3539 a_12891_46348# a_13483_43940# 0.062818f
C3540 a_12549_44172# a_12429_44172# 0.137881f
C3541 a_3090_45724# a_n2661_42834# 0.164804f
C3542 a_11525_45546# a_11688_45572# 0.011381f
C3543 a_4185_45028# a_11827_44484# 0.03083f
C3544 a_526_44458# a_626_44172# 0.180416f
C3545 a_4883_46098# a_11309_47204# 0.012799f
C3546 a_16327_47482# a_19321_45002# 0.925259f
C3547 a_n971_45724# a_4646_46812# 0.303249f
C3548 a_3160_47472# a_2443_46660# 0.019074f
C3549 a_2905_45572# a_2609_46660# 0.027251f
C3550 a_12861_44030# a_n2661_46634# 0.03828f
C3551 a_13507_46334# a_12549_44172# 0.363125f
C3552 a_n1151_42308# a_n2661_46098# 0.024549f
C3553 a_18907_42674# a_19332_42282# 0.017308f
C3554 a_18057_42282# a_18220_42308# 0.01135f
C3555 a_18727_42674# a_18214_42558# 0.035505f
C3556 a_20922_43172# VDD 0.192467f
C3557 a_n1079_45724# VDD 0.172275f
C3558 a_n913_45002# a_7174_31319# 0.02792f
C3559 a_14021_43940# a_22591_43396# 0.057848f
C3560 a_6031_43396# a_7112_43396# 0.101963f
C3561 a_6197_43396# a_6547_43396# 0.216095f
C3562 a_3626_43646# a_3457_43396# 0.067226f
C3563 a_n2017_45002# a_5111_44636# 0.024598f
C3564 a_n37_45144# a_413_45260# 0.021944f
C3565 a_7499_43078# a_n2661_44458# 0.059442f
C3566 a_10227_46804# a_10083_42826# 0.292997f
C3567 a_2324_44458# a_895_43940# 0.011941f
C3568 a_n2312_39304# a_n2293_46098# 0.027561f
C3569 a_7577_46660# a_8492_46660# 0.118423f
C3570 a_4915_47217# a_14275_46494# 0.01257f
C3571 a_10227_46804# a_3483_46348# 0.057984f
C3572 a_7754_38636# a_3754_38470# 0.037604f
C3573 a_n4334_40480# VDD 0.390668f
C3574 a_7754_40130# a_4338_37500# 0.030623f
C3575 a_n1641_43230# a_n1736_43218# 0.049827f
C3576 a_9313_44734# a_22775_42308# 0.011571f
C3577 a_n4318_39768# a_n3674_37592# 0.024842f
C3578 a_7705_45326# VDD 0.211554f
C3579 a_10193_42453# a_17737_43940# 0.02461f
C3580 a_526_44458# a_2813_43396# 0.013054f
C3581 a_20692_30879# a_17538_32519# 0.05141f
C3582 a_n2661_43370# a_n2433_44484# 0.018595f
C3583 a_16922_45042# a_20193_45348# 0.328274f
C3584 a_n2438_43548# a_n2661_45546# 0.065227f
C3585 a_n881_46662# a_6472_45840# 0.179318f
C3586 a_n1613_43370# a_6511_45714# 0.017587f
C3587 a_15559_46634# a_2324_44458# 0.012623f
C3588 a_11453_44696# a_7499_43078# 0.02227f
C3589 a_22591_46660# a_12741_44636# 0.0686f
C3590 a_3090_45724# a_17715_44484# 0.108364f
C3591 a_18083_42858# a_18599_43230# 0.113784f
C3592 a_949_44458# a_1115_44172# 0.016355f
C3593 a_742_44458# a_1467_44172# 0.018499f
C3594 a_3357_43084# a_3626_43646# 0.018539f
C3595 a_2443_46660# a_413_45260# 0.020902f
C3596 a_16327_47482# a_18184_42460# 0.168018f
C3597 a_3090_45724# a_15861_45028# 0.125763f
C3598 a_13661_43548# a_15595_45028# 0.214904f
C3599 a_2982_43646# VDD 1.40372f
C3600 a_20193_45348# a_15743_43084# 0.060559f
C3601 a_n2293_42834# a_n1076_43230# 0.01241f
C3602 a_n2956_38216# a_n3674_37592# 0.025763f
C3603 a_6540_46812# VDD 0.084698f
C3604 a_13747_46662# a_19279_43940# 0.048937f
C3605 a_10903_43370# a_6171_45002# 0.041534f
C3606 a_2711_45572# a_10193_42453# 0.218272f
C3607 a_6511_45714# a_7230_45938# 0.088127f
C3608 a_6667_45809# a_6812_45938# 0.057222f
C3609 a_2324_44458# a_3065_45002# 0.017588f
C3610 a_3483_46348# a_1307_43914# 0.095243f
C3611 a_n1613_43370# a_n2065_43946# 0.30437f
C3612 a_15673_47210# a_16241_47178# 0.183195f
C3613 a_15811_47375# a_16327_47482# 0.038827f
C3614 a_12861_44030# a_18143_47464# 0.394543f
C3615 a_15507_47210# a_16023_47582# 0.109156f
C3616 COMP_P a_n4209_39590# 0.010869f
C3617 a_n913_45002# a_5932_42308# 0.220872f
C3618 a_15493_43940# a_10341_43396# 0.051273f
C3619 a_11967_42832# a_12895_43230# 0.035759f
C3620 a_15682_43940# a_16243_43396# 0.013782f
C3621 a_n1151_42308# a_n901_43156# 0.01984f
C3622 a_20692_30879# a_19721_31679# 0.051673f
C3623 a_n2293_46634# a_3626_43646# 0.012347f
C3624 a_n971_45724# a_n901_46420# 0.021388f
C3625 a_11453_44696# a_15227_44166# 0.979188f
C3626 a_12861_44030# a_765_45546# 0.190301f
C3627 a_2443_46660# a_2609_46660# 0.579196f
C3628 a_8325_42308# VDD 0.313956f
C3629 a_n3565_39590# a_n4209_37414# 0.031279f
C3630 a_n4209_39590# a_n3565_37414# 0.032656f
C3631 a_5742_30871# C0_N_btm 0.014563f
C3632 a_n4064_40160# a_n4064_37440# 0.056406f
C3633 a_n3420_38528# a_n4064_37984# 7.35343f
C3634 a_n4064_38528# a_n3420_37984# 0.044626f
C3635 a_n2946_38778# a_n2946_37984# 0.052227f
C3636 a_19268_43646# a_4190_30871# 0.035721f
C3637 a_3626_43646# a_5342_30871# 0.08847f
C3638 a_n356_44636# a_5742_30871# 0.120133f
C3639 a_18597_46090# a_21195_42852# 0.01512f
C3640 a_413_45260# a_949_44458# 0.018785f
C3641 a_4791_45118# a_6511_45714# 0.034343f
C3642 a_10227_46804# a_n357_42282# 0.103631f
C3643 a_16388_46812# a_16721_46634# 0.222024f
C3644 a_21753_35474# VDD 0.525301f
C3645 a_14539_43914# VDD 0.873589f
C3646 a_2982_43646# a_n784_42308# 0.026817f
C3647 a_20205_31679# a_14209_32519# 0.051418f
C3648 a_n699_43396# a_n2661_43922# 0.053529f
C3649 a_11827_44484# a_11967_42832# 0.095859f
C3650 a_10057_43914# a_9313_44734# 0.139382f
C3651 a_7499_43078# a_9145_43396# 0.040441f
C3652 a_5204_45822# a_5066_45546# 0.402457f
C3653 a_n881_46662# a_n745_45366# 0.152998f
C3654 a_4883_46098# a_6171_45002# 0.020043f
C3655 a_11599_46634# a_15415_45028# 0.013635f
C3656 a_8953_45546# a_526_44458# 0.037032f
C3657 a_18819_46122# a_18985_46122# 0.749955f
C3658 a_765_45546# a_310_45028# 0.012232f
C3659 a_2253_43940# VDD 0.156797f
C3660 a_n699_43396# a_n447_43370# 0.040315f
C3661 a_n1059_45260# a_685_42968# 0.103646f
C3662 a_9313_44734# a_14021_43940# 0.014591f
C3663 a_8953_45546# a_9223_42460# 0.166987f
C3664 a_3316_45546# a_3503_45724# 0.024901f
C3665 a_310_45028# a_509_45822# 0.039722f
C3666 a_n1099_45572# a_n443_42852# 0.026572f
C3667 a_10586_45546# a_11525_45546# 0.115475f
C3668 a_13059_46348# a_14537_43396# 0.30244f
C3669 a_584_46384# a_453_43940# 0.125447f
C3670 a_768_44030# a_5891_43370# 0.050862f
C3671 a_16327_47482# a_20362_44736# 0.213851f
C3672 a_5066_45546# a_8697_45822# 0.033513f
C3673 a_7871_42858# VDD 0.395222f
C3674 a_n971_45724# a_6545_47178# 0.295443f
C3675 a_2952_47436# a_3160_47472# 0.192116f
C3676 a_n1741_47186# a_6575_47204# 0.075265f
C3677 a_5534_30871# C7_P_btm 0.060228f
C3678 a_5267_42460# a_5379_42460# 0.156424f
C3679 a_3318_42354# a_3581_42558# 0.011552f
C3680 a_1755_42282# a_5932_42308# 0.046344f
C3681 a_14021_43940# a_20974_43370# 0.893848f
C3682 a_5891_43370# a_5755_42852# 0.160849f
C3683 a_1823_45246# VDD 1.7584f
C3684 a_n2956_39304# a_n4318_40392# 0.023379f
C3685 a_12741_44636# a_n2293_43922# 0.114756f
C3686 a_n357_42282# a_1307_43914# 0.044512f
C3687 a_2324_44458# a_6298_44484# 0.315008f
C3688 a_7499_43078# a_n1059_45260# 0.277353f
C3689 a_n1613_43370# a_n2129_43609# 0.44294f
C3690 a_2747_46873# a_2959_46660# 0.010672f
C3691 a_12549_44172# a_n743_46660# 0.03191f
C3692 a_4883_46098# a_4955_46873# 0.09516f
C3693 a_n1613_43370# a_288_46660# 0.01808f
C3694 a_n4064_40160# a_n3420_39072# 0.052668f
C3695 a_n4209_39590# a_n4209_39304# 0.045123f
C3696 a_n4315_30879# a_n4064_39072# 0.036792f
C3697 a_2982_43646# a_21487_43396# 0.169809f
C3698 a_3626_43646# a_743_42282# 0.147999f
C3699 a_12427_45724# VDD 0.33808f
C3700 a_n913_45002# a_n2661_43370# 0.031604f
C3701 a_20205_31679# a_17730_32519# 0.051307f
C3702 a_13556_45296# a_14537_43396# 0.590856f
C3703 a_2680_45002# a_2809_45028# 0.062574f
C3704 a_11309_47204# a_11387_46155# 0.061891f
C3705 a_n743_46660# a_1208_46090# 0.045297f
C3706 a_n2293_46634# a_167_45260# 0.087596f
C3707 SMPL_ON_P a_n2810_45572# 0.039568f
C3708 a_171_46873# a_376_46348# 0.080253f
C3709 a_768_44030# a_9290_44172# 0.189655f
C3710 a_7754_39632# VDD 0.205733f
C3711 a_n3420_37984# VREF_GND 0.047887f
C3712 a_22581_37893# a_22537_39537# 1.00904f
C3713 a_22613_38993# a_22889_38993# 0.237336f
C3714 a_22589_40599# a_22629_37990# 0.021352f
C3715 a_n2661_43370# CLK 0.011991f
C3716 a_4905_42826# a_5193_42852# 0.016389f
C3717 a_14309_45028# VDD 0.189806f
C3718 a_8199_44636# a_9127_43156# 0.01079f
C3719 a_n2293_42834# a_n2293_43922# 0.031735f
C3720 a_11691_44458# a_18248_44752# 0.040333f
C3721 a_18184_42460# a_n356_44636# 0.05602f
C3722 a_11827_44484# a_18989_43940# 0.054716f
C3723 a_3483_46348# a_8016_46348# 0.019798f
C3724 a_2952_47436# a_413_45260# 0.026401f
C3725 a_n1151_42308# a_n467_45028# 0.406349f
C3726 a_16327_47482# a_21363_45546# 0.276554f
C3727 a_5068_46348# a_5204_45822# 0.20685f
C3728 a_4646_46812# a_2711_45572# 0.053113f
C3729 a_13717_47436# a_2437_43646# 0.085485f
C3730 a_n881_46662# a_15765_45572# 0.58719f
C3731 a_17595_43084# a_17749_42852# 0.010303f
C3732 a_n3674_39768# VDD 0.398971f
C3733 a_13249_42308# a_13460_43230# 0.014543f
C3734 a_11031_47542# VDD 0.214104f
C3735 a_6545_47178# DATA[3] 0.178561f
C3736 a_5891_43370# a_7845_44172# 0.119969f
C3737 a_4915_47217# CLK 0.198293f
C3738 a_n2661_42834# a_1414_42308# 0.081864f
C3739 a_20640_44752# a_20679_44626# 0.582607f
C3740 a_n2293_42834# a_n97_42460# 0.17628f
C3741 a_n1151_42308# a_n2661_43922# 0.056653f
C3742 a_15227_44166# a_n1059_45260# 0.099892f
C3743 a_2107_46812# a_n2661_43370# 0.02614f
C3744 a_n1613_43370# a_n2129_44697# 0.026334f
C3745 a_6945_45028# a_6511_45714# 0.028815f
C3746 a_n1925_42282# a_n443_42852# 0.02261f
C3747 a_9290_44172# a_11652_45724# 0.020364f
C3748 a_11189_46129# a_11525_45546# 0.085926f
C3749 a_12005_46116# a_10193_42453# 0.016165f
C3750 a_13747_46662# a_21101_45002# 0.081818f
C3751 a_5807_45002# a_11827_44484# 0.022597f
C3752 a_19321_45002# a_20567_45036# 0.205038f
C3753 a_17324_43396# VDD 0.274722f
C3754 a_11341_43940# a_22223_43948# 0.175191f
C3755 a_21115_43940# a_15493_43940# 0.0516f
C3756 a_2711_45572# a_18479_45785# 0.032371f
C3757 a_12465_44636# a_14021_43940# 0.015806f
C3758 a_n2312_38680# a_n3674_39768# 0.023176f
C3759 a_n2840_45546# a_n2840_45002# 0.026152f
C3760 a_n971_45724# a_3877_44458# 0.927248f
C3761 a_2905_45572# a_2443_46660# 0.026052f
C3762 a_13507_46334# a_12891_46348# 0.076674f
C3763 a_16588_47582# a_5807_45002# 0.040789f
C3764 a_18057_42282# a_18214_42558# 0.18824f
C3765 a_19987_42826# VDD 0.588466f
C3766 a_n2293_45546# VDD 2.06545f
C3767 a_14021_43940# a_13887_32519# 0.020984f
C3768 a_6197_43396# a_6765_43638# 0.17072f
C3769 a_6031_43396# a_7287_43370# 0.042271f
C3770 a_4185_45028# a_n2661_42282# 0.833759f
C3771 a_19692_46634# a_20974_43370# 0.012779f
C3772 a_13259_45724# a_13857_44734# 0.03212f
C3773 a_2324_44458# a_2479_44172# 0.010173f
C3774 a_9313_45822# a_9569_46155# 0.019679f
C3775 a_8145_46902# a_7927_46660# 0.209641f
C3776 a_7577_46660# a_8667_46634# 0.041879f
C3777 a_13258_32519# VIN_N 0.137523f
C3778 a_n4315_30879# VDD 4.04834f
C3779 a_7754_40130# a_3726_37500# 0.021358f
C3780 a_6709_45028# VDD 0.390566f
C3781 a_19778_44110# a_21005_45260# 0.135527f
C3782 a_20205_31679# a_17538_32519# 0.051233f
C3783 a_n2661_43370# a_n2661_44458# 1.0558f
C3784 a_16922_45042# a_11691_44458# 0.428229f
C3785 a_2711_45572# a_14021_43940# 0.029672f
C3786 a_n2293_42834# a_742_44458# 0.039916f
C3787 a_4883_46098# a_8746_45002# 0.032616f
C3788 a_10227_46804# a_13249_42308# 0.064815f
C3789 a_n743_46660# a_n2661_45546# 0.013544f
C3790 a_n881_46662# a_6194_45824# 0.063172f
C3791 a_n1613_43370# a_6472_45840# 0.017909f
C3792 a_n2293_46634# a_n863_45724# 0.157683f
C3793 a_22591_46660# a_20820_30879# 0.166885f
C3794 a_11415_45002# a_12741_44636# 1.07921f
C3795 a_7227_42852# a_7573_43172# 0.013377f
C3796 a_n913_45002# a_1568_43370# 0.098659f
C3797 a_n2956_39768# a_n4209_39590# 0.334714f
C3798 a_n2312_38680# a_n4315_30879# 0.024522f
C3799 a_n2442_46660# a_n2302_40160# 0.017419f
C3800 a_167_45260# a_2277_45546# 0.214157f
C3801 a_n1151_42308# a_n452_44636# 0.238824f
C3802 a_17957_46116# a_16375_45002# 0.017118f
C3803 a_16327_47482# a_19778_44110# 0.037655f
C3804 a_3090_45724# a_8696_44636# 0.038457f
C3805 a_13661_43548# a_15415_45028# 0.133591f
C3806 a_2896_43646# VDD 0.208317f
C3807 a_n2293_42282# a_n3674_38216# 0.111055f
C3808 a_5732_46660# VDD 0.277366f
C3809 a_16922_45042# a_4190_30871# 0.353708f
C3810 a_n2293_42834# a_n901_43156# 0.021108f
C3811 a_n2293_43922# a_n2012_43396# 0.011692f
C3812 a_19321_45002# a_20679_44626# 0.023087f
C3813 a_10903_43370# a_3232_43370# 0.114259f
C3814 a_167_45260# a_626_44172# 0.04273f
C3815 a_2711_45572# a_10180_45724# 0.01318f
C3816 a_6472_45840# a_7230_45938# 0.05936f
C3817 a_8953_45546# a_8953_45002# 0.023516f
C3818 a_1823_45246# a_1423_45028# 0.024089f
C3819 a_8199_44636# a_10951_45334# 0.237774f
C3820 a_4915_47217# a_11453_44696# 0.026396f
C3821 a_12861_44030# a_10227_46804# 0.291378f
C3822 a_15507_47210# a_16327_47482# 0.425757f
C3823 a_n1741_47186# a_12891_46348# 0.107238f
C3824 a_n971_45724# a_8128_46384# 0.041637f
C3825 a_n4318_38216# a_n3420_39616# 0.023792f
C3826 a_n3674_38680# a_n4064_39616# 0.019915f
C3827 a_1606_42308# a_7174_31319# 2.41314f
C3828 a_11967_42832# a_13113_42826# 0.021992f
C3829 a_n913_45002# a_6171_42473# 0.034189f
C3830 a_20205_31679# a_19721_31679# 0.052217f
C3831 a_20692_30879# a_18114_32519# 0.051555f
C3832 a_13249_42308# a_1307_43914# 0.056917f
C3833 a_n2497_47436# a_1823_45246# 0.025359f
C3834 a_11453_44696# a_18834_46812# 0.010577f
C3835 a_12861_44030# a_17339_46660# 1.25428f
C3836 a_n1925_46634# a_5907_46634# 0.010645f
C3837 a_13258_32519# CAL_N 0.020535f
C3838 a_2112_39137# a_2113_38308# 0.478223f
C3839 a_n2293_43922# a_5379_42460# 0.4571f
C3840 a_15743_43084# a_4190_30871# 0.290729f
C3841 a_18799_45938# VDD 0.132317f
C3842 a_16751_45260# a_17023_45118# 0.13675f
C3843 a_13259_45724# a_15493_43940# 0.019228f
C3844 a_10193_42453# a_20512_43084# 0.086337f
C3845 a_4791_45118# a_6472_45840# 0.025301f
C3846 a_19692_46634# a_20528_46660# 0.021985f
C3847 a_17609_46634# a_18280_46660# 0.094543f
C3848 a_5257_43370# a_6419_46155# 0.186651f
C3849 C0_dummy_P_btm C0_dummy_N_btm 0.033338f
C3850 C7_P_btm C7_N_btm 0.028901f
C3851 C6_P_btm C6_N_btm 0.019861f
C3852 C5_P_btm C5_N_btm 0.03705f
C3853 C4_P_btm C4_N_btm 0.02642f
C3854 C3_P_btm C3_N_btm 2.90911f
C3855 C2_P_btm C2_N_btm 0.026726f
C3856 C1_P_btm C1_N_btm 0.065833f
C3857 C0_P_btm C0_N_btm 0.044249f
C3858 a_19998_34978# VDD 0.319197f
C3859 a_n1557_42282# a_n1794_35082# 0.865968f
C3860 a_16112_44458# VDD 0.182397f
C3861 a_14579_43548# a_14635_42282# 0.124652f
C3862 a_20692_30879# a_13887_32519# 0.051577f
C3863 a_n699_43396# a_n2661_42834# 0.131393f
C3864 a_4223_44672# a_n2661_43922# 0.059715f
C3865 a_n863_45724# a_743_42282# 0.05133f
C3866 a_10440_44484# a_9313_44734# 0.027369f
C3867 a_n443_42852# a_15743_43084# 0.034562f
C3868 a_5164_46348# a_5066_45546# 0.096188f
C3869 a_n1613_43370# a_n745_45366# 0.012092f
C3870 a_4883_46098# a_3232_43370# 0.017979f
C3871 a_12861_44030# a_1307_43914# 0.038753f
C3872 a_11415_45002# a_16375_45002# 0.080382f
C3873 a_12741_44636# a_13259_45724# 0.113445f
C3874 a_8270_45546# a_7499_43078# 0.063428f
C3875 a_1443_43940# VDD 0.144342f
C3876 a_10341_42308# a_5742_30871# 0.031841f
C3877 a_13467_32519# a_22485_38105# 0.076404f
C3878 a_15928_47570# VDD 0.08228f
C3879 a_768_44030# RST_Z 0.05505f
C3880 a_8199_44636# a_9803_42558# 0.036259f
C3881 a_n1925_42282# COMP_P 0.071512f
C3882 a_n881_46662# CLK 0.023376f
C3883 a_3218_45724# a_3503_45724# 0.099872f
C3884 a_n1099_45572# a_509_45822# 0.026885f
C3885 a_380_45546# a_n443_42852# 0.030032f
C3886 a_10586_45546# a_11322_45546# 0.220166f
C3887 a_13059_46348# a_14180_45002# 0.073427f
C3888 a_12861_44030# a_18579_44172# 0.221909f
C3889 a_16327_47482# a_20159_44458# 0.270426f
C3890 a_584_46384# a_1414_42308# 0.321387f
C3891 a_n1151_42308# a_n809_44244# 0.02481f
C3892 a_11415_45002# a_413_45260# 0.063143f
C3893 a_7227_42852# VDD 0.254613f
C3894 a_2952_47436# a_2905_45572# 0.318161f
C3895 a_n971_45724# a_6151_47436# 0.29974f
C3896 a_2063_45854# a_n1151_42308# 0.425035f
C3897 a_3318_42354# a_3497_42558# 0.010303f
C3898 a_n1794_35082# a_5934_30871# 0.039258f
C3899 a_1755_42282# a_6171_42473# 0.065035f
C3900 a_1606_42308# a_5932_42308# 0.111585f
C3901 a_n2661_42834# a_n4318_38680# 0.102282f
C3902 a_18579_44172# a_19700_43370# 0.175511f
C3903 a_11967_42832# a_16823_43084# 0.093759f
C3904 a_14021_43940# a_14401_32519# 0.059818f
C3905 a_n2017_45002# a_18504_43218# 0.016191f
C3906 a_1138_42852# VDD 0.397518f
C3907 a_5257_43370# a_n2661_42282# 0.01339f
C3908 a_n2293_45546# a_1423_45028# 0.06244f
C3909 a_2324_44458# a_5518_44484# 0.112753f
C3910 a_7499_43078# a_n2017_45002# 0.065458f
C3911 a_n863_45724# a_626_44172# 0.097275f
C3912 a_10809_44734# a_n2661_44458# 0.033319f
C3913 a_10903_43370# a_8975_43940# 0.043009f
C3914 a_n1613_43370# a_n2433_43396# 0.299968f
C3915 a_n881_46662# a_2107_46812# 0.138703f
C3916 a_n1613_43370# a_1983_46706# 0.020434f
C3917 a_19321_45002# a_19594_46812# 0.267862f
C3918 a_12891_46348# a_n743_46660# 0.044305f
C3919 a_14097_32519# C4_N_btm 0.030945f
C3920 a_n1794_35082# a_10890_34112# 0.017188f
C3921 a_11962_45724# VDD 0.210594f
C3922 a_n97_42460# a_n13_43084# 0.13246f
C3923 a_n1059_45260# a_n2661_43370# 0.03635f
C3924 a_2382_45260# a_2809_45028# 0.034331f
C3925 a_3090_45724# a_14205_43396# 0.040425f
C3926 a_9482_43914# a_14537_43396# 0.040878f
C3927 a_5807_45002# a_6419_46155# 0.072498f
C3928 a_12991_46634# a_12816_46660# 0.233657f
C3929 a_n743_46660# a_805_46414# 0.064413f
C3930 a_n881_46662# a_14493_46090# 0.011925f
C3931 a_12549_44172# a_9290_44172# 0.053193f
C3932 a_11309_47204# a_11133_46155# 0.040357f
C3933 a_11453_44696# a_10809_44734# 0.274367f
C3934 a_n2497_47436# a_n2293_45546# 0.307373f
C3935 a_22537_40625# a_22629_38406# 0.066321f
C3936 a_n4064_37984# VIN_P 0.059416f
C3937 a_n3565_38216# VCM 0.03544f
C3938 a_22581_37893# a_22889_38993# 0.112329f
C3939 a_10922_42852# a_10341_42308# 0.053077f
C3940 a_n443_42852# a_3539_42460# 0.02291f
C3941 a_8953_45546# a_8037_42858# 0.017317f
C3942 a_22612_30879# a_14097_32519# 0.059759f
C3943 a_n755_45592# a_8147_43396# 0.134231f
C3944 a_n2293_42834# a_n2661_43922# 0.03113f
C3945 a_11691_44458# a_17970_44736# 0.040435f
C3946 a_n2661_44458# a_5883_43914# 0.010478f
C3947 a_3877_44458# a_2711_45572# 0.099631f
C3948 a_n2293_46634# a_11823_42460# 0.072996f
C3949 a_16327_47482# a_20623_45572# 0.168593f
C3950 a_5068_46348# a_5164_46348# 0.31819f
C3951 a_n1435_47204# a_2437_43646# 0.191468f
C3952 a_n971_45724# a_5111_44636# 0.381443f
C3953 a_n881_46662# a_15903_45785# 0.032602f
C3954 a_743_42282# a_8685_42308# 0.039566f
C3955 a_5649_42852# a_6123_31319# 0.062309f
C3956 a_17595_43084# a_17665_42852# 0.011552f
C3957 a_n4318_39768# VDD 0.469044f
C3958 a_11823_42460# a_5342_30871# 0.044603f
C3959 a_n2661_43370# a_n2840_43370# 0.172532f
C3960 a_11967_42832# a_19279_43940# 0.070262f
C3961 a_17517_44484# a_22315_44484# 0.063928f
C3962 a_n2661_42834# a_1467_44172# 0.028215f
C3963 a_20362_44736# a_20679_44626# 0.102355f
C3964 a_10193_42453# a_18249_42858# 0.038446f
C3965 a_9863_47436# VDD 0.207794f
C3966 a_6151_47436# DATA[3] 0.041263f
C3967 a_10903_43370# a_10193_42453# 0.402091f
C3968 a_11189_46129# a_11322_45546# 0.05577f
C3969 a_n1151_42308# a_n2661_42834# 0.038196f
C3970 a_n1613_43370# a_n2433_44484# 0.29864f
C3971 a_6945_45028# a_6472_45840# 0.034109f
C3972 a_526_44458# a_n443_42852# 2.06448f
C3973 a_13259_45724# a_16375_45002# 0.60955f
C3974 a_13747_46662# a_21005_45260# 0.058269f
C3975 a_19321_45002# a_18494_42460# 0.084551f
C3976 a_4883_46098# a_8975_43940# 0.018394f
C3977 a_17499_43370# VDD 0.453381f
C3978 a_20935_43940# a_15493_43940# 0.037795f
C3979 a_11322_45546# a_11136_45572# 0.044092f
C3980 a_n2312_38680# a_n4318_39768# 0.023285f
C3981 a_8049_45260# a_8191_45002# 0.084237f
C3982 a_17339_46660# a_18287_44626# 0.018815f
C3983 a_3483_46348# a_11827_44484# 0.060892f
C3984 a_n443_46116# a_2107_46812# 0.075963f
C3985 a_16327_47482# a_13747_46662# 0.128159f
C3986 a_16763_47508# a_5807_45002# 0.127783f
C3987 a_18727_42674# a_18907_42674# 0.185422f
C3988 a_19164_43230# VDD 0.278643f
C3989 a_2982_43646# a_3457_43396# 0.074308f
C3990 a_14021_43940# a_22223_43396# 0.028989f
C3991 a_6031_43396# a_6547_43396# 0.105995f
C3992 a_n2956_38216# VDD 0.484692f
C3993 a_n143_45144# a_n37_45144# 0.13675f
C3994 a_n913_45002# a_3537_45260# 0.148413f
C3995 a_20202_43084# a_15493_43940# 0.02138f
C3996 a_9313_45822# a_9625_46129# 0.018694f
C3997 a_7577_46660# a_7927_46660# 0.206455f
C3998 a_4915_47217# a_13925_46122# 0.029041f
C3999 a_7411_46660# a_8492_46660# 0.102325f
C4000 a_22485_38105# RST_Z 0.036748f
C4001 a_n4209_39304# C7_P_btm 0.184297f
C4002 a_n901_43156# a_n13_43084# 0.014329f
C4003 a_n1991_42858# a_n1736_43218# 0.064178f
C4004 a_16137_43396# a_18249_42858# 0.021561f
C4005 a_7229_43940# VDD 0.821851f
C4006 a_413_45260# a_n2661_43922# 0.031184f
C4007 a_18184_42460# a_18494_42460# 1.31047f
C4008 a_19778_44110# a_20567_45036# 0.044967f
C4009 a_7229_43940# a_7640_43914# 0.177622f
C4010 a_20692_30879# a_14401_32519# 0.054254f
C4011 a_n1613_43370# a_8495_42852# 0.012196f
C4012 a_4883_46098# a_10193_42453# 0.040505f
C4013 a_n881_46662# a_5907_45546# 0.070761f
C4014 a_14976_45028# a_2324_44458# 0.086305f
C4015 a_11415_45002# a_20820_30879# 0.056772f
C4016 a_20202_43084# a_12741_44636# 0.22243f
C4017 a_n2312_38680# a_n2956_38216# 0.044798f
C4018 a_9313_45822# a_9159_45572# 0.051702f
C4019 a_3626_43646# a_14113_42308# 0.077829f
C4020 a_n1059_45260# a_1568_43370# 0.011697f
C4021 a_18287_44626# a_18579_44172# 0.107662f
C4022 a_18989_43940# a_19279_43940# 0.053948f
C4023 a_11823_42460# a_743_42282# 0.147603f
C4024 a_3357_43084# a_2982_43646# 0.01988f
C4025 a_584_46384# a_n699_43396# 0.632931f
C4026 a_n443_46116# a_n2661_44458# 0.034876f
C4027 a_167_45260# a_1609_45822# 0.141505f
C4028 a_18189_46348# a_16375_45002# 0.165328f
C4029 a_17957_46116# a_18243_46436# 0.010132f
C4030 a_13661_43548# a_14797_45144# 0.116989f
C4031 a_n2293_42282# a_n2104_42282# 0.058363f
C4032 a_5907_46634# VDD 0.341121f
C4033 a_16922_45042# a_21259_43561# 0.108631f
C4034 a_20512_43084# a_14021_43940# 0.030282f
C4035 a_n2293_42834# a_n1641_43230# 0.014975f
C4036 a_19321_45002# a_20640_44752# 0.034599f
C4037 a_2711_45572# a_10053_45546# 0.018932f
C4038 a_6472_45840# a_6812_45938# 0.027606f
C4039 a_8199_44636# a_10775_45002# 0.064568f
C4040 a_5937_45572# a_8953_45002# 0.062333f
C4041 a_2324_44458# a_2382_45260# 0.044897f
C4042 a_12861_44030# a_17591_47464# 0.079093f
C4043 a_15811_47375# a_15673_47210# 0.281607f
C4044 a_15507_47210# a_16241_47178# 0.06628f
C4045 a_11599_46634# a_16327_47482# 0.526398f
C4046 a_n1741_47186# a_11309_47204# 0.01734f
C4047 a_6151_47436# a_12465_44636# 0.025929f
C4048 a_11323_42473# a_11551_42558# 0.062483f
C4049 a_11341_43940# a_10341_43396# 0.289072f
C4050 a_n1917_43396# a_n1821_43396# 0.013793f
C4051 a_11967_42832# a_12545_42858# 0.028062f
C4052 a_15493_43940# a_14955_43396# 0.013181f
C4053 a_n97_42460# a_104_43370# 0.027998f
C4054 a_n913_45002# a_5755_42308# 0.036226f
C4055 a_10809_44734# EN_OFFSET_CAL 0.035912f
C4056 a_20205_31679# a_18114_32519# 0.051478f
C4057 a_20623_45572# a_20731_45938# 0.057222f
C4058 a_2324_44458# a_15433_44458# 0.021739f
C4059 a_n2293_46634# a_2982_43646# 0.015801f
C4060 a_n2661_46098# a_2443_46660# 0.063999f
C4061 a_n2497_47436# a_1138_42852# 0.144386f
C4062 a_11453_44696# a_17609_46634# 0.079593f
C4063 a_15811_47375# a_16388_46812# 0.010369f
C4064 a_10227_46804# a_14035_46660# 0.035412f
C4065 a_n4315_30879# a_n4064_37440# 0.035563f
C4066 a_n4209_39590# a_n4209_37414# 0.031971f
C4067 a_n4064_40160# a_n3420_37440# 0.062634f
C4068 a_n4064_38528# a_n3565_38216# 0.028041f
C4069 a_n3565_38502# a_n4064_37984# 0.028083f
C4070 a_n3420_38528# a_n3420_37984# 0.113087f
C4071 a_2982_43646# a_5342_30871# 0.178973f
C4072 a_3626_43646# a_5534_30871# 0.082646f
C4073 a_18783_43370# a_4190_30871# 0.044615f
C4074 a_18596_45572# VDD 0.077608f
C4075 a_n2661_42282# a_n2293_42282# 1.04835f
C4076 a_3537_45260# a_n2661_44458# 0.056342f
C4077 a_16751_45260# a_16922_45042# 0.12103f
C4078 a_n755_45592# a_n2661_42282# 0.025718f
C4079 a_18597_46090# a_20922_43172# 0.021228f
C4080 a_6151_47436# a_2711_45572# 0.050517f
C4081 a_17609_46634# a_17639_46660# 0.094289f
C4082 a_5257_43370# a_6165_46155# 0.11382f
C4083 a_19250_34978# VDD 0.323729f
C4084 a_15004_44636# VDD 0.090175f
C4085 a_10334_44484# a_9313_44734# 0.018652f
C4086 a_20205_31679# a_13887_32519# 0.051379f
C4087 a_5518_44484# a_5708_44484# 0.045837f
C4088 a_4223_44672# a_n2661_42834# 0.031905f
C4089 a_n2661_44458# a_11541_44484# 0.053139f
C4090 a_2779_44458# a_n2661_43922# 0.013114f
C4091 a_10193_42453# a_8685_43396# 0.024858f
C4092 a_5068_46348# a_5066_45546# 0.04842f
C4093 a_n881_46662# a_n1059_45260# 0.121542f
C4094 a_2747_46873# a_413_45260# 0.038809f
C4095 a_n1613_43370# a_n913_45002# 0.686014f
C4096 a_8199_44636# a_526_44458# 0.019697f
C4097 a_765_45546# a_380_45546# 0.141908f
C4098 a_8270_45546# a_8568_45546# 0.015327f
C4099 a_1241_43940# VDD 0.162129f
C4100 a_n2293_43922# a_11341_43940# 0.026007f
C4101 a_n699_43396# a_n1177_43370# 0.060973f
C4102 a_768_44030# VDD 1.53454f
C4103 a_8199_44636# a_9223_42460# 0.065156f
C4104 a_8953_45546# a_8685_42308# 0.250058f
C4105 a_n1925_42282# a_n4318_37592# 0.024213f
C4106 a_768_44030# a_7640_43914# 0.036222f
C4107 a_3218_45724# a_3316_45546# 0.162813f
C4108 a_380_45546# a_509_45822# 0.062574f
C4109 a_8049_45260# a_11823_42460# 0.046281f
C4110 a_n863_45724# a_1609_45822# 0.117311f
C4111 a_n2293_46634# a_14539_43914# 0.045317f
C4112 a_8270_45546# a_n2661_43370# 0.022558f
C4113 a_1823_45246# a_3357_43084# 0.062163f
C4114 a_10586_45546# a_10490_45724# 0.235237f
C4115 a_584_46384# a_n1151_42308# 0.047349f
C4116 a_n1741_47186# a_7227_47204# 0.016018f
C4117 a_n237_47217# a_4915_47217# 0.071869f
C4118 a_5755_42852# VDD 0.179985f
C4119 a_21076_30879# VCM 0.097317f
C4120 a_n2661_42834# a_n3674_39304# 0.038671f
C4121 a_1176_45822# VDD 0.781481f
C4122 a_11823_42460# a_15051_42282# 0.367924f
C4123 a_14021_43940# a_21381_43940# 0.022437f
C4124 a_18597_46090# a_2982_43646# 0.239147f
C4125 a_12549_44172# a_19319_43548# 0.024381f
C4126 a_2324_44458# a_5343_44458# 0.255488f
C4127 a_10903_43370# a_10057_43914# 0.052284f
C4128 a_19692_46634# a_20512_43084# 0.387138f
C4129 a_n1613_43370# a_2107_46812# 0.05377f
C4130 a_2747_46873# a_2609_46660# 0.347674f
C4131 a_n1151_42308# a_11901_46660# 0.020194f
C4132 a_4883_46098# a_4646_46812# 0.028054f
C4133 a_9313_45822# a_6755_46942# 0.031706f
C4134 a_n2946_39866# a_n2860_39866# 0.011479f
C4135 a_n4064_39616# a_n2302_39866# 0.239588f
C4136 a_n4064_40160# a_n3565_39304# 0.028096f
C4137 a_n4315_30879# a_n3420_39072# 0.036979f
C4138 a_2982_43646# a_743_42282# 0.047135f
C4139 a_3626_43646# a_4190_30871# 0.070713f
C4140 a_11652_45724# VDD 0.155048f
C4141 a_13556_45296# a_13777_45326# 0.101558f
C4142 a_20273_45572# a_21101_45002# 0.014321f
C4143 a_n2017_45002# a_n2661_43370# 0.038361f
C4144 a_9049_44484# a_9313_44734# 0.034936f
C4145 a_7229_43940# a_1423_45028# 0.024468f
C4146 a_9482_43914# a_14180_45002# 0.022677f
C4147 a_5807_45002# a_6165_46155# 0.039202f
C4148 a_9313_45822# a_8049_45260# 0.086184f
C4149 a_n743_46660# a_472_46348# 0.076758f
C4150 a_n881_46662# a_13925_46122# 0.019683f
C4151 a_11309_47204# a_11189_46129# 0.03753f
C4152 a_n2293_46634# a_1823_45246# 0.230429f
C4153 a_22589_40599# a_22629_38406# 0.032572f
C4154 VDAC_Pi VDD 0.591846f
C4155 a_22527_39145# a_22537_39537# 0.351623f
C4156 a_22581_37893# a_22613_38993# 0.275268f
C4157 a_7754_39964# RST_Z 0.843939f
C4158 a_10991_42826# a_10341_42308# 0.035667f
C4159 a_n443_42852# a_3626_43646# 0.027303f
C4160 a_21588_30879# a_14097_32519# 0.056136f
C4161 a_n2293_42834# a_n2661_42834# 0.202366f
C4162 a_11691_44458# a_17767_44458# 0.060949f
C4163 a_742_44458# a_949_44458# 0.185221f
C4164 a_2063_45854# a_413_45260# 0.031952f
C4165 a_584_46384# a_327_44734# 0.040089f
C4166 a_4791_45118# a_n913_45002# 0.254334f
C4167 a_16327_47482# a_20841_45814# 0.161808f
C4168 a_12741_44636# a_17715_44484# 0.029877f
C4169 a_n881_46662# a_15599_45572# 0.601034f
C4170 a_4361_42308# a_5934_30871# 0.092304f
C4171 a_7845_44172# VDD 0.11772f
C4172 a_743_42282# a_8325_42308# 0.02734f
C4173 a_11967_42832# a_20766_44850# 0.042853f
C4174 a_17517_44484# a_3422_30871# 0.073987f
C4175 a_11823_42460# a_15279_43071# 0.010476f
C4176 a_20159_44458# a_20679_44626# 0.043567f
C4177 a_20362_44736# a_20640_44752# 0.118759f
C4178 a_7640_43914# a_7845_44172# 0.021949f
C4179 a_n2661_42834# a_1115_44172# 0.011443f
C4180 a_10193_42453# a_17333_42852# 0.032471f
C4181 a_9067_47204# VDD 0.47483f
C4182 a_4915_47217# DATA[5] 0.121371f
C4183 a_9290_44172# a_11322_45546# 0.077646f
C4184 a_11387_46155# a_10193_42453# 0.050391f
C4185 a_n1613_43370# a_n2661_44458# 0.05666f
C4186 a_11189_46129# a_10490_45724# 0.03271f
C4187 a_3483_46348# a_10907_45822# 0.140023f
C4188 a_13747_46662# a_20567_45036# 0.026034f
C4189 a_19321_45002# a_18184_42460# 0.094476f
C4190 a_12741_44636# a_15861_45028# 0.075863f
C4191 a_13467_32519# EN_VIN_BSTR_N 0.03202f
C4192 a_16759_43396# VDD 0.191873f
C4193 a_n2293_43922# a_10341_43396# 0.022718f
C4194 a_20623_43914# a_15493_43940# 0.040969f
C4195 a_2711_45572# a_16147_45260# 0.028186f
C4196 a_12549_44172# a_10949_43914# 0.052089f
C4197 a_n1925_42282# a_1307_43914# 0.03653f
C4198 a_n2293_46098# a_n2661_44458# 0.026753f
C4199 a_8049_45260# a_7705_45326# 0.032872f
C4200 a_10490_45724# a_11136_45572# 0.048799f
C4201 a_17339_46660# a_18248_44752# 0.019889f
C4202 a_2324_44458# a_8560_45348# 0.070986f
C4203 a_4791_45118# a_2107_46812# 0.078338f
C4204 a_4883_46098# a_9804_47204# 0.020011f
C4205 a_16327_47482# a_13661_43548# 0.132061f
C4206 a_n2109_47186# a_5385_46902# 0.013334f
C4207 a_19339_43156# VDD 0.338297f
C4208 a_2982_43646# a_2813_43396# 0.096538f
C4209 a_6031_43396# a_6765_43638# 0.053479f
C4210 a_6293_42852# a_6197_43396# 0.213423f
C4211 a_n97_42460# a_10341_43396# 0.917198f
C4212 a_n913_45002# a_13258_32519# 0.025596f
C4213 a_18184_42460# a_22765_42852# 0.012194f
C4214 a_n2472_45546# VDD 0.290266f
C4215 a_19692_46634# a_21381_43940# 0.022586f
C4216 a_n1059_45260# a_3537_45260# 0.162323f
C4217 a_13249_42308# a_11827_44484# 0.029876f
C4218 a_13259_45724# a_13213_44734# 0.020051f
C4219 a_9313_45822# a_8953_45546# 0.038855f
C4220 a_7577_46660# a_8145_46902# 0.170059f
C4221 a_4915_47217# a_13759_46122# 0.024639f
C4222 a_7411_46660# a_8667_46634# 0.043475f
C4223 a_6540_46812# a_6755_46942# 0.057503f
C4224 a_3754_38802# a_3754_38470# 0.02792f
C4225 a_22485_38105# VDD 1.31335f
C4226 a_n901_43156# a_n1076_43230# 0.234322f
C4227 a_n1853_43023# a_n1736_43218# 0.183149f
C4228 a_16137_43396# a_17333_42852# 0.01487f
C4229 a_7276_45260# VDD 0.093163f
C4230 a_413_45260# a_n2661_42834# 0.023284f
C4231 a_n2661_43370# a_n2840_44458# 0.011391f
C4232 a_19778_44110# a_18494_42460# 0.04586f
C4233 a_20205_31679# a_14401_32519# 0.054064f
C4234 a_1823_45246# a_743_42282# 0.06422f
C4235 a_22365_46825# a_12741_44636# 0.062216f
C4236 a_n2293_46634# a_n2293_45546# 0.065405f
C4237 a_n881_46662# a_5263_45724# 0.180025f
C4238 a_11415_45002# a_22591_46660# 0.172844f
C4239 a_15368_46634# a_15015_46420# 0.012546f
C4240 a_3090_45724# a_2324_44458# 0.684819f
C4241 a_14976_45028# a_14840_46494# 0.010576f
C4242 a_17517_44484# VDD 2.99662f
C4243 a_1307_43914# a_3737_43940# 0.058797f
C4244 a_584_46384# a_4223_44672# 0.044788f
C4245 a_4791_45118# a_n2661_44458# 0.095212f
C4246 a_167_45260# a_n443_42852# 0.246952f
C4247 a_5732_46660# a_3357_43084# 0.017659f
C4248 a_768_44030# a_1423_45028# 0.096238f
C4249 a_n1151_42308# a_n1177_44458# 0.021669f
C4250 a_17715_44484# a_16375_45002# 0.026655f
C4251 a_n743_46660# a_6171_45002# 0.140224f
C4252 a_12861_44030# a_11827_44484# 0.466435f
C4253 a_13661_43548# a_14537_43396# 0.505634f
C4254 a_17957_46116# a_18147_46436# 0.011458f
C4255 a_n2293_42834# a_n1423_42826# 0.011631f
C4256 a_n2293_43922# a_n97_42460# 0.136247f
C4257 a_7499_43078# a_7309_42852# 0.011818f
C4258 a_5167_46660# VDD 0.203378f
C4259 a_n2810_45572# a_n3674_37592# 0.025877f
C4260 a_8270_45546# a_5883_43914# 0.20967f
C4261 a_6755_46942# a_14539_43914# 0.094724f
C4262 a_13747_46662# a_20679_44626# 0.030878f
C4263 a_12549_44172# a_3422_30871# 0.148646f
C4264 a_167_45260# a_375_42282# 0.017297f
C4265 a_17339_46660# a_16922_45042# 0.02918f
C4266 a_16375_45002# a_15861_45028# 0.029833f
C4267 a_8199_44636# a_8953_45002# 0.12099f
C4268 a_5937_45572# a_8191_45002# 0.180306f
C4269 a_2711_45572# a_9049_44484# 0.025215f
C4270 a_n237_47217# a_n881_46662# 0.958566f
C4271 a_2905_45572# a_2747_46873# 0.010677f
C4272 a_n2497_47436# a_768_44030# 0.023758f
C4273 a_15507_47210# a_15673_47210# 0.81159f
C4274 a_11323_42473# a_5742_30871# 0.198522f
C4275 a_n3674_38680# a_n3420_39616# 0.020072f
C4276 a_6945_45028# CLK 0.027466f
C4277 a_11967_42832# a_12089_42308# 0.022254f
C4278 a_22223_46124# EN_OFFSET_CAL 0.011048f
C4279 a_21363_45546# a_21188_45572# 0.233657f
C4280 a_20841_45814# a_20731_45938# 0.097745f
C4281 a_20623_45572# a_20528_45572# 0.049827f
C4282 a_4883_46098# a_19692_46634# 0.058277f
C4283 a_n971_45724# a_n1991_46122# 0.010501f
C4284 a_5742_30871# C0_P_btm 0.014563f
C4285 a_n3420_38528# a_n3690_38304# 0.018295f
C4286 a_5891_43370# a_5934_30871# 0.027588f
C4287 a_19256_45572# VDD 0.27151f
C4288 a_17339_46660# a_15743_43084# 0.450316f
C4289 a_13259_45724# a_11341_43940# 0.045479f
C4290 a_19692_46634# a_5649_42852# 0.01341f
C4291 a_n357_42282# a_n2661_42282# 0.055806f
C4292 a_4791_45118# a_5907_45546# 0.02288f
C4293 a_n971_45724# a_7499_43078# 0.857375f
C4294 a_2107_46812# a_6945_45028# 0.028356f
C4295 a_19692_46634# a_21188_46660# 0.022017f
C4296 C0_P_btm C0_dummy_P_btm 7.97415f
C4297 a_18194_34908# VDD 2.25174f
C4298 a_4190_30871# a_21356_42826# 0.011885f
C4299 a_13720_44458# VDD 0.202097f
C4300 a_n1557_42282# a_n3674_37592# 0.022251f
C4301 a_10157_44484# a_9313_44734# 0.026406f
C4302 a_5343_44458# a_5708_44484# 0.048542f
C4303 a_n357_42282# a_16823_43084# 0.016884f
C4304 a_949_44458# a_n2661_43922# 0.055363f
C4305 a_18494_42460# a_20159_44458# 0.024732f
C4306 a_n1613_43370# a_n1059_45260# 0.202724f
C4307 a_n746_45260# a_n2661_43370# 0.060205f
C4308 a_584_46384# a_n2293_42834# 0.049322f
C4309 a_12861_44030# a_15595_45028# 0.012748f
C4310 a_8270_45546# a_8162_45546# 0.170838f
C4311 a_17364_32525# a_13258_32519# 0.053358f
C4312 a_10341_42308# a_10723_42308# 0.024028f
C4313 a_13678_32519# a_22775_42308# 0.024479f
C4314 a_5649_42852# a_21613_42308# 0.02466f
C4315 a_742_44458# a_n97_42460# 0.083982f
C4316 a_14539_43914# a_15037_43940# 0.054182f
C4317 a_n1925_42282# a_n1736_42282# 0.029727f
C4318 a_12549_44172# VDD 3.08339f
C4319 a_n881_46662# DATA[5] 0.082222f
C4320 a_768_44030# a_6109_44484# 0.04198f
C4321 a_8049_45260# a_12427_45724# 0.012343f
C4322 a_16327_47482# a_11967_42832# 0.241578f
C4323 a_n863_45724# a_n443_42852# 0.556081f
C4324 a_13059_46348# a_13556_45296# 0.274813f
C4325 a_167_45260# a_2437_43646# 0.025008f
C4326 a_584_46384# a_1115_44172# 0.174981f
C4327 a_n237_47217# a_n443_46116# 0.110841f
C4328 a_2063_45854# a_2905_45572# 0.037943f
C4329 a_n1741_47186# a_6851_47204# 0.030234f
C4330 a_5111_42852# VDD 0.178652f
C4331 a_n1794_35082# a_6123_31319# 0.036823f
C4332 a_21076_30879# VREF_GND 0.041931f
C4333 a_5111_44636# a_5193_42852# 0.018763f
C4334 a_13249_42308# a_13575_42558# 0.088907f
C4335 a_11823_42460# a_14113_42308# 0.103699f
C4336 a_1208_46090# VDD 0.178097f
C4337 a_n2293_45546# a_626_44172# 0.150062f
C4338 a_4185_45028# a_n356_44636# 1.54308f
C4339 a_2324_44458# a_4743_44484# 0.042685f
C4340 a_n863_45724# a_375_42282# 0.451905f
C4341 a_n1613_43370# a_948_46660# 0.281392f
C4342 a_13747_46662# a_19594_46812# 0.03826f
C4343 a_2747_46873# a_2443_46660# 0.129886f
C4344 a_n1151_42308# a_11813_46116# 0.019835f
C4345 a_n4064_40160# a_n4334_39392# 0.013157f
C4346 a_9803_43646# a_10149_43396# 0.013377f
C4347 a_n97_42460# a_n901_43156# 0.011039f
C4348 a_n2956_37592# a_n3565_38216# 0.074137f
C4349 a_11525_45546# VDD 0.133093f
C4350 a_n2293_43922# a_12800_43218# 0.011493f
C4351 a_9482_43914# a_13777_45326# 0.206086f
C4352 a_3483_46348# a_9801_43940# 0.027985f
C4353 a_7499_43078# a_9313_44734# 0.0624f
C4354 a_3090_45724# a_14579_43548# 0.074713f
C4355 a_n2293_46634# a_1138_42852# 0.023262f
C4356 a_12469_46902# a_12816_46660# 0.051162f
C4357 a_n743_46660# a_376_46348# 0.076781f
C4358 a_n881_46662# a_13759_46122# 0.01582f
C4359 a_11453_44696# a_6945_45028# 0.022389f
C4360 a_n3565_38216# VREF 0.057702f
C4361 CAL_N a_22629_38406# 0.204616f
C4362 a_n3420_37984# VIN_P 0.067554f
C4363 a_7754_39964# VDD 0.848281f
C4364 a_n4209_38216# VCM 0.035453f
C4365 a_22589_40055# a_22537_39537# 0.035975f
C4366 a_22527_39145# a_22889_38993# 0.010853f
C4367 a_19237_31679# a_13258_32519# 0.055803f
C4368 a_10796_42968# a_10341_42308# 0.65943f
C4369 a_10991_42826# a_10922_42852# 0.209641f
C4370 a_8953_45546# a_7871_42858# 0.017048f
C4371 a_11823_42460# a_13565_43940# 0.046344f
C4372 a_13259_45724# a_10341_43396# 0.08137f
C4373 a_11691_44458# a_16979_44734# 0.12231f
C4374 a_11827_44484# a_18287_44626# 0.024541f
C4375 a_584_46384# a_413_45260# 0.164383f
C4376 a_4791_45118# a_n1059_45260# 0.020789f
C4377 a_16327_47482# a_20273_45572# 0.050306f
C4378 a_n1151_42308# a_n967_45348# 0.170453f
C4379 a_7542_44172# VDD 0.412456f
C4380 a_16795_42852# a_16877_42852# 0.171361f
C4381 a_11967_42832# a_20835_44721# 0.033569f
C4382 a_17517_44484# a_21398_44850# 0.01617f
C4383 a_6575_47204# VDD 1.32036f
C4384 a_4915_47217# DATA[4] 0.069022f
C4385 a_11823_42460# a_5534_30871# 0.511874f
C4386 a_20159_44458# a_20640_44752# 0.042415f
C4387 a_7640_43914# a_7542_44172# 0.20977f
C4388 a_10193_42453# a_18083_42858# 0.037244f
C4389 a_16327_47482# a_18989_43940# 0.100946f
C4390 a_11133_46155# a_10193_42453# 0.039441f
C4391 a_9290_44172# a_10490_45724# 0.022805f
C4392 a_19321_45002# a_19778_44110# 0.568668f
C4393 a_12741_44636# a_8696_44636# 2.20704f
C4394 a_4190_30871# C10_P_btm 0.446355f
C4395 a_16977_43638# VDD 0.206333f
C4396 a_20365_43914# a_15493_43940# 0.048673f
C4397 a_13483_43940# a_14021_43940# 0.109097f
C4398 a_n863_45724# a_2437_43646# 0.071802f
C4399 a_526_44458# a_1307_43914# 0.467539f
C4400 a_15227_44166# a_9313_44734# 0.06548f
C4401 a_n2442_46660# a_n3674_39768# 0.023663f
C4402 a_16327_47482# a_5807_45002# 0.451783f
C4403 a_16023_47582# a_16131_47204# 0.057222f
C4404 a_4883_46098# a_8128_46384# 0.010382f
C4405 a_2063_45854# a_2443_46660# 0.017518f
C4406 a_n2109_47186# a_4817_46660# 0.028101f
C4407 a_18599_43230# VDD 0.197104f
C4408 a_18494_42460# a_20356_42852# 0.014237f
C4409 a_18184_42460# a_20753_42852# 0.029113f
C4410 a_14021_43940# a_13678_32519# 0.021333f
C4411 a_6031_43396# a_6197_43396# 0.581047f
C4412 a_n2661_45546# VDD 0.733118f
C4413 a_20202_43084# a_11341_43940# 0.033215f
C4414 a_n2017_45002# a_3537_45260# 0.033622f
C4415 a_11823_42460# a_11691_44458# 0.022559f
C4416 a_n913_45002# a_3065_45002# 0.225034f
C4417 a_9313_45822# a_5937_45572# 0.137696f
C4418 a_7411_46660# a_7927_46660# 0.105839f
C4419 a_7754_38968# a_3754_38470# 0.209356f
C4420 a_n2157_42858# a_n1736_43218# 0.089677f
C4421 a_16409_43396# a_16795_42852# 0.010927f
C4422 a_5205_44484# VDD 0.508148f
C4423 a_13259_45724# a_n97_42460# 0.182889f
C4424 a_19778_44110# a_18184_42460# 0.119002f
C4425 a_765_45546# a_167_45260# 0.276049f
C4426 a_7715_46873# a_5066_45546# 0.020181f
C4427 a_14976_45028# a_15015_46420# 0.012921f
C4428 a_17061_44734# VDD 0.17647f
C4429 a_3422_30871# EN_VIN_BSTR_N 0.182769f
C4430 a_5755_42852# a_6101_43172# 0.013377f
C4431 a_n357_42282# a_12545_42858# 0.042417f
C4432 a_n2661_43922# a_n2293_43922# 0.05908f
C4433 a_n356_44636# a_11967_42832# 0.025796f
C4434 a_n2442_46660# a_n4315_30879# 0.361271f
C4435 a_5907_46634# a_3357_43084# 0.013466f
C4436 a_1823_45246# a_1609_45822# 0.35471f
C4437 a_17957_46116# a_13259_45724# 0.011559f
C4438 a_10809_44734# a_12379_46436# 0.011204f
C4439 a_1427_43646# VDD 0.19291f
C4440 a_n4318_38680# a_n4064_38528# 0.047936f
C4441 a_n2293_42282# a_n2472_42282# 0.163758f
C4442 a_n2293_42834# a_n1991_42858# 0.02898f
C4443 a_5385_46902# VDD 0.203316f
C4444 a_1138_42852# a_626_44172# 0.010739f
C4445 a_8270_45546# a_8701_44490# 0.015888f
C4446 a_6755_46942# a_16112_44458# 0.023983f
C4447 a_19321_45002# a_20159_44458# 0.065041f
C4448 a_13747_46662# a_20640_44752# 0.027627f
C4449 a_n443_42852# a_11823_42460# 0.356965f
C4450 a_8199_44636# a_8191_45002# 0.234072f
C4451 a_16375_45002# a_8696_44636# 0.043034f
C4452 a_5937_45572# a_7705_45326# 0.070066f
C4453 a_9290_44172# a_6171_45002# 0.028032f
C4454 a_13259_45724# a_16020_45572# 0.024851f
C4455 a_19466_46812# a_19929_45028# 0.012303f
C4456 a_15507_47210# a_15811_47375# 0.170975f
C4457 a_11599_46634# a_15673_47210# 0.012504f
C4458 a_n746_45260# a_n881_46662# 0.190303f
C4459 a_n237_47217# a_n1613_43370# 0.034341f
C4460 a_2952_47436# a_2747_46873# 0.078913f
C4461 a_6151_47436# a_4883_46098# 0.032223f
C4462 a_10723_42308# a_5742_30871# 0.185564f
C4463 a_n1917_43396# a_n1809_43762# 0.057222f
C4464 a_11967_42832# a_12379_42858# 0.492977f
C4465 a_n1533_46116# VDD 0.143145f
C4466 a_n1151_42308# a_n1853_43023# 0.021207f
C4467 a_3090_45724# a_19478_44306# 0.027139f
C4468 a_20273_45572# a_20731_45938# 0.034619f
C4469 a_16327_47482# a_16867_43762# 0.012196f
C4470 a_15227_44166# a_17737_43940# 0.013191f
C4471 a_n971_45724# a_n1853_46287# 0.08556f
C4472 a_4883_46098# a_19466_46812# 0.028345f
C4473 a_11599_46634# a_16388_46812# 0.24092f
C4474 a_n237_47217# a_n2293_46098# 0.044593f
C4475 a_n4315_30879# a_n3420_37440# 0.039346f
C4476 a_8515_42308# VDD 0.194691f
C4477 a_5742_30871# C1_P_btm 0.026156f
C4478 a_n4064_40160# a_n3565_37414# 4.2965f
C4479 a_n4209_38502# a_n4064_37984# 0.028133f
C4480 a_n3565_38502# a_n3420_37984# 0.028236f
C4481 a_n4064_38528# a_n4209_38216# 0.028013f
C4482 a_n3420_38528# a_n3565_38216# 0.035254f
C4483 a_n3690_38528# a_n3690_38304# 0.052468f
C4484 a_2982_43646# a_5534_30871# 0.094381f
C4485 a_5891_43370# a_7963_42308# 0.036306f
C4486 a_19431_45546# VDD 0.342308f
C4487 a_20202_43084# a_10341_43396# 0.037863f
C4488 a_17339_46660# a_18783_43370# 0.02025f
C4489 a_3065_45002# a_n2661_44458# 0.027917f
C4490 a_4791_45118# a_5263_45724# 0.021183f
C4491 a_15227_46910# a_13059_46348# 0.043664f
C4492 C1_P_btm C0_dummy_P_btm 1.24905f
C4493 EN_VIN_BSTR_N VDD 1.19259f
C4494 a_13076_44458# VDD 0.180665f
C4495 a_3080_42308# a_n1794_35082# 0.032975f
C4496 a_9838_44484# a_9313_44734# 0.037628f
C4497 a_20692_30879# a_13678_32519# 0.051702f
C4498 a_3232_43370# a_11750_44172# 0.020452f
C4499 a_742_44458# a_n2661_43922# 0.066714f
C4500 a_18184_42460# a_20159_44458# 0.01449f
C4501 a_13507_46334# a_22775_42308# 0.022177f
C4502 SMPL_ON_N a_13258_32519# 0.030848f
C4503 a_4883_46098# a_5111_44636# 0.048482f
C4504 a_10227_46804# a_8953_45002# 0.017713f
C4505 a_11415_45002# a_13259_45724# 0.505354f
C4506 a_n1613_43370# a_n2017_45002# 0.015448f
C4507 a_n971_45724# a_n2661_43370# 0.064346f
C4508 a_768_44030# a_3357_43084# 0.09747f
C4509 a_15227_44166# a_2711_45572# 0.113396f
C4510 a_18189_46348# a_17957_46116# 0.038851f
C4511 a_10341_42308# a_10533_42308# 0.035479f
C4512 a_5649_42852# a_21887_42336# 0.017243f
C4513 a_13678_32519# a_21613_42308# 0.024855f
C4514 a_12891_46348# VDD 1.01428f
C4515 a_n881_46662# DATA[4] 0.087677f
C4516 a_8199_44636# a_8685_42308# 0.114007f
C4517 a_5111_44636# a_5649_42852# 0.121004f
C4518 a_2957_45546# a_3218_45724# 0.063846f
C4519 a_8049_45260# a_11962_45724# 0.019556f
C4520 a_n2293_45546# a_1609_45822# 0.159696f
C4521 a_2202_46116# a_2437_43646# 0.022869f
C4522 a_12861_44030# a_19279_43940# 0.152657f
C4523 a_16327_47482# a_19006_44850# 0.028858f
C4524 a_13059_46348# a_9482_43914# 0.448068f
C4525 a_10586_45546# a_10193_42453# 0.380236f
C4526 a_n755_45592# a_n356_45724# 0.016853f
C4527 a_n746_45260# a_n443_46116# 0.060788f
C4528 a_n971_45724# a_4915_47217# 0.017974f
C4529 a_1431_47204# a_n1151_42308# 0.013895f
C4530 a_n237_47217# a_4791_45118# 0.10712f
C4531 a_n1741_47186# a_6491_46660# 0.023524f
C4532 a_4520_42826# VDD 0.142755f
C4533 a_n913_45002# a_14635_42282# 0.332583f
C4534 a_21076_30879# VREF 0.417978f
C4535 a_13249_42308# a_13070_42354# 0.141799f
C4536 a_805_46414# VDD 0.154663f
C4537 a_10227_46804# a_3626_43646# 0.011826f
C4538 a_2324_44458# a_n699_43396# 0.070009f
C4539 a_n2661_45546# a_1423_45028# 0.020024f
C4540 a_n1613_43370# a_1123_46634# 0.358475f
C4541 a_13747_46662# a_19321_45002# 0.080725f
C4542 a_768_44030# a_n2293_46634# 0.26984f
C4543 a_n1151_42308# a_11735_46660# 0.050593f
C4544 a_16877_42852# VDD 0.192454f
C4545 a_n4064_40160# a_n4209_39304# 0.04848f
C4546 a_n784_42308# EN_VIN_BSTR_N 0.051272f
C4547 a_n2946_39866# a_n4064_39616# 0.053228f
C4548 a_n1794_35082# a_n1057_35014# 0.017188f
C4549 a_n4315_30879# a_n3565_39304# 0.048127f
C4550 a_14955_43396# a_10341_43396# 0.01411f
C4551 a_2982_43646# a_4190_30871# 0.3223f
C4552 a_11322_45546# VDD 0.370908f
C4553 a_n2810_45028# a_n3565_38216# 0.349341f
C4554 a_9482_43914# a_13556_45296# 0.726155f
C4555 a_n967_45348# a_n2293_42834# 0.038042f
C4556 a_n2293_45010# a_n2661_43370# 0.067876f
C4557 a_5205_44484# a_1423_45028# 0.821456f
C4558 a_11901_46660# a_12816_46660# 0.125324f
C4559 a_n2497_47436# a_n2661_45546# 0.030609f
C4560 CAL_N CAL_P 5.92093f
C4561 a_22527_39145# a_22613_38993# 0.12129f
C4562 a_22589_40055# a_22889_38993# 0.19183f
C4563 a_7754_40130# RST_Z 0.022036f
C4564 a_10796_42968# a_10922_42852# 0.170059f
C4565 a_10835_43094# a_10341_42308# 0.541777f
C4566 a_n2661_44458# a_6298_44484# 0.025865f
C4567 a_n443_42852# a_2982_43646# 0.037773f
C4568 a_11691_44458# a_14539_43914# 0.268287f
C4569 a_11415_45002# a_18189_46348# 0.028334f
C4570 a_4791_45118# a_n2017_45002# 0.023951f
C4571 a_n2661_46634# a_11823_42460# 0.331717f
C4572 a_16327_47482# a_20107_45572# 0.674639f
C4573 a_9313_45822# a_2437_43646# 0.045826f
C4574 a_n743_46660# a_10193_42453# 0.25279f
C4575 a_7281_43914# VDD 0.198809f
C4576 a_4361_42308# a_6123_31319# 0.065399f
C4577 a_13249_42308# a_12545_42858# 0.030353f
C4578 a_11967_42832# a_20679_44626# 0.863531f
C4579 a_17517_44484# a_20980_44850# 0.026284f
C4580 a_7903_47542# VDD 0.202868f
C4581 a_11823_42460# a_14543_43071# 0.028488f
C4582 a_4915_47217# DATA[3] 0.07179f
C4583 a_20159_44458# a_20362_44736# 0.233657f
C4584 a_n2661_42834# a_175_44278# 0.010875f
C4585 a_5111_44636# a_8685_43396# 0.078598f
C4586 a_1307_43914# a_3626_43646# 0.012223f
C4587 a_16327_47482# a_18374_44850# 0.16003f
C4588 a_13661_43548# a_18494_42460# 0.049953f
C4589 a_13747_46662# a_18184_42460# 0.123281f
C4590 a_19321_45002# a_18911_45144# 0.050257f
C4591 a_10355_46116# a_10490_45724# 0.01084f
C4592 a_11189_46129# a_10193_42453# 0.123385f
C4593 a_16409_43396# VDD 0.250832f
C4594 a_20269_44172# a_15493_43940# 0.051355f
C4595 a_20935_43940# a_21115_43940# 0.185422f
C4596 a_13483_43940# a_13829_44260# 0.013377f
C4597 a_12359_47026# VDD 0.142103f
C4598 a_n2442_46660# a_n4318_39768# 0.023739f
C4599 a_13507_46334# a_14021_43940# 0.01995f
C4600 a_8049_45260# a_7229_43940# 0.014199f
C4601 a_16327_47482# a_16131_47204# 0.016621f
C4602 a_9313_45822# a_n2661_46634# 0.032598f
C4603 a_13717_47436# a_21588_30879# 0.052863f
C4604 a_11599_46634# a_19321_45002# 0.091019f
C4605 a_2063_45854# a_n2661_46098# 0.021195f
C4606 a_n356_44636# a_n2293_42282# 1.10197f
C4607 a_14021_43940# a_21855_43396# 0.025748f
C4608 a_6031_43396# a_6293_42852# 0.163953f
C4609 a_n913_45002# a_19511_42282# 0.120073f
C4610 a_n2810_45572# VDD 0.557886f
C4611 a_n755_45592# a_n356_44636# 2.42652f
C4612 a_12549_44172# a_20556_43646# 0.125209f
C4613 a_n1059_45260# a_3065_45002# 0.023485f
C4614 a_9313_45822# a_8199_44636# 0.015956f
C4615 a_7715_46873# a_7577_46660# 0.205227f
C4616 a_n237_47217# a_6945_45028# 0.072758f
C4617 a_n1151_42308# a_2324_44458# 0.075066f
C4618 a_7411_46660# a_8145_46902# 0.053385f
C4619 a_5807_45002# a_16721_46634# 0.112018f
C4620 a_13747_46662# a_13059_46348# 0.273684f
C4621 a_3754_38802# VDAC_Ni 0.301032f
C4622 a_n1423_42826# a_n1076_43230# 0.051162f
C4623 a_16137_43396# a_17701_42308# 0.025497f
C4624 a_16547_43609# a_16795_42852# 0.081093f
C4625 a_3422_30871# a_5934_30871# 0.02193f
C4626 a_6431_45366# VDD 0.203167f
C4627 a_n467_45028# a_n2661_43922# 0.024697f
C4628 a_10193_42453# a_11750_44172# 0.01114f
C4629 a_16922_45042# a_11827_44484# 0.032223f
C4630 a_5205_44484# a_6109_44484# 0.029986f
C4631 a_3232_43370# a_5891_43370# 0.137859f
C4632 a_3090_45724# a_15015_46420# 0.019425f
C4633 a_768_44030# a_2277_45546# 0.027945f
C4634 a_n2442_46660# a_n2956_38216# 0.048086f
C4635 a_20202_43084# a_11415_45002# 0.041726f
C4636 a_22365_46825# a_22591_46660# 0.08571f
C4637 a_n2312_38680# a_n2810_45572# 0.062154f
C4638 a_16241_44734# VDD 0.189894f
C4639 a_3422_30871# a_10890_34112# 0.19148f
C4640 a_n357_42282# a_12089_42308# 0.027195f
C4641 a_n2661_42834# a_n2293_43922# 0.034793f
C4642 a_n443_42852# a_7871_42858# 0.013386f
C4643 a_10193_42453# a_4361_42308# 0.274131f
C4644 a_n699_43396# a_n1761_44111# 0.018554f
C4645 a_11599_46634# a_18184_42460# 0.018223f
C4646 a_768_44030# a_626_44172# 0.186913f
C4647 a_584_46384# a_949_44458# 0.011926f
C4648 a_1823_45246# a_n443_42852# 0.125287f
C4649 a_n971_45724# a_5883_43914# 0.027317f
C4650 a_18189_46348# a_13259_45724# 0.016675f
C4651 a_n1557_42282# VDD 0.355513f
C4652 a_4817_46660# VDD 0.370615f
C4653 a_n2293_42834# a_n1853_43023# 0.053782f
C4654 a_19321_45002# a_19615_44636# 0.035767f
C4655 a_8016_46348# a_8953_45002# 0.016464f
C4656 a_5937_45572# a_6709_45028# 0.629301f
C4657 a_2711_45572# a_8568_45546# 0.011004f
C4658 a_3483_46348# a_14537_43396# 0.087339f
C4659 a_9290_44172# a_3232_43370# 0.087744f
C4660 a_13259_45724# a_17478_45572# 0.048668f
C4661 a_11599_46634# a_15811_47375# 0.107881f
C4662 a_n1741_47186# a_9804_47204# 0.010096f
C4663 a_n971_45724# a_n881_46662# 0.236696f
C4664 a_n746_45260# a_n1613_43370# 0.146842f
C4665 a_2553_47502# a_2747_46873# 0.14563f
C4666 a_4915_47217# a_12465_44636# 0.07724f
C4667 a_10533_42308# a_5742_30871# 0.020913f
C4668 a_n4318_37592# a_n4064_40160# 0.079413f
C4669 a_n1917_43396# a_n2012_43396# 0.049827f
C4670 a_n1699_43638# a_n1809_43762# 0.097745f
C4671 a_n913_45002# a_4921_42308# 0.169235f
C4672 a_6945_45028# DATA[5] 0.047689f
C4673 a_2711_45572# a_n2661_43370# 0.112998f
C4674 a_3090_45724# a_15493_43396# 0.134629f
C4675 a_20273_45572# a_20528_45572# 0.064178f
C4676 a_20841_45814# a_21188_45572# 0.051162f
C4677 a_15227_44166# a_15682_43940# 0.072383f
C4678 a_9313_45822# a_765_45546# 0.034184f
C4679 a_11599_46634# a_13059_46348# 0.371555f
C4680 a_n743_46660# a_4646_46812# 0.031686f
C4681 a_n746_45260# a_n2293_46098# 0.027821f
C4682 a_13507_46334# a_19692_46634# 0.823157f
C4683 a_768_44030# a_6755_46942# 0.017611f
C4684 a_n1925_46634# a_4955_46873# 0.033508f
C4685 a_5934_30871# VDD 0.431179f
C4686 a_5742_30871# C2_P_btm 0.030783f
C4687 a_n3420_38528# a_n4334_38304# 0.014479f
C4688 a_1666_39043# a_2113_38308# 0.088649f
C4689 a_16137_43396# a_4361_42308# 0.019831f
C4690 a_5891_43370# a_6123_31319# 0.028865f
C4691 a_3905_42865# a_4649_42852# 0.04156f
C4692 a_18691_45572# VDD 0.191893f
C4693 a_17339_46660# a_18525_43370# 0.060382f
C4694 a_19692_46634# a_21855_43396# 0.016876f
C4695 a_n467_45028# a_n452_44636# 0.092885f
C4696 a_768_44030# a_8049_45260# 0.027975f
C4697 a_n971_45724# a_8162_45546# 0.015463f
C4698 a_19692_46634# a_20623_46660# 0.03624f
C4699 a_4915_47217# a_2711_45572# 0.265557f
C4700 a_15227_44166# a_22000_46634# 0.154332f
C4701 a_5257_43370# a_5164_46348# 0.02844f
C4702 a_16327_47482# a_n357_42282# 0.49929f
C4703 C2_P_btm C0_dummy_P_btm 7.14548f
C4704 C1_P_btm C0_P_btm 11.2332f
C4705 a_10890_34112# VDD 0.345626f
C4706 a_n1557_42282# a_n784_42308# 0.058812f
C4707 a_12883_44458# VDD 0.263743f
C4708 a_18494_42460# a_11967_42832# 0.025796f
C4709 a_5883_43914# a_9313_44734# 0.124999f
C4710 a_20205_31679# a_13678_32519# 0.051502f
C4711 a_8975_43940# a_5891_43370# 0.021307f
C4712 a_742_44458# a_n2661_42834# 0.034578f
C4713 a_13507_46334# a_21613_42308# 0.035917f
C4714 a_12594_46348# a_10809_44734# 0.082565f
C4715 a_14209_32519# a_13258_32519# 0.051594f
C4716 a_10835_43094# a_5742_30871# 0.011953f
C4717 a_13678_32519# a_21887_42336# 0.012293f
C4718 a_4185_45028# a_5742_30871# 0.062132f
C4719 a_11309_47204# VDD 0.358104f
C4720 a_n1925_42282# a_n2104_42282# 0.166917f
C4721 a_n2956_37592# a_n4318_38680# 0.023187f
C4722 a_n809_44244# a_n984_44318# 0.234322f
C4723 a_18597_46090# a_17517_44484# 0.021693f
C4724 a_310_45028# a_n23_45546# 0.022295f
C4725 a_n2293_45546# a_n443_42852# 0.084694f
C4726 a_1823_45246# a_2437_43646# 0.324477f
C4727 a_16327_47482# a_18588_44850# 0.012252f
C4728 a_13059_46348# a_13348_45260# 0.010157f
C4729 a_n1151_42308# a_n1761_44111# 0.642214f
C4730 a_n755_45592# a_3503_45724# 0.163919f
C4731 a_2063_45854# a_2553_47502# 0.040297f
C4732 a_n971_45724# a_n443_46116# 0.129009f
C4733 a_n1741_47186# a_6545_47178# 0.053219f
C4734 a_3935_42891# VDD 0.096403f
C4735 a_n784_42308# a_5934_30871# 0.142087f
C4736 a_18579_44172# a_18525_43370# 0.012789f
C4737 a_472_46348# VDD 0.706547f
C4738 a_n913_45002# a_13291_42460# 0.070562f
C4739 a_n1059_45260# a_14635_42282# 0.063373f
C4740 a_n2956_38216# a_n3565_39304# 0.02162f
C4741 a_21076_30879# VIN_N 0.067776f
C4742 a_20820_30879# VCM 0.05604f
C4743 a_n863_45724# a_1307_43914# 0.050349f
C4744 a_n2293_45546# a_375_42282# 0.104283f
C4745 a_9290_44172# a_8975_43940# 0.114958f
C4746 a_2324_44458# a_4223_44672# 0.56408f
C4747 a_n1613_43370# a_383_46660# 0.182504f
C4748 a_6151_47436# a_8035_47026# 0.038687f
C4749 a_9804_47204# a_n743_46660# 0.295465f
C4750 a_16245_42852# VDD 0.205729f
C4751 a_n3420_39616# a_n4064_39616# 6.66063f
C4752 a_n1794_35082# a_n1696_34930# 0.46221f
C4753 a_15095_43370# a_10341_43396# 0.013375f
C4754 a_10490_45724# VDD 0.162001f
C4755 a_n2956_37592# a_n4209_38216# 0.104159f
C4756 a_2982_43646# a_21259_43561# 0.034927f
C4757 a_13348_45260# a_13556_45296# 0.189446f
C4758 en_comp a_n2293_42834# 0.103485f
C4759 a_n2472_45002# a_n2661_43370# 0.017331f
C4760 a_13017_45260# a_14180_45002# 0.079928f
C4761 a_2324_44458# a_15493_43940# 0.061147f
C4762 a_n1925_42282# a_n2661_42282# 2.27741f
C4763 a_768_44030# a_8953_45546# 0.025581f
C4764 a_12469_46902# a_12251_46660# 0.209641f
C4765 a_11901_46660# a_12991_46634# 0.042415f
C4766 a_12465_44636# a_10809_44734# 0.099854f
C4767 a_n4209_38216# VREF 0.055795f
C4768 a_11206_38545# CAL_P 0.234643f
C4769 a_n3565_38216# VIN_P 0.028666f
C4770 a_7754_40130# VDD 13.6809f
C4771 a_22537_40625# a_22537_39537# 0.604835f
C4772 a_22527_39145# a_22581_37893# 0.076507f
C4773 a_10796_42968# a_10991_42826# 0.206455f
C4774 a_10835_43094# a_10922_42852# 0.053385f
C4775 a_17730_32519# a_13258_32519# 0.05785f
C4776 a_n467_45028# a_n809_44244# 0.010788f
C4777 a_n2661_44458# a_5518_44484# 0.01193f
C4778 a_n2661_45546# a_3457_43396# 0.030099f
C4779 a_11691_44458# a_16112_44458# 0.012386f
C4780 a_11827_44484# a_17970_44736# 0.012326f
C4781 a_11415_45002# a_17715_44484# 0.032854f
C4782 a_n971_45724# a_3537_45260# 0.266743f
C4783 a_4419_46090# a_4704_46090# 0.016592f
C4784 a_n881_46662# a_15037_45618# 0.044816f
C4785 a_12741_44636# a_2324_44458# 0.019655f
C4786 a_6453_43914# VDD 0.194953f
C4787 a_4361_42308# a_7227_42308# 0.01047f
C4788 a_18249_42858# a_18504_43218# 0.05936f
C4789 a_16414_43172# a_16245_42852# 0.08213f
C4790 a_n2661_43922# a_n809_44244# 0.010689f
C4791 a_n2661_42834# a_n984_44318# 0.012148f
C4792 a_11967_42832# a_20640_44752# 0.588649f
C4793 a_7227_47204# VDD 0.430714f
C4794 a_10809_44734# a_2711_45572# 0.037787f
C4795 a_2063_45854# a_n2661_43922# 0.033229f
C4796 a_11415_45002# a_15861_45028# 0.041647f
C4797 a_16327_47482# a_18443_44721# 0.1665f
C4798 a_10903_43370# a_7499_43078# 0.888628f
C4799 a_13747_46662# a_19778_44110# 0.670692f
C4800 a_13661_43548# a_18184_42460# 0.031622f
C4801 a_3483_46348# a_8697_45822# 0.033264f
C4802 a_9290_44172# a_10193_42453# 1.23123f
C4803 a_16547_43609# VDD 0.31275f
C4804 a_19862_44208# a_15493_43940# 0.534481f
C4805 a_12156_46660# VDD 0.082428f
C4806 a_20365_43914# a_11341_43940# 0.010232f
C4807 a_n2661_45546# a_3357_43084# 0.045914f
C4808 a_768_44030# a_9028_43914# 0.113848f
C4809 a_584_46384# a_n97_42460# 0.526796f
C4810 a_2324_44458# a_n2293_42834# 0.168086f
C4811 a_n2293_45546# a_2437_43646# 0.031092f
C4812 a_16241_47178# a_16131_47204# 0.097745f
C4813 a_n2109_47186# a_4651_46660# 0.025236f
C4814 a_15673_47210# a_5807_45002# 0.011029f
C4815 a_12465_44636# a_n881_46662# 0.813228f
C4816 a_18597_46090# a_12549_44172# 0.042681f
C4817 a_584_46384# a_n2661_46098# 0.17431f
C4818 a_18184_42460# a_20256_42852# 0.01674f
C4819 a_n2840_45546# VDD 0.302566f
C4820 a_3357_43084# a_5205_44484# 0.020505f
C4821 a_12549_44172# a_743_42282# 0.119701f
C4822 a_n357_42282# a_n356_44636# 0.308599f
C4823 a_n2312_39304# a_n4318_38680# 0.0235f
C4824 a_n2017_45002# a_3065_45002# 0.043491f
C4825 a_n913_45002# a_2382_45260# 0.021705f
C4826 SMPL_ON_P a_n2956_38680# 0.039338f
C4827 a_7411_46660# a_7577_46660# 0.634781f
C4828 a_13661_43548# a_13059_46348# 0.267127f
C4829 a_5807_45002# a_16388_46812# 0.235518f
C4830 a_n2472_42826# a_n4318_38680# 0.158196f
C4831 a_n1991_42858# a_n1076_43230# 0.123255f
C4832 a_n1853_43023# a_n13_43084# 0.109925f
C4833 a_16547_43609# a_16414_43172# 0.143695f
C4834 a_6171_45002# VDD 0.441339f
C4835 a_3232_43370# a_8375_44464# 0.022129f
C4836 a_10193_42453# a_10807_43548# 0.060211f
C4837 a_n2293_46634# a_n2661_45546# 0.85166f
C4838 a_15009_46634# a_15015_46420# 0.012232f
C4839 a_5257_43370# a_5066_45546# 0.053231f
C4840 a_10227_46804# a_11823_42460# 0.428745f
C4841 a_n881_46662# a_2711_45572# 0.170524f
C4842 a_14673_44172# VDD 0.381917f
C4843 a_17538_32519# a_13258_32519# 0.054578f
C4844 a_1307_43914# a_2455_43940# 0.047238f
C4845 a_n357_42282# a_12379_42858# 0.031137f
C4846 a_n2661_42834# a_n2661_43922# 0.841361f
C4847 w_10694_33990# a_18194_34908# 0.799261f
C4848 SMPL_ON_P a_n1550_35448# 0.012033f
C4849 a_1138_42852# a_n443_42852# 0.14758f
C4850 a_1176_45822# a_1609_45822# 0.010535f
C4851 a_15368_46634# a_15599_45572# 0.100853f
C4852 a_13661_43548# a_13556_45296# 0.559682f
C4853 a_3090_45724# a_15765_45572# 0.046838f
C4854 a_584_46384# a_742_44458# 0.031608f
C4855 a_17715_44484# a_13259_45724# 0.391904f
C4856 a_4955_46873# VDD 0.467566f
C4857 a_n2293_42834# a_n2157_42858# 0.058852f
C4858 a_13259_45724# a_15861_45028# 0.16873f
C4859 a_4646_46812# a_5891_43370# 0.089437f
C4860 a_19321_45002# a_11967_42832# 0.266816f
C4861 a_2324_44458# a_413_45260# 0.021366f
C4862 a_5937_45572# a_7229_43940# 0.126047f
C4863 a_2711_45572# a_8162_45546# 0.019489f
C4864 a_n971_45724# a_n1613_43370# 0.6298f
C4865 a_2063_45854# a_2747_46873# 0.023413f
C4866 a_12861_44030# a_16327_47482# 0.120085f
C4867 a_11599_46634# a_15507_47210# 0.267808f
C4868 a_n2267_43396# a_n1809_43762# 0.034619f
C4869 a_6945_45028# DATA[4] 0.0111f
C4870 a_3090_45724# a_19328_44172# 0.153704f
C4871 a_20107_45572# a_20528_45572# 0.086377f
C4872 a_20273_45572# a_21188_45572# 0.125324f
C4873 a_15227_44166# a_14955_43940# 0.134177f
C4874 a_13249_42308# a_14537_43396# 0.020089f
C4875 a_11823_42460# a_1307_43914# 0.049611f
C4876 a_11453_44696# a_14976_45028# 0.014048f
C4877 a_n743_46660# a_3877_44458# 0.034265f
C4878 a_n2661_46634# a_5732_46660# 0.010632f
C4879 a_n971_45724# a_n2293_46098# 0.110318f
C4880 a_13507_46334# a_19466_46812# 0.03247f
C4881 a_4883_46098# a_15227_44166# 0.176028f
C4882 a_n1925_46634# a_4651_46660# 0.046762f
C4883 a_12549_44172# a_6755_46942# 0.553062f
C4884 a_n4315_30879# a_n3565_37414# 0.037486f
C4885 a_n3565_38502# a_n3565_38216# 0.0433f
C4886 a_n3420_38528# a_n4209_38216# 0.050044f
C4887 a_n4209_38502# a_n3420_37984# 0.028231f
C4888 a_n4064_40160# a_n4209_37414# 0.055461f
C4889 a_7963_42308# VDD 0.266057f
C4890 a_5742_30871# C3_P_btm 0.030866f
C4891 a_19721_31679# a_13258_32519# 0.054727f
C4892 a_15743_43084# a_16823_43084# 0.031733f
C4893 a_3499_42826# a_n2293_42282# 0.058548f
C4894 a_18909_45814# VDD 0.205795f
C4895 a_n913_45002# a_5343_44458# 0.020508f
C4896 a_17339_46660# a_18429_43548# 0.033468f
C4897 a_2382_45260# a_n2661_44458# 0.032484f
C4898 a_12549_44172# a_8049_45260# 0.031115f
C4899 a_n1151_42308# a_6511_45714# 0.044048f
C4900 a_5807_45002# a_5066_45546# 0.027744f
C4901 a_19692_46634# a_20841_46902# 0.025536f
C4902 a_n443_46116# a_2711_45572# 0.060543f
C4903 a_13507_46334# a_20205_31679# 0.023531f
C4904 C3_P_btm C0_dummy_P_btm 0.087354f
C4905 EN_VIN_BSTR_N C10_N_btm 0.320569f
C4906 C2_P_btm C0_P_btm 0.827449f
C4907 a_n217_35014# VDD 0.296751f
C4908 a_n1557_42282# a_196_42282# 0.031105f
C4909 a_12607_44458# VDD 0.188171f
C4910 a_19778_44110# a_19615_44636# 0.012379f
C4911 a_18184_42460# a_11967_42832# 0.024012f
C4912 a_5883_43914# a_9241_44734# 0.010354f
C4913 a_7499_43078# a_8685_43396# 0.153217f
C4914 a_n2293_42834# a_n1761_44111# 0.03111f
C4915 a_10057_43914# a_5891_43370# 0.197199f
C4916 a_3232_43370# a_10949_43914# 0.093316f
C4917 a_16922_45042# a_19279_43940# 0.018289f
C4918 a_20193_45348# a_17517_44484# 0.015762f
C4919 a_12861_44030# a_14537_43396# 0.015677f
C4920 a_n1613_43370# a_n2293_45010# 0.077436f
C4921 a_12005_46116# a_10809_44734# 0.029593f
C4922 a_17715_44484# a_18189_46348# 0.014348f
C4923 a_17583_46090# a_17957_46116# 0.092344f
C4924 a_5649_42852# a_7174_31319# 0.025928f
C4925 a_13467_32519# a_22775_42308# 0.016923f
C4926 a_n967_45348# a_n1076_43230# 0.019022f
C4927 a_n2956_37592# a_n3674_39304# 0.023366f
C4928 a_n2810_45028# a_n4318_38680# 0.023185f
C4929 a_n699_43396# a_n2129_43609# 0.062898f
C4930 a_n755_45592# a_133_42852# 0.020885f
C4931 a_n1099_45572# a_n23_45546# 0.042611f
C4932 a_310_45028# a_n356_45724# 0.12349f
C4933 a_17715_44484# a_17478_45572# 0.017416f
C4934 a_10586_45546# a_10053_45546# 0.024917f
C4935 a_n755_45592# a_3316_45546# 0.045656f
C4936 a_n971_45724# a_4791_45118# 0.025426f
C4937 a_1209_47178# a_n1151_42308# 0.024897f
C4938 a_584_46384# a_2553_47502# 0.100103f
C4939 a_n1741_47186# a_6151_47436# 0.071065f
C4940 a_3681_42891# VDD 0.223661f
C4941 a_5342_30871# EN_VIN_BSTR_N 0.010795f
C4942 a_3537_45260# a_5837_42852# 0.042825f
C4943 a_2711_45572# a_20107_42308# 0.164316f
C4944 a_376_46348# VDD 0.116284f
C4945 a_n1059_45260# a_13291_42460# 0.03043f
C4946 a_n2017_45002# a_14635_42282# 0.025779f
C4947 a_n913_45002# a_13003_42852# 0.026478f
C4948 a_20820_30879# VREF_GND 0.02097f
C4949 a_9290_44172# a_10057_43914# 0.034053f
C4950 a_2324_44458# a_2779_44458# 0.092751f
C4951 a_15861_45028# a_17478_45572# 0.080824f
C4952 a_n1613_43370# a_601_46902# 0.178721f
C4953 a_5807_45002# a_19321_45002# 0.376188f
C4954 a_6151_47436# a_7832_46660# 0.016469f
C4955 a_n3420_39616# a_n2946_39866# 0.236674f
C4956 a_n4315_30879# a_n4209_39304# 0.032541f
C4957 a_n1794_35082# a_n1550_35448# 0.019052f
C4958 a_n3565_39590# a_n2302_39866# 0.044102f
C4959 a_n3690_39616# a_n4064_39616# 0.085414f
C4960 a_14205_43396# a_10341_43396# 0.033299f
C4961 a_8746_45002# VDD 0.970181f
C4962 a_n2810_45028# a_n4209_38216# 0.063751f
C4963 a_13348_45260# a_9482_43914# 0.352976f
C4964 a_13017_45260# a_13777_45326# 0.195607f
C4965 a_15227_44166# a_8685_43396# 0.013522f
C4966 a_20107_45572# a_18494_42460# 0.010062f
C4967 a_526_44458# a_n2661_42282# 0.191497f
C4968 a_n2661_45010# a_n2661_43370# 0.077441f
C4969 a_768_44030# a_5937_45572# 0.05116f
C4970 a_11901_46660# a_12251_46660# 0.219633f
C4971 a_11735_46660# a_12816_46660# 0.102325f
C4972 a_22589_40599# a_22537_39537# 0.380009f
C4973 a_22589_40055# a_22581_37893# 0.461959f
C4974 a_10835_43094# a_10991_42826# 0.105839f
C4975 a_10518_42984# a_10922_42852# 0.051162f
C4976 a_11827_44484# a_17767_44458# 0.014019f
C4977 a_11691_44458# a_15004_44636# 0.221929f
C4978 a_3483_46348# a_5164_46348# 0.025074f
C4979 a_22000_46634# a_10809_44734# 0.012475f
C4980 a_n2109_47186# a_5691_45260# 0.113268f
C4981 a_18597_46090# a_19431_45546# 0.062716f
C4982 a_n2661_46634# a_11962_45724# 0.020358f
C4983 a_n971_45724# a_3429_45260# 0.171338f
C4984 a_15567_42826# a_16245_42852# 0.03084f
C4985 a_5663_43940# VDD 0.133666f
C4986 a_4361_42308# a_6761_42308# 0.042179f
C4987 a_17333_42852# a_18504_43218# 0.157683f
C4988 a_5649_42852# a_5932_42308# 0.126438f
C4989 a_10057_43914# a_10807_43548# 0.039192f
C4990 a_6109_44484# a_6453_43914# 0.165572f
C4991 a_n2661_42834# a_n809_44244# 0.021917f
C4992 a_1307_43914# a_2982_43646# 0.028987f
C4993 a_13249_42308# a_12379_42858# 0.029761f
C4994 a_11967_42832# a_20362_44736# 0.052989f
C4995 a_11823_42460# a_13635_43156# 0.040348f
C4996 a_n2293_42834# a_n2267_43396# 0.010565f
C4997 a_6851_47204# VDD 0.287724f
C4998 a_2063_45854# a_n2661_42834# 0.022984f
C4999 a_584_46384# a_n2661_43922# 0.0255f
C5000 a_11415_45002# a_8696_44636# 0.10924f
C5001 a_16327_47482# a_18287_44626# 0.552724f
C5002 a_768_44030# a_11691_44458# 0.029945f
C5003 a_12549_44172# a_20193_45348# 0.587618f
C5004 a_10227_46804# a_14539_43914# 0.012909f
C5005 a_3090_45724# a_n913_45002# 0.039732f
C5006 a_9290_44172# a_10180_45724# 0.037823f
C5007 a_10355_46116# a_10193_42453# 0.058019f
C5008 a_16243_43396# VDD 0.39865f
C5009 a_19478_44306# a_15493_43940# 0.025498f
C5010 a_13259_45724# a_17303_42282# 0.460497f
C5011 a_20623_43914# a_20935_43940# 0.040559f
C5012 a_n2956_39768# a_n3674_39768# 0.023472f
C5013 a_n1151_42308# a_n2129_43609# 0.019226f
C5014 a_20692_30879# a_20447_31679# 9.02991f
C5015 a_n2109_47186# a_4646_46812# 0.021783f
C5016 a_15673_47210# a_16131_47204# 0.034619f
C5017 a_11599_46634# a_13747_46662# 0.25325f
C5018 a_6151_47436# a_n743_46660# 0.03019f
C5019 a_584_46384# a_1799_45572# 0.179456f
C5020 a_14021_43940# a_13467_32519# 0.016437f
C5021 a_n2312_40392# a_n4318_38680# 0.025333f
C5022 a_n2312_39304# a_n3674_39304# 0.023737f
C5023 a_n1059_45260# a_2382_45260# 0.025598f
C5024 SMPL_ON_P a_n2956_39304# 0.039212f
C5025 a_9313_45822# a_8016_46348# 0.02464f
C5026 a_n971_45724# a_6945_45028# 0.247957f
C5027 a_7411_46660# a_7715_46873# 0.162909f
C5028 a_5807_45002# a_13059_46348# 0.1145f
C5029 a_7754_38968# a_7754_38636# 0.296258f
C5030 a_n4064_39072# EN_VIN_BSTR_P 1.00237f
C5031 a_n2840_42826# a_n4318_38680# 0.044261f
C5032 a_n3674_39768# a_n4318_37592# 0.023075f
C5033 a_n1423_42826# a_n1641_43230# 0.209641f
C5034 a_n1991_42858# a_n901_43156# 0.041762f
C5035 a_n1853_43023# a_n1076_43230# 0.040291f
C5036 a_16137_43396# a_16795_42852# 0.010001f
C5037 a_3232_43370# VDD 2.96597f
C5038 a_3422_30871# a_6123_31319# 0.021957f
C5039 a_15227_44166# a_17333_42852# 0.043277f
C5040 a_1307_43914# a_14539_43914# 0.131617f
C5041 a_10193_42453# a_10949_43914# 0.032349f
C5042 a_5205_44484# a_5289_44734# 0.011388f
C5043 a_22365_46825# a_20202_43084# 0.115624f
C5044 a_n1613_43370# a_2711_45572# 0.028041f
C5045 a_765_45546# a_1138_42852# 0.02041f
C5046 a_n97_42460# a_4958_30871# 0.069553f
C5047 a_3422_30871# EN_VIN_BSTR_P 0.182769f
C5048 a_5111_42852# a_5457_43172# 0.013377f
C5049 a_1307_43914# a_2253_43940# 0.056967f
C5050 a_n357_42282# a_10341_42308# 0.057131f
C5051 w_10694_33990# EN_VIN_BSTR_N 3.97924f
C5052 SMPL_ON_P a_n2002_35448# 0.399437f
C5053 a_n2956_39768# a_n4315_30879# 0.056491f
C5054 a_17583_46090# a_13259_45724# 0.191869f
C5055 a_n2293_46098# a_2711_45572# 0.530463f
C5056 a_1176_45822# a_n443_42852# 0.071187f
C5057 a_13059_46348# a_15143_45578# 0.262261f
C5058 a_13661_43548# a_9482_43914# 0.127225f
C5059 a_5807_45002# a_13556_45296# 0.017285f
C5060 a_n1151_42308# a_n2129_44697# 0.039834f
C5061 a_4883_46098# a_n2661_43370# 0.022462f
C5062 a_4905_42826# VDD 0.439034f
C5063 a_7845_44172# a_8333_44056# 0.065494f
C5064 a_n2293_42834# a_n2472_42826# 0.199703f
C5065 a_4651_46660# VDD 0.457722f
C5066 a_13259_45724# a_8696_44636# 0.259609f
C5067 a_1823_45246# a_1307_43914# 0.013371f
C5068 a_3483_46348# a_13777_45326# 0.027519f
C5069 a_5937_45572# a_7276_45260# 0.052629f
C5070 a_3090_45724# a_n2661_44458# 0.088502f
C5071 a_4915_47217# a_4883_46098# 0.024005f
C5072 a_10533_42308# a_10723_42308# 0.23663f
C5073 a_n3674_38216# a_n4064_40160# 0.02459f
C5074 a_n1177_43370# a_n447_43370# 0.010921f
C5075 a_n2267_43396# a_n2012_43396# 0.064178f
C5076 a_6945_45028# DATA[3] 0.014238f
C5077 a_n913_45002# a_3905_42558# 0.047606f
C5078 a_20107_45572# a_21188_45572# 0.102355f
C5079 a_20273_45572# a_21363_45546# 0.042415f
C5080 a_20841_45814# a_20623_45572# 0.209641f
C5081 a_n357_42282# a_18494_42460# 0.033084f
C5082 a_13249_42308# a_14180_45002# 0.014749f
C5083 a_16327_47482# a_19268_43646# 0.024286f
C5084 a_11453_44696# a_3090_45724# 0.232756f
C5085 a_n1925_46634# a_4646_46812# 0.089593f
C5086 a_12891_46348# a_6755_46942# 0.025465f
C5087 a_12861_44030# a_16721_46634# 0.070721f
C5088 a_6123_31319# VDD 0.533032f
C5089 a_5742_30871# C4_P_btm 0.03103f
C5090 a_18114_32519# a_13258_32519# 0.059438f
C5091 a_5891_43370# a_6761_42308# 0.010358f
C5092 a_18341_45572# VDD 0.2432f
C5093 a_10193_42453# a_3422_30871# 0.404849f
C5094 a_n1059_45260# a_5343_44458# 0.019826f
C5095 a_8696_44636# a_n2661_43922# 0.257466f
C5096 a_19692_46634# a_13467_32519# 0.015407f
C5097 a_12891_46348# a_8049_45260# 0.035062f
C5098 a_n1151_42308# a_6472_45840# 0.01357f
C5099 a_19692_46634# a_20273_46660# 0.02419f
C5100 a_4791_45118# a_2711_45572# 0.160646f
C5101 a_n2438_43548# a_n2956_39304# 0.014879f
C5102 C4_P_btm C0_dummy_P_btm 0.113156f
C5103 EN_VIN_BSTR_N C9_N_btm 0.226529f
C5104 C2_P_btm C1_P_btm 5.24136f
C5105 C3_P_btm C0_P_btm 0.409238f
C5106 EN_VIN_BSTR_P VDD 0.917665f
C5107 a_8975_43940# VDD 0.257588f
C5108 a_n1557_42282# a_n473_42460# 0.077371f
C5109 a_18479_45785# a_19319_43548# 0.102555f
C5110 a_19778_44110# a_11967_42832# 0.024799f
C5111 a_20692_30879# a_13467_32519# 0.051714f
C5112 a_n699_43396# a_3363_44484# 0.07346f
C5113 a_3232_43370# a_10729_43914# 0.090148f
C5114 a_11691_44458# a_17517_44484# 0.058911f
C5115 a_n1177_44458# a_n2661_43922# 0.010791f
C5116 a_n743_46660# a_16147_45260# 0.071228f
C5117 a_10903_43370# a_10809_44734# 0.353301f
C5118 a_3483_46348# a_5066_45546# 0.081087f
C5119 a_768_44030# a_2437_43646# 0.137571f
C5120 a_13887_32519# a_13258_32519# 0.054157f
C5121 a_5342_30871# a_5934_30871# 0.018148f
C5122 a_13467_32519# a_21613_42308# 0.053076f
C5123 a_n2810_45028# a_n3674_39304# 0.023324f
C5124 a_3357_43084# a_3935_42891# 0.025181f
C5125 a_n1331_43914# a_n984_44318# 0.051162f
C5126 a_n357_42282# a_133_42852# 0.011275f
C5127 a_n1099_45572# a_n356_45724# 0.070228f
C5128 a_n1079_45724# a_n1013_45572# 0.010598f
C5129 a_18479_47436# a_17517_44484# 0.017833f
C5130 a_13059_46348# a_13017_45260# 0.022433f
C5131 a_17715_44484# a_15861_45028# 0.184272f
C5132 a_n2661_45546# a_1609_45822# 0.02204f
C5133 a_n755_45592# a_3218_45724# 0.045755f
C5134 a_584_46384# a_2063_45854# 0.406382f
C5135 a_327_47204# a_n1151_42308# 0.013822f
C5136 a_n1741_47186# a_5815_47464# 0.021904f
C5137 a_2905_42968# VDD 0.142081f
C5138 a_n784_42308# a_6123_31319# 0.144274f
C5139 a_5342_30871# a_10890_34112# 0.013129f
C5140 a_3537_45260# a_5193_42852# 0.012016f
C5141 a_2711_45572# a_13258_32519# 0.02914f
C5142 a_n2956_38216# a_n4209_39304# 0.020992f
C5143 a_n1076_46494# VDD 0.294742f
C5144 a_n2017_45002# a_13291_42460# 0.042872f
C5145 a_20820_30879# VREF 0.195875f
C5146 a_n2661_42282# a_3626_43646# 0.02843f
C5147 a_14021_43940# a_19319_43548# 0.026713f
C5148 a_8696_44636# a_17478_45572# 0.185985f
C5149 a_2324_44458# a_949_44458# 0.323116f
C5150 a_n881_46662# a_171_46873# 0.018745f
C5151 a_n1613_43370# a_33_46660# 0.599895f
C5152 a_13661_43548# a_13747_46662# 0.095862f
C5153 a_15597_42852# VDD 0.239357f
C5154 a_n784_42308# EN_VIN_BSTR_P 0.051272f
C5155 a_n3565_39590# a_n4064_39616# 0.231239f
C5156 a_n97_42460# a_n1853_43023# 0.151542f
C5157 a_15095_43370# a_14955_43396# 0.130374f
C5158 a_10193_42453# VDD 2.18892f
C5159 a_13159_45002# a_9482_43914# 0.020865f
C5160 a_13017_45260# a_13556_45296# 0.049621f
C5161 a_3090_45724# a_9145_43396# 0.189557f
C5162 a_3232_43370# a_1423_45028# 0.396815f
C5163 a_768_44030# a_8199_44636# 0.026637f
C5164 a_11735_46660# a_12991_46634# 0.043475f
C5165 a_11901_46660# a_12469_46902# 0.175891f
C5166 a_12465_44636# a_6945_45028# 0.023497f
C5167 a_4883_46098# a_10809_44734# 0.068164f
C5168 a_n4209_38216# VIN_P 0.028615f
C5169 a_3754_39964# VDD 0.033808f
C5170 CAL_N a_22537_39537# 0.02334f
C5171 a_22589_40055# a_22848_40081# 0.010269f
C5172 a_10835_43094# a_10796_42968# 0.671797f
C5173 a_n1177_44458# a_n452_44636# 0.011059f
C5174 a_n913_45002# a_1414_42308# 0.021774f
C5175 a_11827_44484# a_16979_44734# 0.012885f
C5176 a_11691_44458# a_13720_44458# 0.029855f
C5177 a_n2293_45010# a_895_43940# 0.283316f
C5178 a_21188_46660# a_10809_44734# 0.010814f
C5179 a_n2497_47436# a_3232_43370# 0.04813f
C5180 a_4185_45028# a_4419_46090# 0.066314f
C5181 a_n971_45724# a_3065_45002# 0.220337f
C5182 a_5495_43940# VDD 0.173477f
C5183 a_743_42282# a_5934_30871# 0.020602f
C5184 a_18083_42858# a_18504_43218# 0.088127f
C5185 a_n2293_42834# a_n2129_43609# 0.017516f
C5186 a_n2293_43922# a_n1899_43946# 0.013114f
C5187 a_n2661_42834# a_n1549_44318# 0.011433f
C5188 a_n913_45002# a_12281_43396# 0.28203f
C5189 a_11967_42832# a_20159_44458# 0.056889f
C5190 a_6491_46660# VDD 0.436756f
C5191 a_11823_42460# a_12895_43230# 0.0142f
C5192 a_6945_45028# a_2711_45572# 0.036364f
C5193 a_584_46384# a_n2661_42834# 0.079307f
C5194 a_16327_47482# a_18248_44752# 0.050926f
C5195 a_12549_44172# a_11691_44458# 0.025825f
C5196 a_13661_43548# a_18911_45144# 0.03394f
C5197 a_5807_45002# a_19778_44110# 0.032504f
C5198 a_4883_46098# a_5883_43914# 0.01188f
C5199 a_16137_43396# VDD 0.483673f
C5200 a_15493_43396# a_15493_43940# 0.188034f
C5201 a_19862_44208# a_11341_43940# 0.07932f
C5202 a_3422_30871# a_3080_42308# 0.022126f
C5203 a_13259_45724# a_4958_30871# 0.054732f
C5204 a_n2956_39768# a_n4318_39768# 0.023595f
C5205 a_20205_31679# a_20447_31679# 9.01329f
C5206 a_n443_46116# a_171_46873# 0.029327f
C5207 a_6545_47178# a_n1925_46634# 0.02342f
C5208 a_18479_47436# a_12549_44172# 0.015281f
C5209 a_4883_46098# a_n881_46662# 0.193691f
C5210 a_n2109_47186# a_3877_44458# 0.021838f
C5211 a_10227_46804# a_15928_47570# 0.025137f
C5212 a_11599_46634# a_13661_43548# 0.078449f
C5213 a_17303_42282# a_17531_42308# 0.04615f
C5214 a_20692_30879# RST_Z 0.051046f
C5215 a_n2312_40392# a_n3674_39304# 0.025635f
C5216 a_11823_42460# a_11827_44484# 0.024482f
C5217 a_n2017_45002# a_2382_45260# 0.032443f
C5218 a_12549_44172# a_4190_30871# 0.270972f
C5219 a_768_44030# a_765_45546# 0.033731f
C5220 a_22959_47212# a_22959_46660# 0.025171f
C5221 a_12549_44172# a_17829_46910# 0.057751f
C5222 a_22775_42308# VDD 0.426061f
C5223 a_7754_39300# a_3754_38470# 0.082848f
C5224 a_n2840_42826# a_n3674_39304# 0.16082f
C5225 a_n4318_39768# a_n4318_37592# 0.023201f
C5226 a_n1991_42858# a_n1641_43230# 0.229804f
C5227 a_n2157_42858# a_n1076_43230# 0.102325f
C5228 a_n1853_43023# a_n901_43156# 0.081949f
C5229 a_16137_43396# a_16414_43172# 0.179708f
C5230 a_5691_45260# VDD 0.205518f
C5231 en_comp a_n2293_43922# 0.412872f
C5232 a_n967_45348# a_n2661_43922# 0.024232f
C5233 a_1423_45028# a_8975_43940# 0.331942f
C5234 a_1307_43914# a_16112_44458# 0.012033f
C5235 a_3232_43370# a_6109_44484# 0.072011f
C5236 a_10193_42453# a_10729_43914# 0.010339f
C5237 a_18587_45118# a_18911_45144# 0.010993f
C5238 a_5205_44484# a_5205_44734# 0.015405f
C5239 a_5111_44636# a_5891_43370# 0.702087f
C5240 a_21076_30879# a_17364_32525# 0.057544f
C5241 a_n2442_46660# a_n2810_45572# 0.045104f
C5242 a_12549_44172# a_n443_42852# 0.069091f
C5243 a_n2956_39768# a_n2956_38216# 0.043382f
C5244 a_2063_45854# a_8696_44636# 0.029184f
C5245 a_765_45546# a_1176_45822# 0.241847f
C5246 a_13059_46348# a_3483_46348# 0.319214f
C5247 a_14401_32519# a_13258_32519# 0.053694f
C5248 a_3422_30871# a_n1057_35014# 0.041712f
C5249 a_1307_43914# a_1443_43940# 0.042476f
C5250 w_10694_33990# a_10890_34112# 41.728897f
C5251 a_12861_44030# a_18494_42460# 0.021479f
C5252 a_5807_45002# a_9482_43914# 0.018229f
C5253 a_3147_46376# a_3316_45546# 0.012262f
C5254 a_3090_45724# a_15599_45572# 0.022054f
C5255 a_16327_47482# a_16922_45042# 0.060018f
C5256 a_3080_42308# VDD 0.849713f
C5257 a_3422_30871# a_14021_43940# 0.018792f
C5258 a_n2956_38216# a_n4318_37592# 0.023126f
C5259 a_4646_46812# VDD 2.53408f
C5260 a_13259_45724# a_16680_45572# 0.038605f
C5261 a_3483_46348# a_13556_45296# 0.375978f
C5262 a_4646_46812# a_7640_43914# 0.183308f
C5263 a_n2293_46634# a_14673_44172# 0.100552f
C5264 a_13747_46662# a_11967_42832# 0.021948f
C5265 a_1138_42852# a_1307_43914# 0.123153f
C5266 a_5937_45572# a_5205_44484# 0.481405f
C5267 a_9290_44172# a_5111_44636# 0.031975f
C5268 a_n443_46116# a_4883_46098# 0.037308f
C5269 a_14955_47212# a_11599_46634# 0.011007f
C5270 a_n1794_35082# a_7174_31319# 0.035143f
C5271 COMP_P a_22485_38105# 0.062482f
C5272 a_n1177_43370# a_n1352_43396# 0.233657f
C5273 a_n2129_43609# a_n2012_43396# 0.183186f
C5274 a_19862_44208# a_10341_43396# 0.028065f
C5275 a_20273_45572# a_20623_45572# 0.219856f
C5276 a_20107_45572# a_21363_45546# 0.043567f
C5277 a_n357_42282# a_18184_42460# 0.106442f
C5278 a_16327_47482# a_15743_43084# 1.21037f
C5279 a_21076_30879# a_19237_31679# 0.05495f
C5280 a_n1925_42282# a_n356_44636# 0.020589f
C5281 a_n1925_46634# a_3877_44458# 0.070082f
C5282 a_5807_45002# a_7715_46873# 0.029268f
C5283 a_11309_47204# a_6755_46942# 0.09972f
C5284 a_13507_46334# a_15227_44166# 0.235687f
C5285 a_12861_44030# a_16388_46812# 0.11634f
C5286 a_n4315_30879# a_n4209_37414# 0.039099f
C5287 a_n4334_38528# a_n4334_38304# 0.052468f
C5288 a_n3565_38502# a_n4209_38216# 5.84657f
C5289 a_n4209_38502# a_n3565_38216# 0.028468f
C5290 a_n2302_38778# a_n2216_38778# 0.011479f
C5291 a_7227_42308# VDD 0.296912f
C5292 a_5742_30871# C5_P_btm 0.089375f
C5293 a_18479_45785# VDD 0.536075f
C5294 a_n2017_45002# a_5343_44458# 0.027073f
C5295 a_6171_45002# a_16237_45028# 0.05704f
C5296 a_2063_45854# a_7227_45028# 0.021063f
C5297 a_19692_46634# a_20411_46873# 0.215749f
C5298 C5_P_btm C0_dummy_P_btm 0.11375f
C5299 EN_VIN_BSTR_N C8_N_btm 0.090252f
C5300 C3_P_btm C1_P_btm 8.06688f
C5301 C4_P_btm C0_P_btm 0.138331f
C5302 a_n1057_35014# VDD 0.336606f
C5303 a_10057_43914# VDD 0.399284f
C5304 a_n1557_42282# a_n961_42308# 0.041329f
C5305 a_3080_42308# a_n784_42308# 0.170007f
C5306 a_20205_31679# a_13467_32519# 0.051513f
C5307 a_n1917_44484# a_n2661_43922# 0.010578f
C5308 a_13507_46334# a_7174_31319# 0.041342f
C5309 a_n1613_43370# a_n2661_45010# 0.223356f
C5310 a_17583_46090# a_17715_44484# 0.22771f
C5311 a_4361_42308# a_21335_42336# 0.013772f
C5312 a_13467_32519# a_21887_42336# 0.011781f
C5313 a_14021_43940# VDD 1.60583f
C5314 a_3537_45260# a_5649_42852# 0.048691f
C5315 a_n1899_43946# a_n984_44318# 0.118759f
C5316 a_3357_43084# a_3681_42891# 0.052403f
C5317 a_8953_45546# a_5934_30871# 0.113715f
C5318 a_9804_47204# VDD 0.410522f
C5319 a_n2956_38680# a_n3674_37592# 0.026013f
C5320 a_380_45546# a_n356_45724# 0.088749f
C5321 a_n2661_45546# a_n443_42852# 0.141363f
C5322 a_17715_44484# a_8696_44636# 0.017149f
C5323 a_n755_45592# a_2957_45546# 0.044162f
C5324 a_n971_45724# a_4007_47204# 0.01992f
C5325 a_n785_47204# a_n1151_42308# 0.07743f
C5326 a_2124_47436# a_2063_45854# 0.074695f
C5327 a_n1741_47186# a_5129_47502# 0.012935f
C5328 a_n1794_35082# a_5932_42308# 0.033914f
C5329 a_2713_42308# a_2903_42308# 0.23738f
C5330 a_n2293_43922# a_n2157_42858# 0.040551f
C5331 a_11823_42460# a_13575_42558# 0.075921f
C5332 a_3537_45260# a_4649_42852# 0.065656f
C5333 a_2711_45572# a_19647_42308# 0.046367f
C5334 a_n2810_45572# a_n3565_39304# 0.030572f
C5335 a_n901_46420# VDD 0.518805f
C5336 a_20820_30879# VIN_N 0.049113f
C5337 a_21076_30879# EN_OFFSET_CAL 0.2809f
C5338 a_19692_46634# a_3422_30871# 0.208985f
C5339 a_2711_45572# a_3065_45002# 0.012727f
C5340 a_8696_44636# a_15861_45028# 0.26484f
C5341 a_16115_45572# a_16223_45938# 0.057222f
C5342 a_8128_46384# a_n1925_46634# 0.21095f
C5343 a_n1613_43370# a_171_46873# 0.11335f
C5344 a_5807_45002# a_13747_46662# 0.103485f
C5345 a_12549_44172# a_n2661_46634# 0.024531f
C5346 a_2063_45854# a_11813_46116# 0.093948f
C5347 a_n4334_39616# a_n4064_39616# 0.4504f
C5348 a_n4209_39590# a_n2302_39866# 0.406459f
C5349 a_n3565_39590# a_n2946_39866# 0.406088f
C5350 a_n3690_39616# a_n3420_39616# 0.431154f
C5351 a_14579_43548# a_10341_43396# 0.029139f
C5352 a_10695_43548# a_10849_43646# 0.010303f
C5353 a_14205_43396# a_14955_43396# 0.157423f
C5354 a_9145_43396# a_12281_43396# 0.032945f
C5355 a_n4318_39304# a_n4318_38680# 0.059432f
C5356 a_10180_45724# VDD 0.336512f
C5357 en_comp a_1107_38525# 0.206093f
C5358 a_13159_45002# a_13348_45260# 0.105274f
C5359 a_13017_45260# a_9482_43914# 0.048717f
C5360 a_21496_47436# a_10809_44734# 0.0112f
C5361 a_6755_46942# a_12156_46660# 0.013732f
C5362 a_10623_46897# a_10933_46660# 0.013793f
C5363 a_11735_46660# a_12251_46660# 0.105995f
C5364 a_8270_45546# a_3090_45724# 0.046518f
C5365 a_9804_47204# a_9823_46155# 0.063581f
C5366 a_n4064_37440# EN_VIN_BSTR_P 0.03202f
C5367 a_22589_40055# a_22527_39145# 0.130029f
C5368 a_22537_40625# a_22581_37893# 0.656829f
C5369 a_10518_42984# a_10796_42968# 0.118759f
C5370 a_3422_30871# a_21613_42308# 0.027998f
C5371 a_n1059_45260# a_1414_42308# 0.031011f
C5372 a_n1177_44458# a_n1352_44484# 0.233657f
C5373 a_11827_44484# a_14539_43914# 0.044058f
C5374 a_3357_43084# a_5663_43940# 0.015908f
C5375 a_18911_45144# a_18989_43940# 0.016276f
C5376 a_11691_44458# a_13076_44458# 0.03093f
C5377 a_6575_47204# a_2437_43646# 0.029543f
C5378 a_11415_45002# a_2324_44458# 0.097878f
C5379 a_21363_46634# a_10809_44734# 0.012784f
C5380 a_n1151_42308# a_n913_45002# 0.395136f
C5381 a_n971_45724# a_2680_45002# 0.108251f
C5382 a_n2109_47186# a_5111_44636# 0.017519f
C5383 a_13747_46662# a_15143_45578# 0.040557f
C5384 a_15567_42826# a_15597_42852# 0.025037f
C5385 a_5013_44260# VDD 0.198233f
C5386 a_10057_43914# a_10729_43914# 0.063518f
C5387 a_n2661_42834# a_n1331_43914# 0.01077f
C5388 a_3232_43370# a_3457_43396# 0.131408f
C5389 a_3537_45260# a_8685_43396# 0.023888f
C5390 a_n1059_45260# a_12281_43396# 0.025081f
C5391 a_n2293_42834# a_n2433_43396# 0.025997f
C5392 a_6545_47178# VDD 0.386368f
C5393 a_n1151_42308# CLK 0.022274f
C5394 a_6151_47436# RST_Z 0.010195f
C5395 a_11967_42832# a_19615_44636# 0.065767f
C5396 a_13661_43548# a_18587_45118# 0.087703f
C5397 a_6755_46942# a_6171_45002# 0.026424f
C5398 a_16327_47482# a_17970_44736# 0.219775f
C5399 a_n2438_43548# a_n2661_43370# 0.147387f
C5400 a_12891_46348# a_11691_44458# 0.141379f
C5401 a_4646_46812# a_1423_45028# 0.415897f
C5402 a_4190_30871# EN_VIN_BSTR_N 0.043599f
C5403 a_19328_44172# a_15493_43940# 0.062184f
C5404 a_19862_44208# a_21115_43940# 0.064973f
C5405 a_12429_44172# a_12603_44260# 0.011572f
C5406 a_20365_43914# a_20623_43914# 0.22264f
C5407 a_19692_46634# VDD 2.53528f
C5408 a_6755_46942# a_14673_44172# 0.050772f
C5409 a_20692_30879# a_19963_31679# 0.051965f
C5410 a_8049_45260# a_6171_45002# 0.048422f
C5411 a_13259_45724# en_comp 0.19355f
C5412 a_n2661_45546# a_2437_43646# 0.028152f
C5413 a_n971_45724# a_n229_43646# 0.059197f
C5414 a_11962_45724# a_11682_45822# 0.014813f
C5415 a_n1151_42308# a_2107_46812# 0.073605f
C5416 a_6151_47436# a_n1925_46634# 0.052327f
C5417 a_4883_46098# a_n1613_43370# 0.025959f
C5418 a_12861_44030# a_19321_45002# 0.10527f
C5419 a_10227_46804# a_768_44030# 0.050994f
C5420 a_11599_46634# a_5807_45002# 0.303048f
C5421 a_4958_30871# a_17531_42308# 0.192941f
C5422 a_14021_43940# a_21487_43396# 0.023941f
C5423 a_20692_30879# VDD 0.508982f
C5424 a_20205_31679# RST_Z 0.049474f
C5425 a_18184_42460# a_22400_42852# 0.16156f
C5426 a_n967_45348# a_n955_45028# 0.014419f
C5427 a_3357_43084# a_3232_43370# 0.118744f
C5428 a_12549_44172# a_765_45546# 0.118284f
C5429 SMPL_ON_N a_21076_30879# 0.03043f
C5430 a_21613_42308# VDD 0.27399f
C5431 a_n3420_39072# EN_VIN_BSTR_P 0.814839f
C5432 a_n1991_42858# a_n1423_42826# 0.186387f
C5433 a_n2157_42858# a_n901_43156# 0.043475f
C5434 a_n1853_43023# a_n1641_43230# 0.036072f
C5435 a_4927_45028# VDD 0.159822f
C5436 a_n3674_39768# a_n3674_38216# 0.02323f
C5437 a_1414_42308# a_1606_42308# 0.056716f
C5438 a_n967_45348# a_n2661_42834# 0.027185f
C5439 en_comp a_n2661_43922# 0.237031f
C5440 a_16327_47482# a_20256_43172# 0.054992f
C5441 a_15227_44166# a_17701_42308# 0.172697f
C5442 w_1575_34786# a_5934_30871# 0.097232f
C5443 a_327_44734# a_556_44484# 0.033015f
C5444 a_7499_43078# a_11750_44172# 0.195997f
C5445 a_5147_45002# a_5891_43370# 0.049542f
C5446 a_11599_46634# a_15143_45578# 0.028879f
C5447 a_765_45546# a_1208_46090# 0.134766f
C5448 a_1307_43914# a_1241_43940# 0.038832f
C5449 a_3357_43084# a_4905_42826# 0.062628f
C5450 a_7499_43078# a_4361_42308# 0.04291f
C5451 a_n967_45348# a_n1352_43396# 0.010028f
C5452 a_12861_44030# a_18184_42460# 0.266953f
C5453 a_2324_44458# a_13259_45724# 0.068761f
C5454 a_768_44030# a_1307_43914# 1.13357f
C5455 a_n1151_42308# a_n2661_44458# 0.030695f
C5456 a_3147_46376# a_3218_45724# 0.0111f
C5457 a_13059_46348# a_13249_42308# 0.306398f
C5458 a_n2293_46634# a_3232_43370# 0.046281f
C5459 a_n4318_38680# a_n4334_38528# 0.08371f
C5460 a_4699_43561# VDD 0.262218f
C5461 a_7845_44172# a_7911_44260# 0.010598f
C5462 a_n2293_43922# a_n2267_43396# 0.020404f
C5463 a_n357_42282# a_20753_42852# 0.013117f
C5464 a_3877_44458# VDD 0.786903f
C5465 a_13259_45724# a_16855_45546# 0.067694f
C5466 a_3483_46348# a_9482_43914# 0.130172f
C5467 a_8953_45546# a_6171_45002# 0.0298f
C5468 a_5937_45572# a_6431_45366# 0.129839f
C5469 a_4646_46812# a_6109_44484# 0.010238f
C5470 a_13661_43548# a_11967_42832# 0.165876f
C5471 a_4791_45118# a_4883_46098# 0.135093f
C5472 a_4915_47217# a_13507_46334# 0.032373f
C5473 a_12861_44030# a_15811_47375# 0.144648f
C5474 a_10545_42558# a_10533_42308# 0.011812f
C5475 a_n4318_38216# a_n4064_40160# 0.052465f
C5476 a_n1761_44111# a_n901_43156# 0.013702f
C5477 a_n2433_43396# a_n2012_43396# 0.089677f
C5478 a_n1736_46482# VDD 0.083417f
C5479 a_18184_42460# a_22223_42860# 0.03037f
C5480 a_11967_42832# a_10835_43094# 0.263495f
C5481 a_13249_42308# a_13556_45296# 0.059719f
C5482 a_n2293_46634# a_4905_42826# 0.024749f
C5483 a_768_44030# a_9396_43370# 0.010156f
C5484 a_4791_45118# a_5649_42852# 0.075725f
C5485 a_n1613_43370# a_8685_43396# 0.016726f
C5486 a_20107_45572# a_20623_45572# 0.103168f
C5487 a_20273_45572# a_20841_45814# 0.175891f
C5488 a_2324_44458# a_n2661_43922# 0.088002f
C5489 a_526_44458# a_n356_44636# 0.142971f
C5490 a_16327_47482# a_18783_43370# 0.026485f
C5491 a_11309_47204# a_10249_46116# 0.033926f
C5492 a_6575_47204# a_765_45546# 0.061901f
C5493 a_12861_44030# a_13059_46348# 0.504219f
C5494 a_1273_38525# VDAC_Pi 0.035744f
C5495 a_6761_42308# VDD 0.259312f
C5496 a_5742_30871# C6_P_btm 0.170624f
C5497 a_18429_43548# a_16823_43084# 0.130506f
C5498 a_18175_45572# VDD 0.38478f
C5499 a_n1059_45260# a_n699_43396# 0.021143f
C5500 a_327_44734# a_n2661_44458# 0.027103f
C5501 a_19692_46634# a_21487_43396# 0.016698f
C5502 a_5009_45028# a_5093_45028# 0.092725f
C5503 a_14180_46812# a_13059_46348# 0.074456f
C5504 a_2063_45854# a_6598_45938# 0.018518f
C5505 a_19692_46634# a_20107_46660# 0.126737f
C5506 C6_P_btm C0_dummy_P_btm 0.1194f
C5507 EN_VIN_BSTR_N C7_N_btm 0.115875f
C5508 C3_P_btm C2_P_btm 5.99608f
C5509 C5_P_btm C0_P_btm 0.138093f
C5510 C4_P_btm C1_P_btm 0.128167f
C5511 a_n1696_34930# VDD 2.24623f
C5512 a_10440_44484# VDD 0.159539f
C5513 a_n1557_42282# a_n1329_42308# 0.075734f
C5514 a_2779_44458# a_3363_44484# 0.020864f
C5515 a_13747_46662# a_20107_45572# 0.012917f
C5516 a_12861_44030# a_13556_45296# 0.028687f
C5517 a_22959_47212# a_413_45260# 0.024836f
C5518 a_4361_42308# a_7174_31319# 0.024432f
C5519 a_5649_42852# a_13258_32519# 0.040931f
C5520 a_10341_42308# a_9803_42558# 0.108853f
C5521 a_5534_30871# a_5934_30871# 0.018227f
C5522 a_5342_30871# a_6123_31319# 0.018227f
C5523 a_n967_45348# a_n1423_42826# 0.010397f
C5524 a_8128_46384# VDD 0.403575f
C5525 a_n2956_39304# a_n3674_37592# 0.026377f
C5526 a_n1761_44111# a_n984_44318# 0.056404f
C5527 a_n1899_43946# a_n809_44244# 0.042737f
C5528 a_n1331_43914# a_n1549_44318# 0.209641f
C5529 a_3357_43084# a_2905_42968# 0.025927f
C5530 a_13661_43548# a_18989_43940# 0.039099f
C5531 a_n452_45724# a_n356_45724# 0.318161f
C5532 a_n755_45592# a_1848_45724# 0.030306f
C5533 a_5534_30871# a_10890_34112# 0.010397f
C5534 a_n971_45724# a_3815_47204# 0.04068f
C5535 a_2124_47436# a_584_46384# 0.220021f
C5536 a_n1741_47186# a_4915_47217# 0.128899f
C5537 a_1847_42826# VDD 0.527555f
C5538 a_5342_30871# EN_VIN_BSTR_P 0.010795f
C5539 a_n2661_42282# a_2982_43646# 0.076578f
C5540 a_5745_43940# a_5829_43940# 0.092725f
C5541 a_11823_42460# a_13070_42354# 0.077142f
C5542 a_2711_45572# a_19511_42282# 0.234026f
C5543 a_n1641_46494# VDD 0.226065f
C5544 a_n913_45002# a_11136_42852# 0.026537f
C5545 a_22959_46660# EN_OFFSET_CAL 0.050989f
C5546 a_17339_46660# a_17517_44484# 0.020067f
C5547 a_16333_45814# a_16223_45938# 0.097745f
C5548 a_16115_45572# a_16020_45572# 0.049827f
C5549 a_5807_45002# a_13661_43548# 0.062335f
C5550 a_n1613_43370# a_n133_46660# 0.347805f
C5551 a_n881_46662# a_n2438_43548# 0.080298f
C5552 a_n4209_39590# a_n4064_39616# 0.269818f
C5553 a_n3565_39590# a_n3420_39616# 0.281955f
C5554 a_n4318_39304# a_n3674_39304# 2.9537f
C5555 a_4905_42826# a_743_42282# 0.0175f
C5556 a_10695_43548# a_10765_43646# 0.011552f
C5557 a_10053_45546# VDD 0.150582f
C5558 a_14205_43396# a_15095_43370# 0.086245f
C5559 a_7499_43078# a_5891_43370# 1.00892f
C5560 a_13017_45260# a_13348_45260# 0.044101f
C5561 a_10903_43370# a_11173_44260# 0.035423f
C5562 a_n913_45002# a_n2293_42834# 0.055202f
C5563 a_13507_46334# a_10809_44734# 0.603934f
C5564 a_n2438_43548# a_n2157_46122# 0.270054f
C5565 a_768_44030# a_8016_46348# 0.034453f
C5566 a_9804_47204# a_9569_46155# 0.040648f
C5567 a_11813_46116# a_11901_46660# 0.211542f
C5568 a_11735_46660# a_12469_46902# 0.053479f
C5569 a_4883_46098# a_6945_45028# 0.083863f
C5570 a_22589_40599# a_22581_37893# 0.365664f
C5571 CAL_N a_22613_38993# 0.010642f
C5572 a_10518_42984# a_10835_43094# 0.102355f
C5573 a_10083_42826# a_10796_42968# 0.042737f
C5574 a_11691_44458# a_12883_44458# 0.058264f
C5575 a_n2017_45002# a_1414_42308# 0.015426f
C5576 a_n2661_44458# a_4223_44672# 0.019953f
C5577 a_n357_42282# a_6031_43396# 0.012855f
C5578 a_n443_42852# a_n1557_42282# 0.078868f
C5579 a_n2661_45010# a_895_43940# 0.020382f
C5580 a_n2109_47186# a_5147_45002# 0.05864f
C5581 a_13747_46662# a_14495_45572# 0.288916f
C5582 a_n1151_42308# a_n1059_45260# 0.16984f
C5583 a_18597_46090# a_18341_45572# 0.010006f
C5584 a_11599_46634# a_20107_45572# 0.246047f
C5585 a_n2293_46634# a_10193_42453# 0.037794f
C5586 a_3483_46348# a_4419_46090# 0.218073f
C5587 a_n971_45724# a_2382_45260# 0.019144f
C5588 a_n2661_46634# a_11322_45546# 0.059929f
C5589 a_6491_46660# a_3357_43084# 0.014978f
C5590 a_743_42282# a_6123_31319# 0.018532f
C5591 a_4190_30871# a_5934_30871# 0.020923f
C5592 a_5244_44056# VDD 0.146618f
C5593 a_4361_42308# a_5932_42308# 0.072603f
C5594 a_10057_43914# a_10405_44172# 0.028414f
C5595 a_n2293_43922# a_n2065_43946# 0.02752f
C5596 a_n2661_42834# a_n1899_43946# 0.049432f
C5597 a_3232_43370# a_2813_43396# 0.05929f
C5598 a_10193_42453# a_5342_30871# 0.151919f
C5599 a_n2017_45002# a_12281_43396# 0.028019f
C5600 a_17517_44484# a_18579_44172# 0.031747f
C5601 a_11823_42460# a_12545_42858# 0.039145f
C5602 a_375_42282# a_n1557_42282# 0.450989f
C5603 a_6151_47436# VDD 4.39915f
C5604 a_4007_47204# DATA[2] 0.337596f
C5605 a_9290_44172# a_7499_43078# 0.597117f
C5606 a_8953_45546# a_8746_45002# 0.020026f
C5607 a_16327_47482# a_17767_44458# 0.269619f
C5608 a_3877_44458# a_1423_45028# 0.022537f
C5609 a_526_44458# a_3503_45724# 0.06484f
C5610 a_4190_30871# a_10890_34112# 0.032471f
C5611 a_18451_43940# a_15493_43940# 0.051906f
C5612 a_15493_43396# a_11341_43940# 0.020569f
C5613 a_19862_44208# a_20935_43940# 0.03846f
C5614 a_14539_43914# a_16823_43084# 0.058282f
C5615 a_n4318_40392# a_n4318_38680# 0.023692f
C5616 a_12429_44172# a_12495_44260# 0.012714f
C5617 a_19466_46812# VDD 0.664497f
C5618 a_n2956_39304# a_n2302_39072# 0.040755f
C5619 a_20205_31679# a_19963_31679# 9.023429f
C5620 a_10053_45546# a_10306_45572# 0.011897f
C5621 a_3160_47472# a_2107_46812# 0.041673f
C5622 a_n2497_47436# a_3877_44458# 0.024435f
C5623 a_n971_45724# a_3524_46660# 0.016598f
C5624 a_10227_46804# a_12549_44172# 0.360691f
C5625 a_13507_46334# a_n881_46662# 0.019152f
C5626 a_4915_47217# a_n743_46660# 0.026159f
C5627 a_n443_46116# a_n2438_43548# 0.070894f
C5628 a_4958_30871# a_17303_42282# 0.168656f
C5629 a_22959_43948# a_22959_43396# 0.025171f
C5630 a_14021_43940# a_20556_43646# 0.085306f
C5631 a_20205_31679# VDD 0.74083f
C5632 a_n1059_45260# a_18214_42558# 0.020063f
C5633 a_5937_45572# a_6453_43914# 0.144397f
C5634 a_20202_43084# a_19862_44208# 0.058613f
C5635 a_10193_42453# a_16237_45028# 0.049386f
C5636 a_3357_43084# a_5691_45260# 0.011637f
C5637 a_n863_45724# a_n23_44458# 0.056041f
C5638 a_12891_46348# a_765_45546# 0.041192f
C5639 a_12549_44172# a_17339_46660# 0.081298f
C5640 a_4646_46812# a_6969_46634# 0.072545f
C5641 a_n1741_47186# a_10809_44734# 0.332771f
C5642 a_2063_45854# a_2324_44458# 0.028153f
C5643 a_11453_44696# a_12741_44636# 1.02327f
C5644 a_21887_42336# VDD 0.210392f
C5645 a_n2157_42858# a_n1641_43230# 0.110532f
C5646 a_n1853_43023# a_n1423_42826# 0.022091f
C5647 a_413_45260# CLK 0.033653f
C5648 a_5111_44636# VDD 1.28013f
C5649 a_n4318_39768# a_n3674_38216# 0.023361f
C5650 en_comp a_n2661_42834# 0.080292f
C5651 a_16327_47482# a_18707_42852# 0.012993f
C5652 a_15227_44166# a_17595_43084# 0.041195f
C5653 a_18315_45260# a_18587_45118# 0.13675f
C5654 a_16922_45042# a_18494_42460# 0.242236f
C5655 a_n2293_42834# a_n2661_44458# 0.0289f
C5656 a_7499_43078# a_10807_43548# 0.119721f
C5657 a_21076_30879# a_14209_32519# 0.055087f
C5658 a_4520_42826# a_4743_43172# 0.011458f
C5659 a_n357_42282# a_10796_42968# 0.048375f
C5660 a_3357_43084# a_3080_42308# 0.233522f
C5661 a_n967_45348# a_n1177_43370# 0.013627f
C5662 a_10193_42453# a_743_42282# 1.1645f
C5663 a_18989_43940# a_11967_42832# 0.039137f
C5664 a_12861_44030# a_19778_44110# 0.113118f
C5665 a_12549_44172# a_1307_43914# 1.82879f
C5666 a_4185_45028# a_n755_45592# 0.024134f
C5667 a_4646_46812# a_3357_43084# 0.024669f
C5668 a_2107_46812# a_413_45260# 0.032665f
C5669 a_4235_43370# VDD 0.229422f
C5670 a_n4318_38680# a_n4209_38502# 0.105064f
C5671 a_22959_44484# a_22959_43948# 0.026152f
C5672 a_n356_44636# a_3626_43646# 0.073377f
C5673 a_18494_42460# a_15743_43084# 0.027791f
C5674 a_n2293_43922# a_n2129_43609# 0.028035f
C5675 a_n2956_38216# a_n3674_38216# 0.028821f
C5676 a_13259_45724# a_16115_45572# 0.035684f
C5677 a_22959_46124# a_20447_31679# 0.015464f
C5678 a_12549_44172# a_18579_44172# 0.154956f
C5679 a_3483_46348# a_13348_45260# 0.041217f
C5680 a_5937_45572# a_6171_45002# 0.206948f
C5681 a_8953_45546# a_3232_43370# 0.019509f
C5682 a_8049_45260# a_18341_45572# 0.021945f
C5683 a_n1741_47186# a_n881_46662# 0.179671f
C5684 a_n1699_43638# a_n1352_43396# 0.051162f
C5685 a_15493_43396# a_10341_43396# 0.039468f
C5686 a_n2956_38680# VDD 0.871805f
C5687 a_n913_45002# a_5379_42460# 0.179494f
C5688 a_18184_42460# a_22165_42308# 0.026631f
C5689 a_13249_42308# a_9482_43914# 0.061734f
C5690 a_n2293_46634# a_3080_42308# 0.039273f
C5691 a_21076_30879# a_17730_32519# 0.054832f
C5692 a_20107_45572# a_20841_45814# 0.053479f
C5693 a_16327_47482# a_18525_43370# 0.059008f
C5694 a_n2293_46634# a_4646_46812# 0.135642f
C5695 a_n2661_46634# a_4817_46660# 0.047477f
C5696 a_5807_45002# a_5257_43370# 0.683815f
C5697 a_13507_46334# a_17609_46634# 0.01055f
C5698 a_12861_44030# a_15227_46910# 0.050112f
C5699 a_n2497_47436# a_n1641_46494# 0.020605f
C5700 a_n4209_38502# a_n4209_38216# 0.041706f
C5701 a_5742_30871# C7_P_btm 0.04157f
C5702 a_16137_43396# a_743_42282# 0.183525f
C5703 en_comp a_22527_39145# 0.393507f
C5704 a_17324_43396# a_16823_43084# 0.038999f
C5705 a_16147_45260# VDD 0.197706f
C5706 a_3080_42308# a_5342_30871# 0.01896f
C5707 a_413_45260# a_n2661_44458# 0.69469f
C5708 a_n967_45348# a_n1177_44458# 0.012502f
C5709 a_19692_46634# a_20556_43646# 0.118928f
C5710 a_6171_45002# a_11691_44458# 0.022104f
C5711 a_14035_46660# a_13059_46348# 0.072321f
C5712 a_n743_46660# a_10809_44734# 0.032324f
C5713 a_n2312_38680# a_n2956_38680# 6.25577f
C5714 a_2063_45854# a_6667_45809# 0.029741f
C5715 a_19692_46634# a_19551_46910# 0.0536f
C5716 a_11453_44696# a_16375_45002# 0.104273f
C5717 C7_P_btm C0_dummy_P_btm 0.119061f
C5718 EN_VIN_BSTR_N C6_N_btm 0.118916f
C5719 C6_P_btm C0_P_btm 0.139059f
C5720 C5_P_btm C1_P_btm 0.127408f
C5721 C4_P_btm C2_P_btm 7.72909f
C5722 a_n1550_35448# VDD 0.366274f
C5723 a_10334_44484# VDD 0.19332f
C5724 a_n1557_42282# COMP_P 0.123881f
C5725 a_1307_43914# a_7542_44172# 0.022371f
C5726 a_11691_44458# a_14673_44172# 0.371587f
C5727 a_n2267_44484# a_n2661_43922# 0.010057f
C5728 a_14976_45028# a_2711_45572# 0.025742f
C5729 a_12861_44030# a_9482_43914# 0.021886f
C5730 a_15682_46116# a_17583_46090# 0.013015f
C5731 a_11453_44696# a_413_45260# 0.032816f
C5732 a_4361_42308# a_20712_42282# 0.013294f
C5733 a_13678_32519# a_13258_32519# 0.055554f
C5734 a_n967_45348# a_n1991_42858# 0.034664f
C5735 a_n913_45002# a_n13_43084# 0.042137f
C5736 a_n1761_44111# a_n809_44244# 0.038277f
C5737 a_n2065_43946# a_n984_44318# 0.102325f
C5738 a_n1899_43946# a_n1549_44318# 0.218775f
C5739 a_8199_44636# a_5934_30871# 0.159294f
C5740 a_n2293_46634# a_10057_43914# 0.01757f
C5741 a_8049_45260# a_10193_42453# 0.082788f
C5742 a_12861_44030# a_20159_44458# 0.014378f
C5743 a_n755_45592# a_997_45618# 0.133124f
C5744 a_n971_45724# a_3785_47178# 0.032234f
C5745 a_n237_47217# a_n1151_42308# 0.63407f
C5746 a_n1741_47186# a_n443_46116# 0.053258f
C5747 a_n2109_47186# a_5129_47502# 0.021297f
C5748 a_791_42968# VDD 0.128737f
C5749 a_1755_42282# a_5379_42460# 0.045501f
C5750 a_2725_42558# a_2713_42308# 0.01129f
C5751 COMP_P a_5934_30871# 0.028651f
C5752 a_11823_42460# a_12563_42308# 0.039858f
C5753 a_n1423_46090# VDD 0.227012f
C5754 a_12741_44636# EN_OFFSET_CAL 0.230064f
C5755 a_n2810_45572# a_n4209_39304# 0.020327f
C5756 a_15765_45572# a_16223_45938# 0.027606f
C5757 a_n2661_45546# a_1307_43914# 0.021108f
C5758 a_n2293_46634# a_14021_43940# 0.202404f
C5759 a_8953_45546# a_8975_43940# 0.02155f
C5760 a_11309_47204# a_n2661_46634# 0.042272f
C5761 a_2063_45854# a_11186_47026# 0.012485f
C5762 a_n971_45724# a_3090_45724# 0.071442f
C5763 a_n1151_42308# a_8270_45546# 0.01803f
C5764 a_n881_46662# a_n743_46660# 0.527182f
C5765 a_n1613_43370# a_n2438_43548# 1.04064f
C5766 COMP_P a_10890_34112# 0.011687f
C5767 a_n3565_39590# a_n3690_39616# 0.246863f
C5768 a_n4334_39616# a_n3420_39616# 0.015897f
C5769 a_n4209_39590# a_n2946_39866# 0.022704f
C5770 a_3080_42308# a_743_42282# 0.069641f
C5771 a_9049_44484# VDD 0.680993f
C5772 a_3429_45260# a_3495_45348# 0.010598f
C5773 a_13017_45260# a_13159_45002# 0.160415f
C5774 a_5111_44636# a_1423_45028# 0.028542f
C5775 a_10903_43370# a_10555_44260# 0.011277f
C5776 a_21076_30879# a_17538_32519# 0.054805f
C5777 a_526_44458# a_3499_42826# 0.089844f
C5778 a_n1059_45260# a_n2293_42834# 0.035031f
C5779 a_13507_46334# a_22223_46124# 0.024274f
C5780 a_n2438_43548# a_n2293_46098# 0.409291f
C5781 a_9804_47204# a_9625_46129# 0.037672f
C5782 a_11735_46660# a_11901_46660# 0.579036f
C5783 a_13661_43548# a_3483_46348# 0.381471f
C5784 a_4817_46660# a_765_45546# 0.010165f
C5785 a_4883_46098# a_21137_46414# 0.010468f
C5786 CAL_N a_22581_37893# 0.023534f
C5787 a_22537_40625# a_22527_39145# 0.245895f
C5788 a_n3420_37440# EN_VIN_BSTR_P 0.040234f
C5789 a_10083_42826# a_10835_43094# 0.043619f
C5790 a_11691_44458# a_12607_44458# 0.042423f
C5791 a_n1699_44726# a_n1352_44484# 0.051162f
C5792 a_413_45260# a_19237_31679# 0.119197f
C5793 a_n2293_45010# a_453_43940# 0.181603f
C5794 a_13259_45724# a_13667_43396# 0.160676f
C5795 a_n2661_44458# a_2779_44458# 0.011596f
C5796 a_13747_46662# a_13249_42308# 0.134714f
C5797 a_n1151_42308# a_n2017_45002# 0.058036f
C5798 a_n2661_46634# a_10490_45724# 0.01771f
C5799 a_3483_46348# a_4185_45028# 0.430982f
C5800 a_3905_42865# VDD 0.788273f
C5801 a_n2293_43922# a_n2472_43914# 0.189122f
C5802 a_n2661_43922# a_n2065_43946# 0.013023f
C5803 a_n2661_42834# a_n1761_44111# 0.073205f
C5804 a_8975_43940# a_9028_43914# 0.184602f
C5805 a_10057_43914# a_9672_43914# 0.143523f
C5806 a_11823_42460# a_12089_42308# 0.335983f
C5807 a_19006_44850# a_11967_42832# 0.013801f
C5808 a_4185_45028# a_14097_32519# 0.020305f
C5809 a_5815_47464# VDD 0.399354f
C5810 a_3815_47204# DATA[2] 0.022461f
C5811 a_19321_45002# a_16922_45042# 0.493823f
C5812 a_768_44030# a_11827_44484# 0.831344f
C5813 a_8199_44636# a_10490_45724# 0.019372f
C5814 a_5937_45572# a_8746_45002# 0.121678f
C5815 a_19692_46634# a_3357_43084# 0.046179f
C5816 a_526_44458# a_3316_45546# 0.128261f
C5817 a_20269_44172# a_20365_43914# 0.419086f
C5818 a_18326_43940# a_15493_43940# 0.075033f
C5819 a_19862_44208# a_20623_43914# 0.023134f
C5820 a_n4318_40392# a_n3674_39304# 0.024125f
C5821 a_n2956_39304# a_n4064_39072# 0.054199f
C5822 a_19333_46634# VDD 0.199048f
C5823 a_3090_45724# a_9313_44734# 2.43867f
C5824 a_11525_45546# a_11682_45822# 0.18824f
C5825 a_9290_44172# a_n2661_43370# 0.185465f
C5826 a_18597_46090# a_14021_43940# 0.0185f
C5827 a_10053_45546# a_10216_45572# 0.011381f
C5828 a_21076_30879# a_19721_31679# 0.05488f
C5829 a_2905_45572# a_2107_46812# 0.031826f
C5830 a_16023_47582# a_16119_47582# 0.013793f
C5831 a_n971_45724# a_3699_46634# 0.024384f
C5832 a_12861_44030# a_13747_46662# 0.139424f
C5833 a_10227_46804# a_12891_46348# 0.058451f
C5834 a_n443_46116# a_n743_46660# 0.532861f
C5835 a_18494_42460# a_20256_43172# 0.052522f
C5836 a_5937_45572# a_5663_43940# 0.177912f
C5837 a_10193_42453# a_20193_45348# 0.305022f
C5838 a_n863_45724# a_n356_44636# 0.301674f
C5839 a_11309_47204# a_765_45546# 0.03506f
C5840 a_4646_46812# a_6755_46942# 0.362783f
C5841 a_3877_44458# a_6969_46634# 0.101189f
C5842 a_13747_46662# a_14180_46812# 0.021289f
C5843 a_21335_42336# VDD 0.199586f
C5844 a_4958_30871# VCM 0.642743f
C5845 a_7174_31319# RST_Z 0.216004f
C5846 a_n1853_43023# a_n1991_42858# 0.237526f
C5847 a_n2157_42858# a_n1423_42826# 0.07009f
C5848 a_5147_45002# VDD 0.574918f
C5849 a_n3674_39768# a_n4318_38216# 0.032347f
C5850 a_413_45260# EN_OFFSET_CAL 0.114452f
C5851 a_20820_30879# a_17364_32525# 0.055604f
C5852 a_16922_45042# a_18184_42460# 0.028064f
C5853 a_7499_43078# a_10949_43914# 0.152939f
C5854 w_1575_34786# a_6123_31319# 0.024772f
C5855 a_n2956_39768# a_n2810_45572# 0.043168f
C5856 a_4520_42826# a_4649_43172# 0.010132f
C5857 a_n357_42282# a_10835_43094# 0.02434f
C5858 a_18374_44850# a_11967_42832# 0.053726f
C5859 a_18989_43940# a_19006_44850# 0.168452f
C5860 a_4185_45028# a_22959_42860# 0.013205f
C5861 w_1575_34786# EN_VIN_BSTR_P 3.97869f
C5862 a_12861_44030# a_18911_45144# 0.169f
C5863 a_4185_45028# a_n357_42282# 0.023019f
C5864 a_3877_44458# a_3357_43084# 0.02473f
C5865 a_13059_46348# a_13527_45546# 0.017655f
C5866 a_n2661_46634# a_6171_45002# 0.042529f
C5867 a_4093_43548# VDD 0.216874f
C5868 a_n2293_43922# a_n2433_43396# 0.028793f
C5869 a_n2810_45572# a_n4318_37592# 0.023163f
C5870 a_18184_42460# a_15743_43084# 0.182123f
C5871 a_n2661_42834# a_n2267_43396# 0.014077f
C5872 a_13259_45724# a_16333_45814# 0.02201f
C5873 a_3483_46348# a_13159_45002# 0.017316f
C5874 a_5937_45572# a_3232_43370# 0.662525f
C5875 a_8199_44636# a_6171_45002# 0.163434f
C5876 a_22959_46124# a_22959_45572# 0.025171f
C5877 a_12861_44030# a_11599_46634# 0.169929f
C5878 a_n1741_47186# a_n1613_43370# 0.018791f
C5879 a_n3674_38680# a_n4064_40160# 0.022279f
C5880 a_n2267_43396# a_n1352_43396# 0.124988f
C5881 a_n2129_43609# a_n447_43370# 0.119518f
C5882 a_n2956_39304# VDD 0.455981f
C5883 a_n913_45002# a_5267_42460# 0.081794f
C5884 a_18184_42460# a_21671_42860# 0.021213f
C5885 a_16327_47482# a_18429_43548# 0.057366f
C5886 a_20107_45572# a_20273_45572# 0.667378f
C5887 a_3483_46348# a_11967_42832# 0.264293f
C5888 a_20820_30879# a_19237_31679# 0.053048f
C5889 a_9049_44484# a_1423_45028# 0.024539f
C5890 a_1983_46706# a_n2661_46098# 0.147223f
C5891 a_9804_47204# a_6755_46942# 0.028571f
C5892 a_n2661_46634# a_4955_46873# 0.03751f
C5893 a_4883_46098# a_15368_46634# 0.023335f
C5894 a_2107_46812# a_2443_46660# 0.013591f
C5895 a_18597_46090# a_19692_46634# 0.019861f
C5896 a_10227_46804# a_12359_47026# 0.012196f
C5897 a_n4064_38528# a_n2302_38778# 0.239588f
C5898 a_n2946_38778# a_n2860_38778# 0.011479f
C5899 en_comp a_22589_40055# 0.260977f
C5900 a_17499_43370# a_16823_43084# 0.064861f
C5901 a_13259_45724# a_15493_43396# 0.021264f
C5902 a_19692_46634# a_743_42282# 0.150479f
C5903 a_3232_43370# a_11691_44458# 0.251483f
C5904 a_15227_44166# a_20411_46873# 0.041968f
C5905 a_n2312_38680# a_n2956_39304# 5.96956f
C5906 a_5257_43370# a_3483_46348# 0.028522f
C5907 a_2063_45854# a_6511_45714# 0.037319f
C5908 C8_P_btm C0_dummy_P_btm 0.234177f
C5909 EN_VIN_BSTR_N C5_N_btm 0.115337f
C5910 C6_P_btm C1_P_btm 0.127656f
C5911 C7_P_btm C0_P_btm 0.140846f
C5912 C4_P_btm C3_P_btm 9.61674f
C5913 C5_P_btm C2_P_btm 0.13795f
C5914 a_n2002_35448# VDD 0.522945f
C5915 a_10157_44484# VDD 0.174233f
C5916 a_13507_46334# a_13258_32519# 0.049541f
C5917 a_11827_44484# a_17517_44484# 0.05115f
C5918 a_n2433_44484# a_n2293_43922# 0.010009f
C5919 a_5883_43914# a_5891_43370# 0.216958f
C5920 a_10249_46116# a_10193_42453# 0.034764f
C5921 a_9290_44172# a_10809_44734# 0.239594f
C5922 a_3090_45724# a_2711_45572# 0.555348f
C5923 SMPL_ON_N a_413_45260# 0.199669f
C5924 a_5534_30871# a_6123_31319# 0.01835f
C5925 a_4361_42308# a_20107_42308# 0.010379f
C5926 a_n967_45348# a_n1853_43023# 0.021497f
C5927 a_3357_43084# a_1847_42826# 0.010588f
C5928 a_3537_45260# a_4361_42308# 0.017454f
C5929 a_n1059_45260# a_n13_43084# 0.027848f
C5930 a_n913_45002# a_n1076_43230# 0.05439f
C5931 a_n1899_43946# a_n1331_43914# 0.171939f
C5932 a_n2065_43946# a_n809_44244# 0.043475f
C5933 a_n1761_44111# a_n1549_44318# 0.033724f
C5934 a_18494_42460# a_3626_43646# 0.066461f
C5935 a_n755_45592# a_n2293_42282# 0.208531f
C5936 a_2324_44458# a_8696_44636# 0.033373f
C5937 a_13661_43548# a_18443_44721# 0.011774f
C5938 a_n357_42282# a_997_45618# 0.023595f
C5939 a_12861_44030# a_19615_44636# 0.094785f
C5940 a_1431_47204# a_2124_47436# 0.010942f
C5941 a_n746_45260# a_n1151_42308# 0.116939f
C5942 a_n1741_47186# a_4791_45118# 0.024211f
C5943 a_n2109_47186# a_4915_47217# 0.352259f
C5944 a_n237_47217# a_3160_47472# 0.037234f
C5945 a_685_42968# VDD 0.088446f
C5946 a_20820_30879# EN_OFFSET_CAL 0.107181f
C5947 a_11823_42460# a_11633_42558# 0.039752f
C5948 a_n2661_42834# a_n2472_42826# 0.03087f
C5949 a_n1991_46122# VDD 0.581018f
C5950 a_22959_43948# a_17538_32519# 0.168682f
C5951 a_16855_45546# a_8696_44636# 0.112262f
C5952 a_15765_45572# a_16020_45572# 0.056391f
C5953 a_16327_47482# a_2982_43646# 0.030062f
C5954 a_9290_44172# a_5883_43914# 0.026946f
C5955 a_n443_42852# a_3232_43370# 0.02112f
C5956 a_6151_47436# a_6969_46634# 0.030417f
C5957 a_6545_47178# a_6755_46942# 0.022995f
C5958 a_n881_46662# a_n1021_46688# 0.15991f
C5959 a_n1613_43370# a_n743_46660# 0.521102f
C5960 a_18504_43218# VDD 0.077608f
C5961 a_n4209_39590# a_n3420_39616# 0.234699f
C5962 a_n2302_40160# a_n2302_39866# 0.050477f
C5963 a_4958_30871# a_n4064_38528# 0.030901f
C5964 a_14579_43548# a_15095_43370# 0.109081f
C5965 a_9803_43646# a_10341_43396# 0.11445f
C5966 a_14358_43442# a_14205_43396# 0.163543f
C5967 a_7499_43078# VDD 1.87959f
C5968 a_n357_42282# a_11967_42832# 0.153035f
C5969 a_5147_45002# a_1423_45028# 0.017515f
C5970 a_7499_43078# a_7640_43914# 0.021219f
C5971 a_6171_45002# a_16751_45260# 0.104212f
C5972 a_n2017_45002# a_n2293_42834# 0.28698f
C5973 a_13507_46334# a_6945_45028# 0.187229f
C5974 a_n743_46660# a_n2293_46098# 0.213418f
C5975 a_n2438_43548# a_n2472_46090# 0.020059f
C5976 a_n1925_46634# a_n1853_46287# 0.012373f
C5977 a_11735_46660# a_11813_46116# 0.162547f
C5978 a_5807_45002# a_3483_46348# 0.018693f
C5979 a_4883_46098# a_20708_46348# 0.014516f
C5980 a_22589_40599# a_22527_39145# 1.41544f
C5981 a_22537_40625# a_22589_40055# 0.076642f
C5982 a_3422_30871# a_7174_31319# 2.22059f
C5983 a_10083_42826# a_10518_42984# 0.234322f
C5984 a_1307_43914# a_16241_44734# 0.010259f
C5985 a_n2129_44697# a_n452_44636# 0.079904f
C5986 a_n2267_44484# a_n1352_44484# 0.118759f
C5987 a_11691_44458# a_8975_43940# 0.048259f
C5988 a_413_45260# a_22959_44484# 0.202222f
C5989 a_n967_45348# a_n1899_43946# 0.025102f
C5990 a_n2661_45010# a_2127_44172# 0.096614f
C5991 a_n443_42852# a_4905_42826# 0.037419f
C5992 a_n2661_44458# a_949_44458# 0.041721f
C5993 a_13661_43548# a_13249_42308# 0.486588f
C5994 a_5807_45002# a_14495_45572# 0.012666f
C5995 a_13747_46662# a_13904_45546# 0.031534f
C5996 a_19692_46634# a_8049_45260# 0.045516f
C5997 a_20273_46660# a_10809_44734# 0.027345f
C5998 a_n237_47217# a_413_45260# 0.030002f
C5999 a_n746_45260# a_327_44734# 0.256943f
C6000 a_3483_46348# a_3699_46348# 0.06281f
C6001 a_6151_47436# a_3357_43084# 0.025786f
C6002 a_3600_43914# VDD 0.22716f
C6003 a_743_42282# a_6761_42308# 0.01018f
C6004 a_5649_42852# a_4921_42308# 0.133152f
C6005 a_4190_30871# a_6123_31319# 0.018095f
C6006 a_4361_42308# a_5755_42308# 0.010214f
C6007 a_16795_42852# a_17141_43172# 0.013377f
C6008 a_20193_45348# a_14021_43940# 0.118757f
C6009 a_n2661_43922# a_n2472_43914# 0.068474f
C6010 a_n2661_42834# a_n2065_43946# 0.035267f
C6011 a_n913_45002# a_10341_43396# 0.032712f
C6012 a_11823_42460# a_12379_42858# 0.033971f
C6013 a_10193_42453# a_5534_30871# 0.136243f
C6014 a_10903_43370# a_13291_42460# 0.135558f
C6015 a_4185_45028# a_22400_42852# 0.105559f
C6016 a_5129_47502# VDD 0.20906f
C6017 a_3785_47178# DATA[2] 0.119025f
C6018 a_12549_44172# a_11827_44484# 1.40268f
C6019 a_9625_46129# a_10053_45546# 0.086776f
C6020 a_8199_44636# a_8746_45002# 0.680077f
C6021 a_16327_47482# a_14539_43914# 0.031714f
C6022 a_2324_44458# a_7227_45028# 0.035814f
C6023 a_526_44458# a_3218_45724# 0.032949f
C6024 a_15781_43660# VDD 0.196099f
C6025 a_4190_30871# EN_VIN_BSTR_P 0.043599f
C6026 a_18079_43940# a_15493_43940# 0.040279f
C6027 a_19862_44208# a_20365_43914# 0.075162f
C6028 a_9313_44734# a_12281_43396# 0.027032f
C6029 a_n2956_39304# a_n2946_39072# 0.150476f
C6030 a_15227_44166# VDD 2.69945f
C6031 a_11322_45546# a_11682_45822# 0.034435f
C6032 a_5066_45546# a_8953_45002# 0.013782f
C6033 a_20692_30879# a_19479_31679# 0.051569f
C6034 a_21076_30879# a_18114_32519# 0.054909f
C6035 a_16023_47582# a_15928_47570# 0.049827f
C6036 a_12861_44030# a_13661_43548# 0.8566f
C6037 a_4791_45118# a_n743_46660# 0.080217f
C6038 a_10227_46804# a_11309_47204# 0.026748f
C6039 a_14021_43940# a_20301_43646# 0.024612f
C6040 en_comp a_4958_30871# 0.086457f
C6041 a_18184_42460# a_20256_43172# 0.043416f
C6042 a_3357_43084# a_5111_44636# 0.318002f
C6043 a_n745_45366# a_n467_45028# 0.110406f
C6044 a_13661_43548# a_19700_43370# 0.042923f
C6045 a_10193_42453# a_11691_44458# 0.046462f
C6046 SMPL_ON_N a_20820_30879# 0.029764f
C6047 a_n743_46660# a_16292_46812# 0.064277f
C6048 a_3877_44458# a_6755_46942# 0.388535f
C6049 a_n1741_47186# a_6945_45028# 2.51584f
C6050 a_13747_46662# a_14035_46660# 0.040628f
C6051 a_7174_31319# VDD 0.670206f
C6052 a_4958_30871# VREF_GND 0.054206f
C6053 a_3422_30871# a_5932_42308# 0.022048f
C6054 a_n2157_42858# a_n1991_42858# 0.905962f
C6055 a_4558_45348# VDD 0.25277f
C6056 a_n4318_39768# a_n4318_38216# 0.023318f
C6057 a_413_45260# DATA[5] 0.0381f
C6058 a_3537_45260# a_5891_43370# 0.359819f
C6059 a_14537_43396# a_14539_43914# 0.135541f
C6060 a_n913_45002# a_n2293_43922# 0.019153f
C6061 a_526_44458# a_6293_42852# 0.029694f
C6062 a_17719_45144# a_18315_45260# 0.017382f
C6063 a_16922_45042# a_19778_44110# 0.026041f
C6064 a_7499_43078# a_10729_43914# 0.23002f
C6065 a_21076_30879# a_13887_32519# 0.055154f
C6066 a_10227_46804# a_10490_45724# 0.031f
C6067 VREF_GND VCM 2.79113f
C6068 a_3626_43646# a_5742_30871# 0.168508f
C6069 a_n357_42282# a_10518_42984# 0.010947f
C6070 w_1575_34786# a_n1057_35014# 41.7287f
C6071 a_n1917_44484# a_n1899_43946# 0.012479f
C6072 a_18443_44721# a_11967_42832# 0.035979f
C6073 a_10193_42453# a_4190_30871# 0.305842f
C6074 a_n913_45002# a_n97_42460# 0.109647f
C6075 a_12861_44030# a_18587_45118# 0.011009f
C6076 a_n971_45724# a_n699_43396# 0.139047f
C6077 a_n2293_46634# a_5111_44636# 0.130609f
C6078 a_1756_43548# VDD 0.138878f
C6079 a_1307_43914# a_3935_42891# 0.318189f
C6080 a_n356_44636# a_2982_43646# 0.434193f
C6081 a_n2956_38216# a_n4318_38216# 0.023519f
C6082 a_n443_42852# a_10193_42453# 0.026599f
C6083 a_3483_46348# a_13017_45260# 0.51131f
C6084 a_13259_45724# a_15765_45572# 0.025388f
C6085 a_8199_44636# a_3232_43370# 0.32342f
C6086 a_5937_45572# a_5691_45260# 0.061637f
C6087 a_19692_46634# a_20193_45348# 0.060606f
C6088 a_8049_45260# a_18175_45572# 0.014402f
C6089 a_n2109_47186# a_n881_46662# 0.023562f
C6090 a_n784_42308# a_7174_31319# 1.93626f
C6091 a_11341_43940# a_9145_43396# 0.017582f
C6092 a_15493_43396# a_14955_43396# 0.076347f
C6093 a_n2267_43396# a_n1177_43370# 0.041762f
C6094 a_n1699_43638# a_n1917_43396# 0.209641f
C6095 a_n2129_43609# a_n1352_43396# 0.041828f
C6096 a_6945_45028# SINGLE_ENDED 0.021393f
C6097 a_n913_45002# a_3823_42558# 0.029622f
C6098 a_18184_42460# a_21195_42852# 0.017258f
C6099 a_22959_46124# VDD 0.309939f
C6100 a_16327_47482# a_17324_43396# 0.216094f
C6101 a_4791_45118# a_4361_42308# 0.111224f
C6102 a_n2293_46634# a_4235_43370# 0.012147f
C6103 a_7499_43078# a_1423_45028# 0.020575f
C6104 a_2107_46812# a_n2661_46098# 0.037509f
C6105 a_1983_46706# a_1799_45572# 0.089984f
C6106 a_n2661_46634# a_4651_46660# 0.020633f
C6107 a_11309_47204# a_10467_46802# 0.023291f
C6108 a_9804_47204# a_10249_46116# 0.034717f
C6109 a_8128_46384# a_6755_46942# 0.01823f
C6110 a_n2497_47436# a_n1991_46122# 0.037858f
C6111 a_11599_46634# a_14035_46660# 0.021792f
C6112 a_4883_46098# a_14976_45028# 0.019383f
C6113 a_13507_46334# a_15559_46634# 0.216791f
C6114 a_18597_46090# a_19466_46812# 0.074092f
C6115 a_10227_46804# a_12156_46660# 0.025653f
C6116 a_5934_30871# C5_N_btm 0.139996f
C6117 a_5932_42308# VDD 0.534594f
C6118 a_3080_42308# a_5534_30871# 0.019853f
C6119 a_16759_43396# a_16823_43084# 0.038761f
C6120 a_16137_43396# a_4190_30871# 0.113768f
C6121 a_20193_45348# a_21613_42308# 0.137559f
C6122 a_16327_47482# a_19987_42826# 0.053812f
C6123 a_13249_42308# a_11967_42832# 0.023012f
C6124 a_n913_45002# a_742_44458# 0.302053f
C6125 a_19692_46634# a_20301_43646# 0.110092f
C6126 a_19333_46634# a_19551_46910# 0.08213f
C6127 a_n743_46660# a_6945_45028# 0.029165f
C6128 a_2063_45854# a_6472_45840# 0.545607f
C6129 a_4646_46812# a_5937_45572# 0.105447f
C6130 C9_P_btm C0_dummy_P_btm 0.111645f
C6131 EN_VIN_BSTR_N C4_N_btm 0.116925f
C6132 C6_P_btm C2_P_btm 0.137206f
C6133 C7_P_btm C1_P_btm 0.128479f
C6134 C8_P_btm C0_P_btm 0.146541f
C6135 C5_P_btm C3_P_btm 0.135528f
C6136 a_9838_44484# VDD 0.242131f
C6137 a_n1557_42282# a_n1736_42282# 0.170341f
C6138 a_n443_42852# a_16137_43396# 0.020044f
C6139 a_n2433_44484# a_n2661_43922# 0.075698f
C6140 a_16922_45042# a_20159_44458# 0.012027f
C6141 a_742_44458# a_556_44484# 0.044092f
C6142 a_2324_44458# a_15682_46116# 0.343876f
C6143 a_4419_46090# a_n1925_42282# 0.056546f
C6144 a_10227_46804# a_6171_45002# 0.087616f
C6145 a_4361_42308# a_13258_32519# 0.076336f
C6146 a_n967_45348# a_n2157_42858# 0.02564f
C6147 a_5111_44636# a_743_42282# 0.024053f
C6148 a_n913_45002# a_n901_43156# 0.075029f
C6149 a_n2065_43946# a_n1549_44318# 0.110816f
C6150 a_n1761_44111# a_n1331_43914# 0.043168f
C6151 a_18184_42460# a_3626_43646# 0.052679f
C6152 a_n881_46662# RST_Z 0.351994f
C6153 a_n357_42282# a_n2293_42282# 0.01064f
C6154 a_n1613_43370# a_5891_43370# 0.064769f
C6155 a_15682_46116# a_16855_45546# 0.011741f
C6156 a_13661_43548# a_18287_44626# 0.021421f
C6157 a_n357_42282# a_n755_45592# 0.664842f
C6158 a_10227_46804# a_14673_44172# 0.012944f
C6159 a_12861_44030# a_11967_42832# 0.209245f
C6160 a_n971_45724# a_n1151_42308# 0.682801f
C6161 a_1209_47178# a_584_46384# 0.104123f
C6162 a_n237_47217# a_2905_45572# 0.025329f
C6163 a_n2109_47186# a_n443_46116# 0.080373f
C6164 COMP_P a_6123_31319# 0.028802f
C6165 a_n784_42308# a_5932_42308# 0.151611f
C6166 a_n913_45002# a_12800_43218# 0.016338f
C6167 a_n2661_42834# a_n2840_42826# 0.174935f
C6168 a_22591_46660# EN_OFFSET_CAL 0.047938f
C6169 a_11823_42460# a_11551_42558# 0.138126f
C6170 a_n1853_46287# VDD 0.645231f
C6171 a_15493_43940# a_17538_32519# 0.013565f
C6172 a_16855_45546# a_16680_45572# 0.233657f
C6173 a_15903_45785# a_16020_45572# 0.157972f
C6174 a_8199_44636# a_8975_43940# 0.028334f
C6175 a_6151_47436# a_6755_46942# 0.361724f
C6176 a_n881_46662# a_n1925_46634# 0.467945f
C6177 a_n4209_39590# a_n3690_39616# 0.045251f
C6178 a_3080_42308# a_4190_30871# 0.01835f
C6179 a_9803_43646# a_9885_43646# 0.171361f
C6180 a_9145_43396# a_10341_43396# 0.085699f
C6181 a_14579_43548# a_14205_43396# 0.066243f
C6182 a_742_44458# a_1755_42282# 0.013027f
C6183 a_8568_45546# VDD 0.182812f
C6184 a_18479_45785# a_11691_44458# 0.025645f
C6185 a_6171_45002# a_1307_43914# 0.037515f
C6186 a_21076_30879# a_14401_32519# 0.057698f
C6187 CAL_N a_22527_39145# 0.010004f
C6188 a_22589_40599# a_22589_40055# 0.086408f
C6189 a_n4064_38528# VREF_GND 0.034351f
C6190 a_n3565_37414# EN_VIN_BSTR_P 0.095737f
C6191 a_3422_30871# a_20712_42282# 0.016384f
C6192 a_n2661_43370# VDD 1.53673f
C6193 a_1307_43914# a_14673_44172# 0.012594f
C6194 a_n913_45002# a_n984_44318# 0.013973f
C6195 a_n2267_44484# a_n1177_44458# 0.042415f
C6196 a_n1699_44726# a_n1917_44484# 0.209641f
C6197 a_n2129_44697# a_n1352_44484# 0.048248f
C6198 a_n2661_44458# a_742_44458# 0.026794f
C6199 a_413_45260# a_17730_32519# 0.026007f
C6200 a_n967_45348# a_n1761_44111# 0.015839f
C6201 a_n443_42852# a_3080_42308# 0.029846f
C6202 a_3357_43084# a_3905_42865# 0.125186f
C6203 a_5807_45002# a_13249_42308# 0.725941f
C6204 a_19466_46812# a_8049_45260# 0.061209f
C6205 a_20841_46902# a_6945_45028# 0.013693f
C6206 a_20411_46873# a_10809_44734# 0.010692f
C6207 a_n746_45260# a_413_45260# 0.031693f
C6208 a_n1151_42308# a_n2293_45010# 0.020357f
C6209 a_n1925_46634# a_8162_45546# 0.104508f
C6210 a_n2661_46634# a_10193_42453# 0.351509f
C6211 a_4646_46812# a_n443_42852# 0.038263f
C6212 a_16327_47482# a_18799_45938# 0.013823f
C6213 a_5815_47464# a_3357_43084# 0.029103f
C6214 a_2998_44172# VDD 0.362233f
C6215 a_n2661_42834# a_n2472_43914# 0.012267f
C6216 a_n1059_45260# a_10341_43396# 0.037338f
C6217 a_18479_45785# a_4190_30871# 0.123942f
C6218 a_17517_44484# a_19279_43940# 0.020718f
C6219 a_n2661_43922# a_n2840_43914# 0.171265f
C6220 a_4915_47217# VDD 3.43172f
C6221 a_12891_46348# a_11827_44484# 0.020579f
C6222 a_8199_44636# a_10193_42453# 0.236934f
C6223 a_18285_46348# a_18175_45572# 0.010439f
C6224 a_8049_45260# a_20205_31679# 0.301209f
C6225 a_11415_45002# a_15903_45785# 0.02962f
C6226 a_12861_44030# a_18989_43940# 0.047422f
C6227 a_4791_45118# a_5891_43370# 0.066388f
C6228 a_15681_43442# VDD 0.159054f
C6229 a_4190_30871# a_n1057_35014# 0.027898f
C6230 a_19862_44208# a_20269_44172# 0.049487f
C6231 a_n2293_43922# a_9145_43396# 0.019866f
C6232 a_17973_43940# a_15493_43940# 0.028173f
C6233 a_n2956_39304# a_n3420_39072# 0.208204f
C6234 a_18834_46812# VDD 0.116625f
C6235 a_13259_45724# a_n913_45002# 0.142601f
C6236 a_20205_31679# a_19479_31679# 0.06173f
C6237 a_10490_45724# a_11682_45822# 0.014138f
C6238 a_n2293_46634# a_3905_42865# 0.039006f
C6239 a_n443_46116# a_n1925_46634# 0.080855f
C6240 a_6491_46660# a_n2661_46634# 0.013828f
C6241 a_12861_44030# a_5807_45002# 0.214011f
C6242 a_n3674_37592# a_n4064_37984# 0.020548f
C6243 a_20447_31679# a_13258_32519# 0.054935f
C6244 a_14021_43940# a_4190_30871# 0.086029f
C6245 a_n1059_45260# a_18727_42674# 0.20226f
C6246 a_n443_42852# a_10057_43914# 0.06562f
C6247 a_13661_43548# a_19268_43646# 0.136251f
C6248 a_3357_43084# a_5147_45002# 0.09352f
C6249 a_11453_44696# a_11415_45002# 0.123733f
C6250 SMPL_ON_N a_22591_46660# 0.011048f
C6251 a_13747_46662# a_13885_46660# 0.028801f
C6252 a_n4064_39616# C9_P_btm 0.215899f
C6253 a_7754_39964# a_7754_38470# 0.241119f
C6254 a_20712_42282# VDD 0.282526f
C6255 a_3754_39134# a_3754_38802# 0.296258f
C6256 a_n2157_42858# a_n1853_43023# 0.290902f
C6257 a_n3674_39768# a_n3674_38680# 0.035445f
C6258 a_4574_45260# VDD 0.122256f
C6259 a_1414_42308# a_1184_42692# 0.115223f
C6260 a_413_45260# DATA[4] 0.037695f
C6261 a_3537_45260# a_8375_44464# 0.10437f
C6262 a_1423_45028# a_9838_44484# 0.254741f
C6263 a_14537_43396# a_16112_44458# 0.093722f
C6264 a_20820_30879# a_14209_32519# 0.053104f
C6265 a_n913_45002# a_n2661_43922# 0.024256f
C6266 a_n1059_45260# a_n2293_43922# 0.02309f
C6267 a_16922_45042# a_18911_45144# 0.042178f
C6268 a_15227_44166# a_15567_42826# 0.075768f
C6269 a_n443_42852# a_14021_43940# 0.05804f
C6270 a_7499_43078# a_10405_44172# 0.132405f
C6271 a_n1613_43370# a_8292_43218# 0.011565f
C6272 a_10227_46804# a_8746_45002# 0.117547f
C6273 a_3090_45724# a_10903_43370# 0.031245f
C6274 VREF VCM 44.262398f
C6275 a_n357_42282# a_10083_42826# 0.017324f
C6276 a_3357_43084# a_4093_43548# 0.031759f
C6277 w_1575_34786# a_n1696_34930# 0.799379f
C6278 a_18287_44626# a_11967_42832# 0.789765f
C6279 a_18374_44850# a_18588_44850# 0.097745f
C6280 a_18443_44721# a_19006_44850# 0.049827f
C6281 a_n1059_45260# a_n97_42460# 0.869353f
C6282 a_14275_46494# a_14383_46116# 0.057222f
C6283 a_1823_45246# a_3503_45724# 0.295715f
C6284 a_1568_43370# VDD 0.433732f
C6285 a_22959_42860# a_14097_32519# 0.166017f
C6286 a_n2661_42834# a_n2433_43396# 0.02044f
C6287 a_1307_43914# a_3681_42891# 0.236785f
C6288 a_n2810_45572# a_n3674_38216# 0.023322f
C6289 a_8953_45546# a_5111_44636# 0.181796f
C6290 a_2107_46812# a_n2661_43922# 0.027806f
C6291 a_12549_44172# a_19279_43940# 0.062614f
C6292 a_3483_46348# a_11963_45334# 0.016005f
C6293 a_13259_45724# a_15903_45785# 0.064252f
C6294 a_8016_46348# a_6171_45002# 0.022961f
C6295 a_6511_45714# a_7227_45028# 0.213161f
C6296 a_6667_45809# a_6598_45938# 0.209641f
C6297 a_n1151_42308# a_12465_44636# 0.02014f
C6298 a_n2109_47186# a_n1613_43370# 0.054203f
C6299 a_12861_44030# a_14311_47204# 0.037394f
C6300 a_n1761_44111# a_n1853_43023# 0.019636f
C6301 a_n2267_43396# a_n1917_43396# 0.227165f
C6302 a_n2129_43609# a_n1177_43370# 0.08445f
C6303 a_6945_45028# START 0.029602f
C6304 a_n2433_43396# a_n1352_43396# 0.102325f
C6305 a_n913_45002# a_3318_42354# 0.03912f
C6306 a_18184_42460# a_21356_42826# 0.016504f
C6307 a_10809_44734# VDD 2.67671f
C6308 a_16327_47482# a_17499_43370# 0.34052f
C6309 a_20820_30879# a_17730_32519# 0.052913f
C6310 a_3090_45724# a_14955_43940# 0.018423f
C6311 a_10193_42453# a_16751_45260# 0.048213f
C6312 a_2107_46812# a_1799_45572# 0.079386f
C6313 a_948_46660# a_n2661_46098# 0.018472f
C6314 a_n2661_46634# a_4646_46812# 0.087334f
C6315 a_11309_47204# a_10428_46928# 0.025525f
C6316 a_n2497_47436# a_n1853_46287# 0.029452f
C6317 a_6491_46660# a_765_45546# 0.042766f
C6318 a_18479_47436# a_19692_46634# 0.078022f
C6319 a_13507_46334# a_15368_46634# 0.023781f
C6320 a_4883_46098# a_3090_45724# 0.052016f
C6321 a_n2946_38778# a_n4064_38528# 0.053228f
C6322 a_5934_30871# C4_N_btm 0.030578f
C6323 a_6171_42473# VDD 0.184622f
C6324 a_16977_43638# a_16823_43084# 0.022663f
C6325 a_n2293_43922# a_1606_42308# 0.080878f
C6326 a_20193_45348# a_21887_42336# 0.169001f
C6327 en_comp a_22537_40625# 0.021487f
C6328 a_16327_47482# a_19164_43230# 0.292734f
C6329 a_1423_45028# a_n2661_43370# 0.027675f
C6330 a_413_45260# a_19721_31679# 0.116395f
C6331 a_14180_45002# a_14309_45028# 0.062574f
C6332 a_n467_45028# a_n2661_44458# 0.031118f
C6333 a_n1059_45260# a_742_44458# 0.030569f
C6334 a_19692_46634# a_4190_30871# 0.013919f
C6335 a_19333_46634# a_19123_46287# 0.113955f
C6336 a_15227_44166# a_19551_46910# 0.018691f
C6337 a_11453_44696# a_13259_45724# 0.251534f
C6338 a_2063_45854# a_6194_45824# 0.041827f
C6339 a_n2442_46660# a_n2956_38680# 0.047296f
C6340 a_n1151_42308# a_2711_45572# 0.039506f
C6341 C10_P_btm C0_dummy_P_btm 0.749362f
C6342 EN_VIN_BSTR_N C3_N_btm 0.100325f
C6343 C6_P_btm C3_P_btm 0.133742f
C6344 C7_P_btm C2_P_btm 0.138288f
C6345 C5_P_btm C4_P_btm 18.6196f
C6346 C9_P_btm C0_P_btm 0.146135f
C6347 C8_P_btm C1_P_btm 0.129306f
C6348 a_5883_43914# VDD 0.859221f
C6349 a_3080_42308# COMP_P 4.43537f
C6350 a_8103_44636# a_5891_43370# 0.029956f
C6351 a_1307_43914# a_5663_43940# 0.11718f
C6352 a_n2661_44458# a_n2661_43922# 6.64988f
C6353 a_18287_44626# a_18989_43940# 0.193279f
C6354 a_18443_44721# a_18374_44850# 0.209641f
C6355 a_4419_46090# a_526_44458# 0.099848f
C6356 a_4185_45028# a_n1925_42282# 0.638728f
C6357 a_12861_44030# a_13017_45260# 0.032265f
C6358 a_n2497_47436# a_n2661_43370# 0.031125f
C6359 a_n971_45724# a_n2293_42834# 0.088674f
C6360 a_10227_46804# a_3232_43370# 0.028168f
C6361 a_13467_32519# a_13258_32519# 11.0084f
C6362 a_n1059_45260# a_n901_43156# 0.021049f
C6363 a_n881_46662# VDD 2.6692f
C6364 a_n1761_44111# a_n1899_43946# 0.737653f
C6365 a_n2065_43946# a_n1331_43914# 0.053479f
C6366 a_310_45028# a_n755_45592# 0.02846f
C6367 a_20202_43084# a_n913_45002# 0.322116f
C6368 a_13661_43548# a_18248_44752# 0.019034f
C6369 a_1239_47204# a_1431_47204# 0.219138f
C6370 a_n971_45724# a_3160_47472# 0.011577f
C6371 a_1209_47178# a_2124_47436# 0.095065f
C6372 a_n1741_47186# a_4007_47204# 0.012359f
C6373 a_n2109_47186# a_4791_45118# 0.34446f
C6374 a_7845_44172# a_7287_43370# 0.011834f
C6375 a_15493_43940# a_20974_43370# 0.069596f
C6376 a_3499_42826# a_2982_43646# 0.018486f
C6377 a_11415_45002# EN_OFFSET_CAL 0.14622f
C6378 a_n2157_46122# VDD 0.42567f
C6379 a_3175_45822# a_413_45260# 0.011644f
C6380 a_1138_42852# a_n356_44636# 0.29814f
C6381 a_15599_45572# a_16020_45572# 0.086708f
C6382 a_8199_44636# a_10057_43914# 0.113262f
C6383 a_6151_47436# a_10249_46116# 0.056387f
C6384 a_n1613_43370# a_n1925_46634# 0.33524f
C6385 a_9804_47204# a_n2661_46634# 0.02862f
C6386 a_n4064_40160# a_n4064_39616# 5.80519f
C6387 a_n4209_39590# a_n3565_39590# 6.15218f
C6388 a_4958_30871# a_n3420_38528# 0.030871f
C6389 a_n2956_37592# a_n4064_38528# 0.015398f
C6390 a_8162_45546# VDD 0.266272f
C6391 a_9145_43396# a_9885_43646# 0.052876f
C6392 a_13667_43396# a_14205_43396# 0.076384f
C6393 a_14579_43548# a_14358_43442# 0.142377f
C6394 a_8953_45002# a_9482_43914# 0.010057f
C6395 a_2680_45002# a_2903_45348# 0.011458f
C6396 a_18479_45785# a_19113_45348# 0.013845f
C6397 a_3232_43370# a_1307_43914# 0.14252f
C6398 a_6171_45002# a_16019_45002# 0.01229f
C6399 a_20820_30879# a_17538_32519# 0.052874f
C6400 a_3090_45724# a_8685_43396# 2.11639f
C6401 a_11453_44696# a_18189_46348# 0.534507f
C6402 a_20990_47178# a_6945_45028# 0.026188f
C6403 a_n1925_46634# a_n2293_46098# 0.077794f
C6404 a_n2293_46634# a_n1991_46122# 0.0181f
C6405 a_4883_46098# a_20075_46420# 0.014562f
C6406 a_9313_45822# a_5066_45546# 0.019449f
C6407 a_n2302_37984# VDD 0.350854f
C6408 a_3726_37500# CAL_P 0.102027f
C6409 a_n2433_44484# a_n1352_44484# 0.102355f
C6410 a_n2661_45010# a_1414_42308# 0.059385f
C6411 a_n2293_45010# a_1115_44172# 0.09282f
C6412 a_n2267_44484# a_n1917_44484# 0.212549f
C6413 a_n2129_44697# a_n1177_44458# 0.027646f
C6414 a_13259_45724# a_9145_43396# 0.155949f
C6415 a_413_45260# a_22591_44484# 0.024147f
C6416 a_n967_45348# a_n2065_43946# 0.02253f
C6417 a_6545_47178# a_2437_43646# 0.010642f
C6418 a_20273_46660# a_6945_45028# 0.02808f
C6419 a_20107_46660# a_10809_44734# 0.026612f
C6420 a_n971_45724# a_413_45260# 0.937818f
C6421 a_n746_45260# a_n37_45144# 0.031257f
C6422 a_3147_46376# a_3483_46348# 0.207919f
C6423 a_n2293_46634# a_7499_43078# 0.14773f
C6424 a_2889_44172# VDD 0.1447f
C6425 a_17517_44484# a_20766_44850# 0.018462f
C6426 a_n2661_42834# a_n2840_43914# 0.014735f
C6427 a_n443_46116# VDD 3.87014f
C6428 a_2063_45854# CLK 0.271193f
C6429 a_n1151_42308# DATA[2] 0.01294f
C6430 a_19692_46634# a_2437_43646# 0.293918f
C6431 a_15227_44166# a_3357_43084# 0.026794f
C6432 a_13661_43548# a_16922_45042# 0.080391f
C6433 a_3483_46348# a_13249_42308# 0.338396f
C6434 a_8199_44636# a_10180_45724# 0.216999f
C6435 a_8016_46348# a_8746_45002# 0.078716f
C6436 a_10227_46804# a_8975_43940# 0.037352f
C6437 a_8953_45546# a_9049_44484# 0.03092f
C6438 a_17339_46660# a_18341_45572# 0.015732f
C6439 a_4791_45118# a_8375_44464# 0.010645f
C6440 a_17737_43940# a_15493_43940# 0.037029f
C6441 a_10807_43548# a_11173_44260# 0.05223f
C6442 a_n2956_39304# a_n3690_39392# 0.016795f
C6443 a_n2956_38680# a_n3565_39304# 0.068534f
C6444 a_17609_46634# VDD 0.501057f
C6445 a_11322_45546# a_10907_45822# 0.012408f
C6446 a_20820_30879# a_19721_31679# 0.052985f
C6447 a_13249_42308# a_14495_45572# 0.027073f
C6448 a_13259_45724# a_n1059_45260# 0.390886f
C6449 a_584_46384# a_1983_46706# 0.062968f
C6450 a_2063_45854# a_2107_46812# 0.214026f
C6451 a_4791_45118# a_n1925_46634# 0.026798f
C6452 a_6545_47178# a_n2661_46634# 0.022455f
C6453 a_n237_47217# a_n2661_46098# 0.01906f
C6454 a_14021_43940# a_21259_43561# 0.021338f
C6455 a_19443_46116# VDD 0.132317f
C6456 a_n1059_45260# a_18057_42282# 0.141112f
C6457 a_n2956_37592# en_comp 0.013325f
C6458 a_13661_43548# a_15743_43084# 0.092364f
C6459 a_4646_46812# a_6452_43396# 0.013786f
C6460 a_n1059_45260# a_n467_45028# 0.229142f
C6461 a_n743_46660# a_15368_46634# 0.026392f
C6462 a_9804_47204# a_765_45546# 0.028432f
C6463 a_22731_47423# a_22591_46660# 0.011433f
C6464 a_12465_44636# a_12741_44636# 0.914049f
C6465 a_12861_44030# a_3483_46348# 0.06952f
C6466 a_5807_45002# a_14035_46660# 0.025174f
C6467 a_n3420_39616# C8_P_btm 0.090298f
C6468 a_13258_32519# RST_Z 0.059325f
C6469 a_7754_40130# a_8530_39574# 0.013981f
C6470 VDAC_Pi a_3754_38470# 0.389564f
C6471 a_n2302_37984# a_n2302_37690# 0.050477f
C6472 a_4958_30871# VIN_N 0.025339f
C6473 a_20107_42308# VDD 0.284252f
C6474 a_n4318_39768# a_n3674_38680# 0.027425f
C6475 a_413_45260# DATA[3] 0.037695f
C6476 a_3537_45260# VDD 3.9063f
C6477 a_2711_45572# a_15493_43940# 0.128282f
C6478 a_1423_45028# a_5883_43914# 0.067915f
C6479 a_4185_45028# a_15743_43084# 0.061074f
C6480 a_14537_43396# a_15004_44636# 0.047224f
C6481 a_n1059_45260# a_n2661_43922# 0.034597f
C6482 a_n913_45002# a_n2661_42834# 0.027216f
C6483 a_n2017_45002# a_n2293_43922# 0.654835f
C6484 a_17613_45144# a_17719_45144# 0.080654f
C6485 a_16922_45042# a_18587_45118# 0.021516f
C6486 a_15227_44166# a_5342_30871# 0.01169f
C6487 a_20528_46660# a_12741_44636# 0.018376f
C6488 a_10227_46804# a_10193_42453# 0.039217f
C6489 VREF VREF_GND 44.051197f
C6490 VIN_N VCM 1.7189f
C6491 a_2982_43646# a_5742_30871# 0.196805f
C6492 a_4361_42308# a_14635_42282# 0.018479f
C6493 a_n357_42282# a_8952_43230# 0.011989f
C6494 a_n967_45348# a_n2129_43609# 0.021282f
C6495 en_comp a_n2267_43396# 0.028399f
C6496 a_7499_43078# a_743_42282# 0.087933f
C6497 a_n1059_45260# a_n447_43370# 0.018401f
C6498 a_n2017_45002# a_n97_42460# 0.169401f
C6499 a_18443_44721# a_18588_44850# 0.057222f
C6500 a_18287_44626# a_19006_44850# 0.086658f
C6501 a_18248_44752# a_11967_42832# 0.500539f
C6502 a_14493_46090# a_14383_46116# 0.097745f
C6503 a_12741_44636# a_2711_45572# 0.044854f
C6504 a_17339_46660# a_10193_42453# 0.023481f
C6505 a_2063_45854# a_n2661_44458# 0.029811f
C6506 a_13059_46348# a_11823_42460# 0.256727f
C6507 a_1823_45246# a_3316_45546# 0.099099f
C6508 a_1049_43396# VDD 0.196328f
C6509 a_5342_30871# a_7174_31319# 0.046616f
C6510 a_n2661_42834# a_n4318_39304# 0.041301f
C6511 a_22485_44484# a_15493_43940# 0.087012f
C6512 a_n2956_38216# a_n3674_38680# 0.022975f
C6513 a_5937_45572# a_5111_44636# 0.06133f
C6514 a_2107_46812# a_n2661_42834# 0.028012f
C6515 a_3483_46348# a_11787_45002# 0.019413f
C6516 a_13259_45724# a_15599_45572# 0.205417f
C6517 a_8016_46348# a_3232_43370# 0.025981f
C6518 a_n357_42282# a_13249_42308# 0.024753f
C6519 a_6511_45714# a_6598_45938# 0.06628f
C6520 a_6472_45840# a_7227_45028# 0.208286f
C6521 a_12861_44030# a_13487_47204# 0.127147f
C6522 a_n2267_43396# a_n1699_43638# 0.179796f
C6523 a_n2129_43609# a_n1917_43396# 0.036131f
C6524 a_n2433_43396# a_n1177_43370# 0.043475f
C6525 a_6945_45028# RST_Z 0.022027f
C6526 a_n913_45002# a_2903_42308# 0.041908f
C6527 a_22223_46124# VDD 0.300745f
C6528 a_18184_42460# a_20922_43172# 0.018236f
C6529 a_18494_42460# a_19987_42826# 0.098055f
C6530 a_16327_47482# a_16759_43396# 0.152273f
C6531 a_10193_42453# a_1307_43914# 0.054328f
C6532 a_1123_46634# a_n2661_46098# 0.041919f
C6533 a_n2661_46634# a_3877_44458# 0.010452f
C6534 a_6545_47178# a_765_45546# 0.035873f
C6535 a_13507_46334# a_14976_45028# 0.020647f
C6536 a_18597_46090# a_15227_44166# 0.150202f
C6537 a_n2497_47436# a_n2157_46122# 0.034181f
C6538 a_12861_44030# a_14513_46634# 0.036912f
C6539 a_n3420_38528# a_n4064_38528# 8.203589f
C6540 a_n4064_39072# a_n4064_37984# 0.044699f
C6541 a_2112_39137# a_2684_37794# 0.091415f
C6542 a_5934_30871# C3_N_btm 0.011274f
C6543 a_5755_42308# VDD 0.229304f
C6544 a_6123_31319# C5_N_btm 0.022099f
C6545 a_4958_30871# CAL_N 0.039702f
C6546 en_comp a_22589_40599# 0.021612f
C6547 a_16409_43396# a_16823_43084# 0.020816f
C6548 a_16759_43396# a_16855_43396# 0.013793f
C6549 a_6171_45002# a_11827_44484# 0.09294f
C6550 a_413_45260# a_18114_32519# 0.053981f
C6551 a_10193_42453# a_18579_44172# 0.12582f
C6552 a_4185_45028# a_3539_42460# 0.065262f
C6553 en_comp a_n2267_44484# 0.029536f
C6554 a_n967_45348# a_n2129_44697# 0.017689f
C6555 a_n1059_45260# a_n452_44636# 0.010366f
C6556 a_19692_46634# a_21259_43561# 0.014184f
C6557 a_16327_47482# a_19339_43156# 0.346029f
C6558 a_15227_44166# a_19123_46287# 0.069758f
C6559 a_14180_46812# a_14513_46634# 0.253235f
C6560 a_2063_45854# a_5907_45546# 0.023999f
C6561 a_n1925_46634# a_6945_45028# 0.028603f
C6562 a_2905_45572# a_3175_45822# 0.046585f
C6563 a_n2442_46660# a_n2956_39304# 0.046604f
C6564 EN_VIN_BSTR_N C2_N_btm 0.118072f
C6565 C6_P_btm C4_P_btm 0.143514f
C6566 C7_P_btm C3_P_btm 0.134911f
C6567 C10_P_btm C0_P_btm 0.365593f
C6568 C9_P_btm C1_P_btm 0.132506f
C6569 C8_P_btm C2_P_btm 0.138777f
C6570 a_22725_37990# VDD 0.085163f
C6571 a_8701_44490# VDD 0.164475f
C6572 a_3422_30871# a_n4064_37984# 0.031408f
C6573 a_8103_44636# a_8375_44464# 0.13675f
C6574 a_1307_43914# a_5495_43940# 0.024105f
C6575 a_16922_45042# a_11967_42832# 0.019919f
C6576 a_11827_44484# a_14673_44172# 0.150125f
C6577 a_5111_44636# a_8333_44056# 0.280148f
C6578 a_18287_44626# a_18374_44850# 0.053385f
C6579 a_18248_44752# a_18989_43940# 0.207562f
C6580 a_5883_43914# a_6109_44484# 0.078113f
C6581 a_4185_45028# a_526_44458# 0.162857f
C6582 a_3699_46348# a_n1925_42282# 0.011511f
C6583 a_12465_44636# a_413_45260# 0.28925f
C6584 a_n443_46116# a_1423_45028# 0.022652f
C6585 a_5342_30871# a_5932_42308# 0.01856f
C6586 a_4361_42308# a_19511_42282# 0.071032f
C6587 en_comp a_n2472_42826# 0.019667f
C6588 a_18184_42460# a_2982_43646# 0.020575f
C6589 a_5891_43370# a_10555_44260# 0.015358f
C6590 a_n1613_43370# VDD 4.75085f
C6591 a_n2065_43946# a_n1899_43946# 0.614122f
C6592 a_n1099_45572# a_n755_45592# 0.193775f
C6593 a_310_45028# a_n357_42282# 0.113929f
C6594 a_380_45546# a_997_45618# 0.070624f
C6595 a_15682_46116# a_16333_45814# 0.011944f
C6596 a_n746_45260# a_175_44278# 0.159759f
C6597 a_16327_47482# a_17517_44484# 0.090308f
C6598 a_768_44030# a_n356_44636# 0.098499f
C6599 a_n2497_47436# a_n443_46116# 0.026321f
C6600 a_n971_45724# a_2905_45572# 0.118495f
C6601 a_n815_47178# a_n1151_42308# 0.011772f
C6602 a_1209_47178# a_1431_47204# 0.095209f
C6603 a_n1741_47186# a_3815_47204# 0.023296f
C6604 a_n2109_47186# a_4700_47436# 0.038955f
C6605 a_n1533_42852# VDD 0.142813f
C6606 a_15493_43940# a_14401_32519# 0.052433f
C6607 a_11967_42832# a_15743_43084# 0.180938f
C6608 a_n913_45002# a_11554_42852# 0.016237f
C6609 a_n2293_46098# VDD 1.7963f
C6610 a_2711_45572# a_413_45260# 0.022324f
C6611 a_16333_45814# a_16680_45572# 0.051162f
C6612 a_n443_42852# a_5111_44636# 0.584506f
C6613 a_15903_45785# a_15861_45028# 0.232345f
C6614 a_8016_46348# a_8975_43940# 0.01976f
C6615 a_8128_46384# a_n2661_46634# 0.029397f
C6616 a_n1794_35082# CAL_P 0.016411f
C6617 a_n4209_39590# a_n4334_39616# 0.25243f
C6618 a_9145_43396# a_14955_43396# 0.06858f
C6619 a_8685_43396# a_12281_43396# 0.038443f
C6620 a_7230_45938# VDD 0.077608f
C6621 a_2680_45002# a_2809_45348# 0.010132f
C6622 a_3357_43084# a_n2661_43370# 0.030835f
C6623 a_11787_45002# a_11963_45334# 0.185422f
C6624 a_6171_45002# a_15595_45028# 0.012742f
C6625 a_3537_45260# a_1423_45028# 0.046355f
C6626 a_n2104_46634# a_n2157_46122# 0.013135f
C6627 a_11453_44696# a_17715_44484# 0.036977f
C6628 a_20894_47436# a_6945_45028# 0.016564f
C6629 a_6755_46942# a_15227_44166# 0.288173f
C6630 a_n2293_46634# a_n1853_46287# 0.014216f
C6631 a_22589_40599# a_22537_40625# 1.96968f
C6632 a_n3420_38528# VREF_GND 0.047244f
C6633 a_n4064_37984# VDD 1.70643f
C6634 a_9127_43156# a_10083_42826# 0.011187f
C6635 a_3422_30871# a_13258_32519# 0.410904f
C6636 a_n2433_44484# a_n1177_44458# 0.043567f
C6637 a_n1059_45260# a_n809_44244# 0.021842f
C6638 a_n2293_45010# a_644_44056# 0.014621f
C6639 a_n443_42852# a_4235_43370# 0.026532f
C6640 a_3357_43084# a_2998_44172# 0.119142f
C6641 a_n2267_44484# a_n1699_44726# 0.172319f
C6642 a_n2129_44697# a_n1917_44484# 0.030172f
C6643 a_11827_44484# a_12607_44458# 0.023193f
C6644 a_11453_44696# a_15861_45028# 0.044605f
C6645 a_6151_47436# a_2437_43646# 0.017593f
C6646 a_n746_45260# a_n143_45144# 0.043399f
C6647 a_n1151_42308# a_n2661_45010# 0.155007f
C6648 a_15227_44166# a_8049_45260# 0.036339f
C6649 a_16327_47482# a_19256_45572# 0.235006f
C6650 a_4915_47217# a_3357_43084# 0.028255f
C6651 a_2675_43914# VDD 0.200923f
C6652 a_4361_42308# a_4921_42308# 0.472085f
C6653 a_743_42282# a_5932_42308# 0.024532f
C6654 a_17517_44484# a_20835_44721# 0.029603f
C6655 a_1307_43914# a_3080_42308# 0.01819f
C6656 a_4791_45118# VDD 3.05095f
C6657 a_n1925_42282# a_n2293_42282# 0.234055f
C6658 a_19692_46634# a_21513_45002# 0.098725f
C6659 a_n2293_46634# a_n2661_43370# 2.59564f
C6660 a_5807_45002# a_16922_45042# 0.030945f
C6661 a_8016_46348# a_10193_42453# 0.125497f
C6662 a_8199_44636# a_10053_45546# 0.014322f
C6663 a_3483_46348# a_13904_45546# 0.125708f
C6664 a_4791_45118# a_7640_43914# 0.027432f
C6665 a_10227_46804# a_10057_43914# 0.054198f
C6666 a_n1925_42282# a_n755_45592# 0.020368f
C6667 a_4646_46812# a_1307_43914# 0.031289f
C6668 a_5937_45572# a_9049_44484# 0.311862f
C6669 a_8953_45546# a_7499_43078# 0.108436f
C6670 a_17339_46660# a_18479_45785# 0.027772f
C6671 a_15682_43940# a_15493_43940# 0.067033f
C6672 a_16292_46812# VDD 0.123916f
C6673 a_n2956_39304# a_n3565_39304# 0.307358f
C6674 a_13259_45724# a_n2017_45002# 0.065062f
C6675 a_10227_46804# a_14021_43940# 0.062062f
C6676 a_13059_46348# a_14539_43914# 0.05997f
C6677 a_n2293_46634# a_2998_44172# 0.06774f
C6678 a_8568_45546# a_9159_45572# 0.011449f
C6679 a_20820_30879# a_18114_32519# 0.053f
C6680 a_13904_45546# a_14495_45572# 0.092344f
C6681 a_10193_42453# a_11682_45822# 0.032292f
C6682 a_10490_45724# a_10907_45822# 0.229517f
C6683 a_8270_45546# a_n2661_43922# 0.025118f
C6684 a_n971_45724# a_104_43370# 0.156156f
C6685 a_n237_47217# a_1799_45572# 0.417887f
C6686 a_n746_45260# a_n2661_46098# 0.049386f
C6687 a_16327_47482# a_12549_44172# 0.123271f
C6688 a_6151_47436# a_n2661_46634# 0.140541f
C6689 a_15673_47210# a_15928_47570# 0.064178f
C6690 a_n3674_37592# a_n3420_37984# 0.172946f
C6691 a_17124_42282# a_17303_42282# 0.172579f
C6692 a_20692_30879# C6_N_btm 0.080378f
C6693 a_n913_45002# a_17303_42282# 1.81467f
C6694 a_19963_31679# a_13258_32519# 0.054679f
C6695 a_13661_43548# a_18783_43370# 0.057336f
C6696 a_n745_45366# a_n967_45348# 0.010748f
C6697 a_17339_46660# a_14021_43940# 0.037923f
C6698 a_n2661_45010# a_327_44734# 0.04375f
C6699 a_15227_44166# a_15037_43940# 0.010516f
C6700 a_8128_46384# a_765_45546# 0.03129f
C6701 a_n743_46660# a_14976_45028# 0.024461f
C6702 a_5807_45002# a_13885_46660# 0.014137f
C6703 a_4958_30871# VIN_P 0.025339f
C6704 a_7754_40130# a_7754_38470# 0.112286f
C6705 a_7754_39964# a_3754_38470# 0.081868f
C6706 a_7754_39300# a_7754_38968# 0.296258f
C6707 a_13258_32519# VDD 3.19378f
C6708 a_n2472_42826# a_n2157_42858# 0.080495f
C6709 a_3429_45260# VDD 0.142923f
C6710 a_413_45260# DATA[2] 0.048779f
C6711 a_1414_42308# a_1067_42314# 0.100434f
C6712 a_1423_45028# a_8701_44490# 0.063232f
C6713 a_20820_30879# a_13887_32519# 0.053104f
C6714 a_n2017_45002# a_n2661_43922# 0.034672f
C6715 a_n1059_45260# a_n2661_42834# 0.029616f
C6716 a_526_44458# a_648_43396# 0.04105f
C6717 a_16922_45042# a_18315_45260# 0.065907f
C6718 a_18479_45785# a_18579_44172# 0.045071f
C6719 a_21076_30879# a_13678_32519# 0.05537f
C6720 a_13556_45296# a_14539_43914# 0.025347f
C6721 a_1307_43914# a_10057_43914# 0.03199f
C6722 a_22000_46634# a_12741_44636# 0.044691f
C6723 a_12991_46634# a_13351_46090# 0.011685f
C6724 a_4646_46812# a_8034_45724# 0.014576f
C6725 a_10227_46804# a_10180_45724# 0.03118f
C6726 VIN_N VREF_GND 16.4969f
C6727 VIN_P VCM 1.7189f
C6728 a_4361_42308# a_13291_42460# 0.029279f
C6729 a_n357_42282# a_9127_43156# 0.021342f
C6730 a_n755_45592# a_8387_43230# 0.010497f
C6731 a_1307_43914# a_14021_43940# 0.017312f
C6732 a_n443_42852# a_791_42968# 0.04806f
C6733 a_n913_45002# a_n1177_43370# 0.014185f
C6734 a_18248_44752# a_19006_44850# 0.056391f
C6735 a_13925_46122# a_14383_46116# 0.027606f
C6736 a_12549_44172# a_14537_43396# 0.037266f
C6737 a_584_46384# a_n2661_44458# 0.031143f
C6738 a_167_45260# a_1848_45724# 0.359783f
C6739 a_n1613_43370# a_1423_45028# 0.023846f
C6740 a_n746_45260# a_742_44458# 0.0971f
C6741 a_22223_42860# a_22400_42852# 0.154104f
C6742 a_1209_43370# VDD 0.191694f
C6743 a_20922_43172# a_20753_42852# 0.08213f
C6744 a_n2661_42834# a_n2840_43370# 0.026572f
C6745 a_6453_43914# a_n2661_42282# 0.122766f
C6746 a_22485_44484# a_22223_43948# 0.016889f
C6747 a_20512_43084# a_15493_43940# 0.021257f
C6748 a_1307_43914# a_2075_43172# 0.077359f
C6749 a_n2810_45572# a_n4318_38216# 0.023144f
C6750 a_18579_44172# a_14021_43940# 0.033047f
C6751 a_8199_44636# a_5111_44636# 0.024227f
C6752 a_10809_44734# a_3357_43084# 0.035293f
C6753 a_13059_46348# a_14309_45028# 0.050896f
C6754 a_3483_46348# a_10951_45334# 0.027449f
C6755 a_n2293_46098# a_1423_45028# 0.017396f
C6756 a_6511_45714# a_6667_45809# 0.113977f
C6757 a_6472_45840# a_6598_45938# 0.178024f
C6758 a_11459_47204# a_11599_46634# 0.019787f
C6759 a_n2497_47436# a_n1613_43370# 0.402561f
C6760 a_n1151_42308# a_4883_46098# 0.407909f
C6761 a_13717_47436# a_13487_47204# 0.061247f
C6762 a_9803_42558# a_9885_42558# 0.171361f
C6763 a_n784_42308# a_13258_32519# 0.140549f
C6764 a_n2129_43609# a_n1699_43638# 0.022218f
C6765 a_n2433_43396# a_n1917_43396# 0.108815f
C6766 a_n913_45002# a_2713_42308# 0.291963f
C6767 a_n2017_45002# a_3318_42354# 0.01513f
C6768 a_6945_45028# VDD 1.30257f
C6769 a_18184_42460# a_19987_42826# 0.208392f
C6770 a_16327_47482# a_16977_43638# 0.15941f
C6771 a_13163_45724# a_13159_45002# 0.010135f
C6772 a_10907_45822# a_6171_45002# 0.024408f
C6773 a_11823_42460# a_9482_43914# 0.033152f
C6774 a_1123_46634# a_1799_45572# 0.037438f
C6775 a_6151_47436# a_765_45546# 0.191559f
C6776 a_13507_46334# a_3090_45724# 0.020036f
C6777 a_18597_46090# a_18834_46812# 0.010699f
C6778 a_n2497_47436# a_n2293_46098# 0.039224f
C6779 a_10227_46804# a_19692_46634# 0.239326f
C6780 a_12861_44030# a_14180_46812# 0.238709f
C6781 a_n3420_38528# a_n2946_38778# 0.236674f
C6782 a_n3690_38528# a_n4064_38528# 0.085414f
C6783 a_n3565_38502# a_n2302_38778# 0.044367f
C6784 a_5934_30871# C2_N_btm 0.011047f
C6785 a_6123_31319# C4_N_btm 0.132906f
C6786 a_10341_43396# a_22591_43396# 0.172197f
C6787 en_comp CAL_N 0.023818f
C6788 a_16547_43609# a_16823_43084# 0.08061f
C6789 a_n913_45002# a_n1177_44458# 0.017911f
C6790 a_3232_43370# a_11827_44484# 0.094278f
C6791 a_3357_43084# a_5883_43914# 0.046158f
C6792 a_4185_45028# a_3626_43646# 0.035503f
C6793 a_14797_45144# a_15060_45348# 0.010598f
C6794 a_n443_42852# a_3905_42865# 0.043488f
C6795 a_16327_47482# a_18599_43230# 0.182696f
C6796 a_18834_46812# a_19123_46287# 0.039405f
C6797 a_15227_44166# a_18285_46348# 0.097182f
C6798 a_2063_45854# a_5263_45724# 0.030969f
C6799 a_2905_45572# a_2711_45572# 0.041827f
C6800 EN_VIN_BSTR_N C1_N_btm 0.110046f
C6801 C6_P_btm C5_P_btm 22.305399f
C6802 C7_P_btm C4_P_btm 0.145303f
C6803 C10_P_btm C1_P_btm 0.31753f
C6804 C9_P_btm C2_P_btm 0.141891f
C6805 C8_P_btm C3_P_btm 0.134581f
C6806 a_22629_37990# VDD 0.079474f
C6807 a_n3674_39768# a_n4064_39616# 0.464693f
C6808 a_8103_44636# VDD 0.124028f
C6809 a_1307_43914# a_5013_44260# 0.358053f
C6810 a_8103_44636# a_7640_43914# 0.101633f
C6811 a_18287_44626# a_18443_44721# 0.10279f
C6812 a_18248_44752# a_18374_44850# 0.170059f
C6813 a_15015_46420# a_2324_44458# 0.027704f
C6814 a_3483_46348# a_n1925_42282# 0.536704f
C6815 a_4791_45118# a_1423_45028# 0.721318f
C6816 a_n2312_40392# en_comp 0.036842f
C6817 a_n2312_39304# a_n2956_37592# 0.047801f
C6818 a_n881_46662# a_3357_43084# 0.028875f
C6819 a_2107_46812# a_8696_44636# 0.025973f
C6820 a_n2065_43946# a_n1761_44111# 0.617556f
C6821 a_n2017_45002# a_n1641_43230# 0.011397f
C6822 a_n913_45002# a_n1991_42858# 0.024791f
C6823 a_n1099_45572# a_n357_42282# 0.013419f
C6824 a_n1613_43370# a_6109_44484# 0.099934f
C6825 a_15682_46116# a_15765_45572# 0.015911f
C6826 a_1209_47178# a_1239_47204# 0.264529f
C6827 a_n971_45724# a_2952_47436# 0.019506f
C6828 a_n237_47217# a_2063_45854# 0.947844f
C6829 a_n1741_47186# a_3785_47178# 0.047034f
C6830 a_n2109_47186# a_4007_47204# 0.047269f
C6831 a_11341_43940# a_20974_43370# 0.013722f
C6832 a_22223_43948# a_14401_32519# 0.157135f
C6833 a_15493_43940# a_21381_43940# 0.02116f
C6834 a_22365_46825# EN_OFFSET_CAL 0.195393f
C6835 a_n2472_46090# VDD 0.224658f
C6836 a_15765_45572# a_16680_45572# 0.118759f
C6837 a_8016_46348# a_10057_43914# 0.09388f
C6838 a_8049_45260# a_n2661_43370# 0.013528f
C6839 a_6575_47204# a_8667_46634# 0.01088f
C6840 a_4915_47217# a_6755_46942# 0.260675f
C6841 a_2063_45854# a_8270_45546# 0.017994f
C6842 a_n881_46662# a_n2293_46634# 0.026189f
C6843 a_n4315_30879# a_n4064_39616# 0.034877f
C6844 a_n4064_40160# a_n3420_39616# 0.0583f
C6845 a_9145_43396# a_15095_43370# 0.213415f
C6846 a_6812_45938# VDD 0.132317f
C6847 a_20820_30879# a_14401_32519# 0.055735f
C6848 a_8696_44636# a_n2661_44458# 1.37553f
C6849 a_n2293_46634# a_n2157_46122# 0.04308f
C6850 a_8128_46384# a_8349_46414# 0.101217f
C6851 a_4915_47217# a_8049_45260# 0.022494f
C6852 a_18597_46090# a_10809_44734# 0.036294f
C6853 a_n2946_37984# VDD 0.38275f
C6854 a_n3565_38502# VCM 0.035399f
C6855 a_n4064_38528# VIN_P 0.04356f
C6856 a_9127_43156# a_8952_43230# 0.234322f
C6857 a_3539_42460# a_n2293_42282# 0.010651f
C6858 a_n97_42460# a_7309_42852# 0.024142f
C6859 en_comp a_n2472_43914# 0.014244f
C6860 a_n2433_44484# a_n1917_44484# 0.113784f
C6861 w_1575_34786# a_7174_31319# 0.01195f
C6862 a_n2293_45010# a_175_44278# 0.030523f
C6863 a_n443_42852# a_4093_43548# 0.028988f
C6864 a_n2129_44697# a_n1699_44726# 0.018607f
C6865 a_11827_44484# a_8975_43940# 0.076327f
C6866 a_1823_45246# a_4704_46090# 0.164557f
C6867 a_11453_44696# a_8696_44636# 2.67247f
C6868 a_20107_46660# a_6945_45028# 0.024966f
C6869 a_n746_45260# a_n467_45028# 0.054826f
C6870 a_13747_46662# a_11823_42460# 0.521845f
C6871 a_2804_46116# a_3147_46376# 0.017019f
C6872 a_16327_47482# a_19431_45546# 0.344862f
C6873 a_895_43940# VDD 0.318652f
C6874 a_5111_44636# a_6452_43396# 0.024938f
C6875 a_17517_44484# a_20679_44626# 0.031895f
C6876 a_n1059_45260# a_15095_43370# 0.108103f
C6877 a_21076_30879# a_n1794_35082# 0.032543f
C6878 a_n1151_42308# DATA[0] 0.088597f
C6879 a_4700_47436# VDD 0.086132f
C6880 a_526_44458# a_n2293_42282# 0.010969f
C6881 a_9290_44172# a_13291_42460# 0.078684f
C6882 a_12549_44172# a_20567_45036# 0.176249f
C6883 a_8016_46348# a_10180_45724# 0.259851f
C6884 a_n746_45260# a_n2661_43922# 0.037244f
C6885 a_10227_46804# a_10440_44484# 0.025362f
C6886 a_526_44458# a_n755_45592# 0.065199f
C6887 a_n1925_42282# a_n357_42282# 0.023161f
C6888 a_8953_45546# a_8568_45546# 0.136365f
C6889 a_8199_44636# a_9049_44484# 0.029722f
C6890 a_5937_45572# a_7499_43078# 0.033831f
C6891 a_12861_44030# a_18287_44626# 0.029719f
C6892 a_17339_46660# a_18175_45572# 0.019286f
C6893 a_n2956_38680# a_n4209_39304# 0.021073f
C6894 a_n1761_44111# a_n2129_43609# 0.029483f
C6895 a_9313_44734# a_10341_43396# 0.175125f
C6896 a_10729_43914# a_11173_44260# 0.057346f
C6897 a_10949_43914# a_10555_44260# 0.034175f
C6898 a_14955_43940# a_15493_43940# 0.110232f
C6899 a_15559_46634# VDD 0.301657f
C6900 a_8568_45546# a_8791_45572# 0.011458f
C6901 a_768_44030# a_3499_42826# 0.034429f
C6902 a_13904_45546# a_13249_42308# 0.13587f
C6903 a_10490_45724# a_10210_45822# 0.014252f
C6904 a_8270_45546# a_n2661_42834# 0.034362f
C6905 a_8953_45546# a_n2661_43370# 0.02624f
C6906 a_n971_45724# a_n97_42460# 0.581616f
C6907 a_n971_45724# a_n2661_46098# 0.023255f
C6908 a_2124_47436# a_2107_46812# 0.010665f
C6909 a_n443_46116# a_n2293_46634# 0.050675f
C6910 a_15811_47375# a_15928_47570# 0.161235f
C6911 a_17124_42282# a_4958_30871# 0.20224f
C6912 a_22223_43948# a_22223_43396# 0.025171f
C6913 a_20974_43370# a_10341_43396# 0.08579f
C6914 a_n913_45002# a_4958_30871# 0.058702f
C6915 a_3357_43084# a_3537_45260# 0.026461f
C6916 a_10193_42453# a_11827_44484# 0.121679f
C6917 a_16147_45260# a_16751_45260# 0.054632f
C6918 a_13661_43548# a_18525_43370# 0.031188f
C6919 a_n913_45002# a_n967_45348# 1.00127f
C6920 a_n2810_45028# a_n2956_37592# 6.13705f
C6921 a_n1151_42308# a_11387_46155# 0.195225f
C6922 a_n743_46660# a_3090_45724# 0.050883f
C6923 a_12549_44172# a_16721_46634# 0.013883f
C6924 a_4883_46098# a_12741_44636# 0.076276f
C6925 a_n3565_39590# C8_P_btm 0.384801f
C6926 VDAC_Pi VDAC_Ni 3.18068f
C6927 a_n4064_37984# a_n4064_37440# 0.061238f
C6928 a_19647_42308# VDD 0.227331f
C6929 a_3065_45002# VDD 0.501045f
C6930 a_2711_45572# a_11341_43940# 1.54309f
C6931 a_n2017_45002# a_n2661_42834# 0.037965f
C6932 a_16922_45042# a_17719_45144# 0.22253f
C6933 a_1423_45028# a_8103_44636# 0.064947f
C6934 a_21188_46660# a_12741_44636# 0.052893f
C6935 a_12861_44030# a_13904_45546# 0.027907f
C6936 a_6755_46942# a_10809_44734# 0.042402f
C6937 VIN_P VREF_GND 16.4969f
C6938 VIN_N VREF 0.775904f
C6939 a_n443_42852# a_685_42968# 0.104532f
C6940 en_comp a_n2433_43396# 0.036527f
C6941 a_9313_44734# a_n2293_43922# 0.026681f
C6942 a_18248_44752# a_18588_44850# 0.027606f
C6943 a_167_45260# a_997_45618# 0.052039f
C6944 a_768_44030# a_13777_45326# 0.011242f
C6945 a_n2293_46634# a_3537_45260# 0.155982f
C6946 a_10809_44734# a_8049_45260# 0.059599f
C6947 a_n746_45260# a_n452_44636# 0.042999f
C6948 a_458_43396# VDD 0.431902f
C6949 a_5534_30871# a_7174_31319# 0.038837f
C6950 a_19987_42826# a_20753_42852# 0.07365f
C6951 a_9313_44734# a_n97_42460# 1.76217f
C6952 a_1307_43914# a_1847_42826# 0.428505f
C6953 a_3067_47026# VDD 0.132018f
C6954 a_15227_44166# a_11691_44458# 0.443265f
C6955 a_3483_46348# a_10775_45002# 0.025931f
C6956 a_n443_42852# a_7499_43078# 0.375366f
C6957 a_6194_45824# a_6598_45938# 0.051162f
C6958 a_6472_45840# a_6667_45809# 0.215953f
C6959 a_6151_47436# a_10227_46804# 0.032659f
C6960 a_n1435_47204# a_13487_47204# 0.135076f
C6961 a_13717_47436# a_12861_44030# 0.319645f
C6962 a_n2129_43609# a_n2267_43396# 0.230013f
C6963 a_n2433_43396# a_n1699_43638# 0.062578f
C6964 a_n2017_45002# a_2903_42308# 0.013263f
C6965 a_21137_46414# VDD 0.219745f
C6966 a_16327_47482# a_16409_43396# 0.022593f
C6967 a_n971_45724# a_n901_43156# 0.019025f
C6968 SMPL_ON_P a_n4318_38680# 0.039103f
C6969 a_13747_46662# a_2982_43646# 0.010585f
C6970 a_n881_46662# a_6755_46942# 0.063288f
C6971 a_5815_47464# a_765_45546# 0.01398f
C6972 a_18479_47436# a_15227_44166# 0.199537f
C6973 a_18780_47178# a_18834_46812# 0.010748f
C6974 a_12861_44030# a_14035_46660# 0.153051f
C6975 a_n3565_38502# a_n4064_38528# 0.228245f
C6976 a_n4064_39072# a_n3420_37984# 0.045543f
C6977 a_n3420_39072# a_n4064_37984# 0.045827f
C6978 a_5934_30871# C1_N_btm 0.011025f
C6979 a_6123_31319# C3_N_btm 0.011333f
C6980 a_4958_30871# VDAC_P 0.017827f
C6981 a_10341_43396# a_13887_32519# 0.030175f
C6982 a_19268_43646# a_19700_43370# 0.017165f
C6983 a_16243_43396# a_16823_43084# 0.05964f
C6984 a_15743_43084# a_16664_43396# 0.01372f
C6985 a_20193_45348# a_20712_42282# 0.010791f
C6986 a_13259_45724# a_17973_43940# 0.025372f
C6987 en_comp a_n2433_44484# 0.029809f
C6988 a_n967_45348# a_n2661_44458# 0.0255f
C6989 a_18834_46812# a_18285_46348# 0.144972f
C6990 a_13885_46660# a_14513_46634# 0.101344f
C6991 a_n881_46662# a_8049_45260# 0.025172f
C6992 a_n443_46116# a_2277_45546# 0.048113f
C6993 a_4883_46098# a_16375_45002# 0.01007f
C6994 a_n2956_39768# a_n2956_38680# 0.043291f
C6995 VDAC_P VCM 11.743501f
C6996 EN_VIN_BSTR_N C0_N_btm 0.12803f
C6997 C7_P_btm C5_P_btm 0.151416f
C6998 C10_P_btm C2_P_btm 0.327137f
C6999 C9_P_btm C3_P_btm 0.137552f
C7000 C8_P_btm C4_P_btm 0.145646f
C7001 a_22725_38406# VDD 0.085997f
C7002 a_n4318_39768# a_n4064_39616# 0.047349f
C7003 a_6298_44484# VDD 1.21616f
C7004 a_3422_30871# a_n3420_37984# 0.031681f
C7005 a_5343_44458# a_5891_43370# 1.06553f
C7006 a_n443_42852# a_15781_43660# 0.22553f
C7007 a_526_44458# a_10083_42826# 0.012145f
C7008 a_18494_42460# a_17517_44484# 0.022635f
C7009 a_6298_44484# a_7640_43914# 0.031665f
C7010 a_1307_43914# a_5244_44056# 0.025291f
C7011 a_18248_44752# a_18443_44721# 0.206455f
C7012 a_17970_44736# a_18374_44850# 0.051162f
C7013 a_n357_42282# a_15743_43084# 0.055032f
C7014 a_2711_45572# a_10341_43396# 0.03441f
C7015 a_15015_46420# a_14840_46494# 0.233657f
C7016 a_3483_46348# a_526_44458# 0.134907f
C7017 a_n2312_39304# a_n2810_45028# 0.043636f
C7018 a_n2312_40392# a_n2956_37592# 0.060336f
C7019 a_n1613_43370# a_3357_43084# 0.228593f
C7020 a_15227_44166# a_n443_42852# 0.023429f
C7021 a_4190_30871# a_7174_31319# 0.153555f
C7022 a_5534_30871# a_5932_42308# 0.025879f
C7023 a_22165_42308# a_22223_42860# 0.171681f
C7024 a_n913_45002# a_n1853_43023# 0.094845f
C7025 a_3537_45260# a_743_42282# 0.033447f
C7026 a_n2956_38680# a_n4318_37592# 0.02321f
C7027 a_380_45546# a_n357_42282# 0.071576f
C7028 a_n2293_46098# a_3357_43084# 0.16657f
C7029 a_12465_44636# a_n2293_43922# 0.025736f
C7030 a_n452_45724# a_n755_45592# 0.03904f
C7031 a_n1099_45572# a_310_45028# 0.333219f
C7032 a_15682_46116# a_15903_45785# 0.011633f
C7033 a_n2497_47436# a_895_43940# 0.0309f
C7034 a_8049_45260# a_8162_45546# 0.057007f
C7035 a_n237_47217# a_584_46384# 0.645142f
C7036 a_n971_45724# a_2553_47502# 0.23907f
C7037 a_n1741_47186# a_3381_47502# 0.011573f
C7038 a_n2109_47186# a_3815_47204# 0.045952f
C7039 a_17364_32525# VCM 0.035838f
C7040 a_15493_43940# a_19741_43940# 0.027038f
C7041 a_10193_42453# a_13575_42558# 0.175489f
C7042 a_11967_42832# a_18525_43370# 0.010117f
C7043 a_n2840_46090# VDD 0.295278f
C7044 a_8953_45546# a_5883_43914# 0.262126f
C7045 a_16333_45814# a_16115_45572# 0.209641f
C7046 a_n443_46116# a_2813_43396# 0.124521f
C7047 a_15765_45572# a_16855_45546# 0.042415f
C7048 a_n1613_43370# a_n2293_46634# 0.103089f
C7049 a_14635_42282# VDD 0.369964f
C7050 a_9145_43396# a_14205_43396# 0.13322f
C7051 a_5111_44636# a_1307_43914# 0.114933f
C7052 a_2382_45260# a_2304_45348# 0.045704f
C7053 a_3065_45002# a_1423_45028# 0.017813f
C7054 a_18479_45785# a_11827_44484# 0.03055f
C7055 a_n2293_46634# a_n2293_46098# 0.062583f
C7056 a_8128_46384# a_8016_46348# 0.09182f
C7057 a_4883_46098# a_18985_46122# 0.027089f
C7058 a_n3420_37984# VDD 0.931101f
C7059 a_n2661_42282# a_6123_31319# 0.017717f
C7060 a_n97_42460# a_5837_42852# 0.011979f
C7061 a_3422_30871# a_19511_42282# 0.025144f
C7062 a_n357_42282# a_3539_42460# 0.019382f
C7063 a_n755_45592# a_3626_43646# 0.095572f
C7064 a_n2433_44484# a_n1699_44726# 0.058433f
C7065 a_n913_45002# a_n1899_43946# 0.017336f
C7066 a_n2293_45010# a_n984_44318# 0.048428f
C7067 a_2711_45572# a_n97_42460# 0.137121f
C7068 a_n2129_44697# a_n2267_44484# 0.698671f
C7069 a_1823_45246# a_4419_46090# 0.340207f
C7070 a_20411_46873# a_20708_46348# 0.081063f
C7071 a_18285_46348# a_10809_44734# 0.014976f
C7072 a_13661_43548# a_11823_42460# 0.116839f
C7073 a_16327_47482# a_18691_45572# 0.162157f
C7074 a_4791_45118# a_3357_43084# 0.144996f
C7075 a_n2497_47436# a_3065_45002# 0.022803f
C7076 a_2479_44172# VDD 0.431428f
C7077 a_5649_42852# a_5379_42460# 0.35554f
C7078 a_19237_31679# VCM 0.03748f
C7079 a_4190_30871# a_5932_42308# 0.018227f
C7080 a_1307_43914# a_4235_43370# 0.016608f
C7081 a_5111_44636# a_9396_43370# 0.203348f
C7082 a_5883_43914# a_9028_43914# 0.05428f
C7083 a_17517_44484# a_20640_44752# 0.54753f
C7084 a_4007_47204# VDD 0.41212f
C7085 a_12549_44172# a_18494_42460# 0.331306f
C7086 a_8016_46348# a_10053_45546# 0.017312f
C7087 a_n746_45260# a_n2661_42834# 0.01463f
C7088 a_n971_45724# a_n2661_43922# 0.052944f
C7089 a_15227_44166# a_2437_43646# 0.167451f
C7090 a_10227_46804# a_10334_44484# 0.020432f
C7091 a_526_44458# a_n357_42282# 0.220537f
C7092 a_5937_45572# a_8568_45546# 0.028968f
C7093 a_8199_44636# a_7499_43078# 0.859274f
C7094 a_12861_44030# a_18248_44752# 0.072535f
C7095 a_5342_30871# a_n4064_37984# 0.028465f
C7096 a_15493_43396# a_19478_44306# 0.154347f
C7097 a_10729_43914# a_10555_44260# 0.038445f
C7098 a_15682_43940# a_11341_43940# 0.021147f
C7099 a_n2956_39304# a_n4209_39304# 0.328727f
C7100 a_15368_46634# VDD 0.324877f
C7101 a_8746_45002# a_10210_45822# 0.013725f
C7102 a_n2293_46634# a_2675_43914# 0.026226f
C7103 a_8568_45546# a_8697_45572# 0.010132f
C7104 a_3090_45724# a_5891_43370# 0.166094f
C7105 a_5937_45572# a_n2661_43370# 0.202031f
C7106 a_n971_45724# a_n447_43370# 0.113797f
C7107 a_n1151_42308# a_n2438_43548# 0.093859f
C7108 a_15507_47210# a_15928_47570# 0.089677f
C7109 a_584_46384# a_1123_46634# 0.370049f
C7110 a_n2312_40392# a_n2312_39304# 0.057374f
C7111 a_4791_45118# a_n2293_46634# 0.030843f
C7112 a_16522_42674# a_4958_30871# 0.020415f
C7113 a_14401_32519# a_10341_43396# 0.133035f
C7114 a_5343_44458# a_8292_43218# 0.01105f
C7115 a_13259_45724# a_9313_44734# 0.048952f
C7116 a_13661_43548# a_18429_43548# 0.010678f
C7117 a_n1059_45260# a_n967_45348# 0.081574f
C7118 a_16147_45260# a_1307_43914# 0.150161f
C7119 a_n1151_42308# a_11133_46155# 0.162011f
C7120 a_12549_44172# a_16388_46812# 0.03419f
C7121 a_768_44030# a_13059_46348# 0.062321f
C7122 a_12465_44636# a_11415_45002# 0.375509f
C7123 a_7754_39964# VDAC_Ni 0.207118f
C7124 a_7754_40130# a_3754_38470# 0.191861f
C7125 a_19511_42282# VDD 0.244902f
C7126 a_2680_45002# VDD 0.145087f
C7127 a_n2293_45010# a_n2661_43922# 0.030818f
C7128 a_16922_45042# a_17613_45144# 0.10967f
C7129 a_13556_45296# a_15004_44636# 0.127354f
C7130 a_1423_45028# a_6298_44484# 0.103777f
C7131 a_n1151_42308# a_n1794_35082# 0.056434f
C7132 a_21363_46634# a_12741_44636# 0.053741f
C7133 a_12861_44030# a_13527_45546# 0.274077f
C7134 a_6969_46634# a_6945_45028# 0.017662f
C7135 a_12251_46660# a_12594_46348# 0.011817f
C7136 a_3090_45724# a_9290_44172# 0.196232f
C7137 a_22612_30879# a_20692_30879# 0.07827f
C7138 VIN_P VREF 0.775904f
C7139 a_15743_43084# a_22400_42852# 0.010325f
C7140 a_10193_42453# a_16823_43084# 0.03411f
C7141 a_n755_45592# a_8037_42858# 0.033004f
C7142 a_n357_42282# a_8605_42826# 0.011429f
C7143 a_9313_44734# a_n2661_43922# 0.028486f
C7144 a_12861_44030# a_16922_45042# 0.120012f
C7145 a_167_45260# a_n755_45592# 1.02724f
C7146 a_n2438_43548# a_327_44734# 0.013318f
C7147 a_8270_45546# a_8696_44636# 0.023406f
C7148 a_12594_46348# a_13259_45724# 0.012487f
C7149 a_768_44030# a_13556_45296# 0.267809f
C7150 a_11415_45002# a_2711_45572# 0.337384f
C7151 a_1823_45246# a_1848_45724# 0.028459f
C7152 a_4915_47217# a_11691_44458# 0.020788f
C7153 a_n229_43646# VDD 0.278436f
C7154 a_3080_42308# C3_N_btm 0.027071f
C7155 a_5342_30871# a_13258_32519# 0.030303f
C7156 a_19987_42826# a_20356_42852# 0.014848f
C7157 a_5663_43940# a_6101_44260# 0.013015f
C7158 a_20512_43084# a_11341_43940# 0.02996f
C7159 a_n356_44636# a_n1557_42282# 0.017569f
C7160 a_2864_46660# VDD 0.076834f
C7161 a_n2810_45572# a_n3674_38680# 0.023027f
C7162 a_19692_46634# a_11827_44484# 0.04136f
C7163 a_3483_46348# a_8953_45002# 0.121322f
C7164 a_6945_45028# a_3357_43084# 0.033591f
C7165 a_13259_45724# a_15037_45618# 0.098143f
C7166 a_6472_45840# a_6511_45714# 0.781352f
C7167 a_19321_45002# a_17517_44484# 0.264473f
C7168 a_n971_45724# a_2747_46873# 0.047519f
C7169 a_13381_47204# a_13487_47204# 0.152045f
C7170 a_n1435_47204# a_12861_44030# 0.036547f
C7171 a_1606_42308# a_4958_30871# 0.019472f
C7172 a_9223_42460# a_9377_42558# 0.010303f
C7173 COMP_P a_7174_31319# 0.029084f
C7174 a_20708_46348# VDD 0.093079f
C7175 a_2324_44458# CLK 0.035116f
C7176 a_n2433_43396# a_n2267_43396# 0.756435f
C7177 a_n2017_45002# a_2713_42308# 0.011694f
C7178 a_n443_42852# a_n2661_43370# 0.082119f
C7179 a_3090_45724# a_10807_43548# 0.031941f
C7180 SMPL_ON_P a_n3674_39304# 0.040131f
C7181 a_12861_44030# a_15743_43084# 0.01437f
C7182 a_4791_45118# a_743_42282# 0.053017f
C7183 a_12861_44030# a_13885_46660# 0.042236f
C7184 a_n4334_38528# a_n4064_38528# 0.449049f
C7185 a_n3690_38528# a_n3420_38528# 0.431104f
C7186 a_n3565_38502# a_n2946_38778# 0.406164f
C7187 a_n4209_38502# a_n2302_38778# 0.406492f
C7188 a_5934_30871# C0_N_btm 0.015126f
C7189 a_6123_31319# C2_N_btm 0.01106f
C7190 a_1606_42308# VCM 0.152876f
C7191 a_1273_38525# a_2113_38308# 0.325472f
C7192 a_4921_42308# VDD 0.214995f
C7193 a_10341_43396# a_22223_43396# 0.038582f
C7194 a_12281_43396# a_4361_42308# 0.021275f
C7195 a_6293_42852# a_5755_42852# 0.114235f
C7196 a_16137_43396# a_16823_43084# 0.038492f
C7197 a_n356_44636# a_5934_30871# 0.095373f
C7198 a_n2661_45010# a_949_44458# 0.071688f
C7199 a_375_42282# a_n2661_43370# 0.012518f
C7200 a_13259_45724# a_17737_43940# 0.016944f
C7201 en_comp a_n2661_44458# 0.030481f
C7202 a_4185_45028# a_2982_43646# 0.243496f
C7203 a_11823_42460# a_11967_42832# 0.573139f
C7204 a_13885_46660# a_14180_46812# 0.150851f
C7205 a_17609_46634# a_18285_46348# 0.115413f
C7206 a_n443_46116# a_1609_45822# 0.096281f
C7207 a_12465_44636# a_13259_45724# 0.096616f
C7208 a_n2956_39768# a_n2956_39304# 0.098523f
C7209 a_2107_46812# a_2324_44458# 0.051531f
C7210 a_22629_38406# VDD 0.315181f
C7211 VDAC_P VREF_GND 0.203715f
C7212 EN_VIN_BSTR_N C0_dummy_N_btm 0.026355f
C7213 C7_P_btm C6_P_btm 26.0771f
C7214 C8_P_btm C5_P_btm 0.145019f
C7215 C10_P_btm C3_P_btm 0.321945f
C7216 C9_P_btm C4_P_btm 0.154834f
C7217 CAL_P RST_Z 0.551895f
C7218 a_n3674_39768# a_n3420_39616# 0.073948f
C7219 a_5518_44484# VDD 0.40715f
C7220 a_15743_43084# a_22223_42860# 0.021215f
C7221 a_n443_42852# a_15681_43442# 0.035093f
C7222 a_526_44458# a_8952_43230# 0.039329f
C7223 a_18184_42460# a_17517_44484# 0.020871f
C7224 a_6298_44484# a_6109_44484# 0.068396f
C7225 a_1307_43914# a_3905_42865# 0.224019f
C7226 a_18248_44752# a_18287_44626# 0.633819f
C7227 a_18597_46090# a_13258_32519# 0.023292f
C7228 a_3147_46376# a_526_44458# 0.352f
C7229 a_13747_46662# a_18799_45938# 0.028671f
C7230 a_n2312_40392# a_n2810_45028# 0.055228f
C7231 a_743_42282# a_13258_32519# 0.030886f
C7232 a_n2472_43914# a_n2065_43946# 0.039807f
C7233 a_n863_45724# a_n2293_42282# 0.028166f
C7234 a_n2017_45002# a_n1991_42858# 0.053113f
C7235 a_n1059_45260# a_n1853_43023# 0.03561f
C7236 a_n2956_39304# a_n4318_37592# 0.023347f
C7237 a_n357_42282# a_21195_42852# 0.09377f
C7238 a_13661_43548# a_14539_43914# 0.193767f
C7239 a_n2661_45546# a_3316_45546# 0.027868f
C7240 a_12465_44636# a_n2661_43922# 0.17969f
C7241 a_380_45546# a_310_45028# 0.057269f
C7242 a_n863_45724# a_n755_45592# 1.76733f
C7243 a_13259_45724# a_2711_45572# 1.26722f
C7244 a_2324_44458# a_15903_45785# 0.017867f
C7245 a_21076_30879# a_20447_31679# 0.055814f
C7246 a_n1741_47186# a_n1151_42308# 2.98024f
C7247 a_n971_45724# a_2063_45854# 0.164981f
C7248 a_n2109_47186# a_3785_47178# 0.190973f
C7249 a_n746_45260# a_584_46384# 0.491308f
C7250 a_17364_32525# VREF_GND 0.048253f
C7251 COMP_P a_5932_42308# 0.02968f
C7252 a_n2661_42282# a_3080_42308# 0.161683f
C7253 a_11341_43940# a_21381_43940# 0.034147f
C7254 a_20512_43084# a_10341_43396# 0.758407f
C7255 a_11967_42832# a_18429_43548# 0.019775f
C7256 a_5937_45572# a_5883_43914# 0.454323f
C7257 a_8199_44636# a_9838_44484# 0.024921f
C7258 a_4646_46812# a_n2661_42282# 0.025072f
C7259 a_10809_44734# a_11691_44458# 0.354084f
C7260 a_20202_43084# a_9313_44734# 0.044152f
C7261 a_15765_45572# a_16115_45572# 0.20669f
C7262 a_15599_45572# a_16680_45572# 0.102355f
C7263 a_2324_44458# a_n2661_44458# 0.134417f
C7264 a_12549_44172# a_19321_45002# 0.238866f
C7265 a_n4315_30879# a_n3420_39616# 0.03477f
C7266 a_n4064_40160# a_n3565_39590# 0.031111f
C7267 a_13291_42460# VDD 0.546706f
C7268 a_9145_43396# a_14358_43442# 0.053427f
C7269 a_n2956_37592# a_n3565_38502# 0.024508f
C7270 a_5147_45002# a_1307_43914# 0.032106f
C7271 a_2274_45254# a_2304_45348# 0.062682f
C7272 a_6171_45002# a_14537_43396# 0.054973f
C7273 a_20202_43084# a_20974_43370# 0.026132f
C7274 a_2437_43646# a_n2661_43370# 0.033415f
C7275 a_10903_43370# a_11341_43940# 0.061205f
C7276 a_n1151_42308# a_10586_45546# 0.02493f
C7277 a_11453_44696# a_2324_44458# 0.023884f
C7278 a_8128_46384# a_7920_46348# 0.197919f
C7279 a_n881_46662# a_5937_45572# 0.195456f
C7280 a_n1613_43370# a_8953_45546# 0.024821f
C7281 a_18597_46090# a_6945_45028# 0.049383f
C7282 a_18479_47436# a_10809_44734# 0.04504f
C7283 a_4883_46098# a_18819_46122# 0.054304f
C7284 a_n3690_38304# VDD 0.363068f
C7285 a_n4209_38502# VCM 0.035344f
C7286 a_n3565_38502# VREF 0.056031f
C7287 a_n3420_38528# VIN_P 0.052378f
C7288 a_8605_42826# a_8952_43230# 0.051162f
C7289 a_n357_42282# a_3626_43646# 0.020238f
C7290 a_n2433_44484# a_n2267_44484# 0.730194f
C7291 a_14537_43396# a_14673_44172# 0.044194f
C7292 a_n913_45002# a_n1761_44111# 0.036392f
C7293 a_n2293_45010# a_n809_44244# 0.041966f
C7294 a_n443_42852# a_1568_43370# 0.038016f
C7295 a_1823_45246# a_4185_45028# 0.081652f
C7296 a_4915_47217# a_2437_43646# 0.114772f
C7297 a_17829_46910# a_10809_44734# 0.02024f
C7298 a_5807_45002# a_11823_42460# 0.022934f
C7299 a_16327_47482# a_18909_45814# 0.16767f
C7300 a_2698_46116# a_2804_46116# 0.313533f
C7301 a_2127_44172# VDD 0.138239f
C7302 a_5649_42852# a_5267_42460# 0.016079f
C7303 a_5111_44636# a_8791_43396# 0.05316f
C7304 a_5883_43914# a_8333_44056# 0.152643f
C7305 a_17517_44484# a_20362_44736# 0.047565f
C7306 a_3815_47204# VDD 0.260661f
C7307 a_n913_45002# a_14579_43548# 0.239851f
C7308 a_12549_44172# a_18184_42460# 0.03123f
C7309 a_n971_45724# a_n2661_42834# 0.165951f
C7310 a_n2438_43548# a_n2293_42834# 0.138621f
C7311 a_8199_44636# a_8568_45546# 0.141772f
C7312 a_19328_44172# a_19478_44306# 0.188181f
C7313 a_10405_44172# a_10555_44260# 0.085098f
C7314 a_14976_45028# VDD 0.484864f
C7315 a_11823_42460# a_15143_45578# 0.120787f
C7316 a_10193_42453# a_10210_45822# 0.026406f
C7317 a_n2497_47436# a_n229_43646# 0.022782f
C7318 a_13507_46334# a_15493_43940# 0.021188f
C7319 a_8199_44636# a_n2661_43370# 0.126664f
C7320 a_n1151_42308# a_n743_46660# 0.195953f
C7321 a_15811_47375# a_12549_44172# 0.024519f
C7322 a_9313_45822# a_5807_45002# 0.031627f
C7323 a_16104_42674# a_4958_30871# 0.029272f
C7324 a_19479_31679# a_13258_32519# 0.054577f
C7325 a_20205_31679# C4_N_btm 0.042623f
C7326 a_n2017_45002# a_4958_30871# 0.053522f
C7327 a_11341_43940# a_5649_42852# 0.01232f
C7328 a_18051_46116# VDD 0.189782f
C7329 a_21381_43940# a_10341_43396# 0.03047f
C7330 a_n2017_45002# a_n967_45348# 0.095287f
C7331 a_3357_43084# a_3065_45002# 0.316449f
C7332 a_4646_46812# a_7112_43396# 0.07278f
C7333 a_16147_45260# a_16019_45002# 0.186254f
C7334 a_n1151_42308# a_11189_46129# 0.12414f
C7335 a_13507_46334# a_12741_44636# 0.137731f
C7336 a_6545_47178# a_6419_46155# 0.080336f
C7337 a_12549_44172# a_13059_46348# 0.808395f
C7338 a_22223_47212# a_22365_46825# 0.011422f
C7339 a_n3420_37984# a_n4064_37440# 7.43287f
C7340 a_n2946_37984# a_n2946_37690# 0.050477f
C7341 a_n4064_37984# a_n3420_37440# 0.053897f
C7342 a_2382_45260# VDD 1.6285f
C7343 a_9290_44172# a_12281_43396# 0.36475f
C7344 a_10903_43370# a_10341_43396# 0.042836f
C7345 a_20820_30879# a_13678_32519# 0.053259f
C7346 a_n2293_45010# a_n2661_42834# 0.083461f
C7347 a_16922_45042# a_17023_45118# 0.099834f
C7348 a_18479_45785# a_19279_43940# 0.019159f
C7349 a_21076_30879# a_13467_32519# 0.055522f
C7350 a_9482_43914# a_15004_44636# 0.34299f
C7351 a_13556_45296# a_13720_44458# 0.212774f
C7352 a_1423_45028# a_5518_44484# 0.047243f
C7353 a_10227_46804# a_7499_43078# 0.033512f
C7354 a_20623_46660# a_12741_44636# 0.034292f
C7355 a_12861_44030# a_13163_45724# 0.098707f
C7356 a_768_44030# a_2957_45546# 0.027276f
C7357 a_6755_46942# a_6945_45028# 0.024014f
C7358 a_22612_30879# a_20205_31679# 0.111294f
C7359 a_21588_30879# a_20692_30879# 0.056225f
C7360 a_3422_30871# CAL_P 0.083836f
C7361 a_15433_44458# VDD 0.201121f
C7362 a_n2956_37592# a_n4318_39304# 0.023222f
C7363 a_n2017_45002# a_n1917_43396# 0.01343f
C7364 a_2437_43646# a_1568_43370# 0.058471f
C7365 a_14539_43914# a_11967_42832# 0.512158f
C7366 a_n357_42282# a_8037_42858# 0.048934f
C7367 a_9313_44734# a_n2661_42834# 0.02321f
C7368 a_167_45260# a_n357_42282# 0.148401f
C7369 a_n2438_43548# a_413_45260# 0.032468f
C7370 a_n2293_46634# a_3065_45002# 0.102991f
C7371 a_12549_44172# a_13556_45296# 0.030045f
C7372 a_12891_46348# a_13777_45326# 0.03955f
C7373 a_768_44030# a_9482_43914# 0.77718f
C7374 a_n746_45260# a_n1177_44458# 0.064145f
C7375 a_19987_42826# a_20256_42852# 0.015204f
C7376 a_3080_42308# C2_N_btm 0.108823f
C7377 a_3524_46660# VDD 0.278519f
C7378 a_3483_46348# a_8191_45002# 0.081038f
C7379 a_12549_44172# a_20362_44736# 0.015111f
C7380 a_22223_46124# a_22223_45572# 0.025171f
C7381 a_10809_44734# a_2437_43646# 0.13907f
C7382 a_6194_45824# a_6511_45714# 0.102325f
C7383 a_n1435_47204# a_13717_47436# 0.196889f
C7384 a_9223_42460# a_9293_42558# 0.011552f
C7385 a_n2433_43396# a_n2129_43609# 0.283605f
C7386 a_19900_46494# VDD 0.279179f
C7387 en_comp a_1606_42308# 0.022666f
C7388 a_16327_47482# a_16243_43396# 0.295263f
C7389 a_10903_43370# a_n2293_43922# 0.029114f
C7390 a_11823_42460# a_13017_45260# 0.030503f
C7391 a_7499_43078# a_1307_43914# 0.109806f
C7392 a_8049_45260# a_8103_44636# 0.012205f
C7393 a_10227_46804# a_15227_44166# 0.013242f
C7394 a_171_46873# a_n2661_46098# 0.168482f
C7395 a_383_46660# a_479_46660# 0.013793f
C7396 a_9804_47204# a_9863_46634# 0.017882f
C7397 a_4915_47217# a_765_45546# 0.169406f
C7398 a_n1925_46634# a_3699_46634# 0.014429f
C7399 a_5742_30871# EN_VIN_BSTR_N 0.643089f
C7400 a_1666_39043# a_2684_37794# 0.193789f
C7401 a_n4209_38502# a_n4064_38528# 0.265711f
C7402 a_n3565_38502# a_n3420_38528# 0.278952f
C7403 a_n3565_39304# a_n4064_37984# 0.028081f
C7404 a_n4064_39072# a_n3565_38216# 0.030681f
C7405 a_n3420_39072# a_n3420_37984# 0.046468f
C7406 a_6123_31319# C1_N_btm 0.011005f
C7407 a_4958_30871# VDAC_N 0.021971f
C7408 a_15743_43084# a_19268_43646# 0.010228f
C7409 a_10341_43396# a_5649_42852# 0.049047f
C7410 a_n2661_45010# a_742_44458# 0.694478f
C7411 a_n2293_45010# a_n1352_44484# 0.020183f
C7412 a_n2017_45002# a_n1917_44484# 0.012037f
C7413 a_10903_43370# a_n97_42460# 0.021999f
C7414 a_n2661_46634# a_10809_44734# 0.023983f
C7415 a_13885_46660# a_14035_46660# 0.25868f
C7416 a_17609_46634# a_17829_46910# 0.111805f
C7417 a_15227_44166# a_17339_46660# 0.524034f
C7418 a_n971_45724# a_3775_45552# 0.091275f
C7419 a_n443_46116# a_n443_42852# 0.145452f
C7420 a_2063_45854# a_2711_45572# 0.185507f
C7421 CAL_P VDD 22.475801f
C7422 VDAC_N VCM 11.7445f
C7423 C9_P_btm C5_P_btm 0.150576f
C7424 C10_P_btm C4_P_btm 0.703336f
C7425 C8_P_btm C6_P_btm 0.163943f
C7426 a_n3674_39768# a_n3690_39616# 0.07198f
C7427 a_5343_44458# VDD 0.49245f
C7428 a_526_44458# a_9127_43156# 0.054699f
C7429 a_626_44172# a_895_43940# 0.038336f
C7430 a_19778_44110# a_17517_44484# 0.018823f
C7431 a_5518_44484# a_6109_44484# 0.050093f
C7432 a_5343_44458# a_7640_43914# 0.152634f
C7433 a_17970_44736# a_18287_44626# 0.102355f
C7434 a_11691_44458# a_11541_44484# 0.037586f
C7435 a_3537_45260# a_8333_44056# 0.012371f
C7436 a_1307_43914# a_3600_43914# 0.153686f
C7437 a_14493_46090# a_14840_46494# 0.051162f
C7438 a_19321_45002# a_19431_45546# 0.029441f
C7439 a_13747_46662# a_18596_45572# 0.01625f
C7440 a_n881_46662# a_2437_43646# 0.084076f
C7441 a_8199_44636# a_10809_44734# 0.022266f
C7442 a_14209_32519# a_4958_30871# 0.030901f
C7443 a_n2956_38680# a_n3674_38216# 0.02335f
C7444 a_3065_45002# a_743_42282# 0.040577f
C7445 a_n2017_45002# a_n1853_43023# 0.03086f
C7446 a_n357_42282# a_21356_42826# 0.156735f
C7447 a_5807_45002# a_14539_43914# 0.066683f
C7448 a_13661_43548# a_16112_44458# 0.053099f
C7449 a_n2661_45546# a_3218_45724# 0.010947f
C7450 a_n1079_45724# a_n755_45592# 0.109544f
C7451 a_n863_45724# a_n357_42282# 0.172013f
C7452 a_380_45546# a_n1099_45572# 0.148825f
C7453 a_2324_44458# a_15599_45572# 0.042604f
C7454 a_15227_44166# a_1307_43914# 0.059667f
C7455 a_n971_45724# a_584_46384# 0.152617f
C7456 a_n237_47217# a_1431_47204# 0.045044f
C7457 a_n1741_47186# a_3160_47472# 0.012286f
C7458 a_n2109_47186# a_3381_47502# 0.035813f
C7459 a_2123_42473# a_2351_42308# 0.084895f
C7460 a_21115_43940# a_21381_43940# 0.073198f
C7461 a_n2293_43922# a_5649_42852# 1.78418f
C7462 a_21076_30879# RST_Z 0.052228f
C7463 a_5937_45572# a_8701_44490# 0.022661f
C7464 a_8016_46348# a_10157_44484# 0.016596f
C7465 a_3483_46348# a_16979_44734# 0.173123f
C7466 a_15765_45572# a_16333_45814# 0.17072f
C7467 a_15599_45572# a_16855_45546# 0.043567f
C7468 a_n2312_39304# a_n4318_39304# 0.023404f
C7469 a_n443_42852# a_3537_45260# 0.567413f
C7470 a_7903_47542# a_8145_46902# 0.010369f
C7471 a_n881_46662# a_n2661_46634# 0.035376f
C7472 a_768_44030# a_13747_46662# 0.434325f
C7473 a_13003_42852# VDD 0.132655f
C7474 a_n4064_40160# a_n4334_39616# 0.014656f
C7475 a_n2810_45028# a_n3565_38502# 0.031875f
C7476 a_9145_43396# a_14579_43548# 0.024497f
C7477 a_8685_43396# a_10341_43396# 2.41562f
C7478 a_17715_44484# a_17737_43940# 0.289085f
C7479 a_10775_45002# a_10951_45334# 0.185422f
C7480 a_2382_45260# a_1423_45028# 0.036767f
C7481 a_6171_45002# a_14180_45002# 0.012672f
C7482 a_n1613_43370# a_5937_45572# 0.117604f
C7483 a_18780_47178# a_6945_45028# 0.013003f
C7484 a_4883_46098# a_17957_46116# 0.013641f
C7485 a_n3565_38216# VDD 0.903914f
C7486 a_11206_38545# CAL_N 0.050483f
C7487 a_8037_42858# a_8952_43230# 0.118759f
C7488 a_2982_43646# a_n2293_42282# 0.010686f
C7489 a_n2661_44458# a_n2267_44484# 0.046548f
C7490 a_n2433_44484# a_n2129_44697# 0.130072f
C7491 a_n913_45002# a_n2065_43946# 0.018244f
C7492 a_n2293_45010# a_n1549_44318# 0.014826f
C7493 a_n2017_45002# a_n1899_43946# 0.017371f
C7494 a_n443_42852# a_1049_43396# 0.047375f
C7495 a_n1059_45260# a_n1761_44111# 0.535535f
C7496 a_n755_45592# a_2982_43646# 0.221452f
C7497 a_3357_43084# a_2479_44172# 0.0305f
C7498 a_11415_45002# a_10903_43370# 0.085164f
C7499 a_n746_45260# a_n967_45348# 0.028689f
C7500 a_n443_46116# a_2437_43646# 0.410719f
C7501 a_n1741_47186# a_413_45260# 0.026099f
C7502 a_584_46384# a_n2293_45010# 0.02901f
C7503 a_11599_46634# a_18596_45572# 0.01377f
C7504 a_16327_47482# a_18341_45572# 0.04767f
C7505 a_n2497_47436# a_2382_45260# 0.042349f
C7506 a_n2293_46098# a_5937_45572# 0.078393f
C7507 a_765_45546# a_10809_44734# 2.52248f
C7508 a_453_43940# VDD 0.225569f
C7509 a_19237_31679# VREF 0.046045f
C7510 a_5342_30871# a_14635_42282# 0.012123f
C7511 a_17730_32519# VCM 0.068103f
C7512 a_n4318_38680# a_n3674_37592# 0.02489f
C7513 a_1307_43914# a_1756_43548# 0.267667f
C7514 a_5111_44636# a_8147_43396# 0.08322f
C7515 a_3537_45260# a_6655_43762# 0.031868f
C7516 a_626_44172# a_458_43396# 0.065365f
C7517 a_17517_44484# a_20159_44458# 0.026718f
C7518 a_n1059_45260# a_14579_43548# 0.250544f
C7519 SMPL_ON_N a_22537_40625# 0.028814f
C7520 a_3785_47178# VDD 0.387755f
C7521 a_12549_44172# a_19778_44110# 0.294084f
C7522 a_3483_46348# a_11823_42460# 0.377948f
C7523 a_8199_44636# a_8162_45546# 0.119979f
C7524 a_5534_30871# a_n4064_37984# 0.047233f
C7525 a_5342_30871# a_n3420_37984# 0.028488f
C7526 a_9313_44734# a_15095_43370# 0.039448f
C7527 a_n2293_43922# a_8685_43396# 0.026511f
C7528 a_19328_44172# a_15493_43396# 0.019584f
C7529 a_7542_44172# a_7499_43940# 0.157633f
C7530 a_n755_45592# a_8325_42308# 0.040306f
C7531 a_3090_45724# VDD 2.05725f
C7532 a_11823_42460# a_14495_45572# 0.023559f
C7533 a_8162_45546# a_8192_45572# 0.134163f
C7534 a_2711_45572# a_15861_45028# 0.02395f
C7535 a_3090_45724# a_7640_43914# 0.020595f
C7536 a_5937_45572# a_8704_45028# 0.010036f
C7537 a_n971_45724# a_n1177_43370# 0.014733f
C7538 a_3160_47472# a_n743_46660# 0.011563f
C7539 a_11599_46634# a_768_44030# 0.018831f
C7540 a_1431_47204# a_1123_46634# 0.012069f
C7541 a_n1151_42308# a_n1021_46688# 0.105326f
C7542 a_13717_47436# a_13759_47204# 0.013673f
C7543 a_13487_47204# a_13569_47204# 0.014524f
C7544 a_n443_46116# a_n2661_46634# 0.121882f
C7545 a_4646_46812# a_7287_43370# 0.07176f
C7546 a_n2661_45010# a_n467_45028# 0.227953f
C7547 a_12891_46348# a_13059_46348# 0.372745f
C7548 a_n1151_42308# a_9290_44172# 0.10853f
C7549 a_n881_46662# a_765_45546# 0.333008f
C7550 a_2063_45854# a_12005_46116# 0.051126f
C7551 a_4791_45118# a_5937_45572# 0.151145f
C7552 a_20916_46384# a_19692_46634# 0.117693f
C7553 a_9313_45822# a_3483_46348# 0.087132f
C7554 a_n4209_39590# C9_P_btm 0.786375f
C7555 a_2274_45254# VDD 0.256655f
C7556 a_413_45260# SINGLE_ENDED 0.037852f
C7557 a_n1925_42282# a_3539_42460# 0.024736f
C7558 a_n2661_45010# a_n2661_43922# 0.111071f
C7559 a_9482_43914# a_13720_44458# 0.188323f
C7560 a_1423_45028# a_5343_44458# 0.128331f
C7561 a_n743_46660# a_16375_45002# 0.03035f
C7562 a_8270_45546# a_2324_44458# 0.039817f
C7563 a_20841_46902# a_12741_44636# 0.043075f
C7564 a_16327_47482# a_10193_42453# 0.163668f
C7565 a_n1613_43370# a_n443_42852# 0.062474f
C7566 a_22000_46634# a_20202_43084# 0.154237f
C7567 a_21588_30879# a_20205_31679# 0.058932f
C7568 a_12861_44030# a_12791_45546# 0.248928f
C7569 a_743_42282# a_14635_42282# 0.02914f
C7570 a_14815_43914# VDD 0.307386f
C7571 a_n913_45002# a_n2129_43609# 0.023791f
C7572 a_n755_45592# a_7871_42858# 0.033537f
C7573 a_n357_42282# a_7765_42852# 0.042157f
C7574 a_n2810_45028# a_n4318_39304# 0.023142f
C7575 a_1823_45246# a_n2293_42282# 0.03994f
C7576 a_n743_46660# a_413_45260# 0.031499f
C7577 a_n2293_46634# a_2680_45002# 0.017731f
C7578 a_10227_46804# a_n2661_43370# 0.033611f
C7579 a_526_44458# a_n1925_42282# 0.213917f
C7580 a_12549_44172# a_9482_43914# 0.06308f
C7581 a_12891_46348# a_13556_45296# 0.29495f
C7582 a_167_45260# a_310_45028# 0.035247f
C7583 a_1823_45246# a_n755_45592# 0.390511f
C7584 a_10903_43370# a_13259_45724# 0.600111f
C7585 a_n2293_46098# a_n443_42852# 0.086171f
C7586 a_5534_30871# a_13258_32519# 0.04166f
C7587 a_4190_30871# a_n4064_37984# 0.032018f
C7588 a_3080_42308# C1_N_btm 0.011373f
C7589 a_17538_32519# VCM 0.0424f
C7590 a_3699_46634# VDD 0.347281f
C7591 a_2711_45572# a_3775_45552# 0.044123f
C7592 a_n357_42282# a_11823_42460# 0.063073f
C7593 a_20708_46348# a_3357_43084# 0.017189f
C7594 a_8199_44636# a_3537_45260# 0.199536f
C7595 a_5907_45546# a_6511_45714# 0.043475f
C7596 a_6194_45824# a_6472_45840# 0.118423f
C7597 a_13747_46662# a_17517_44484# 0.022087f
C7598 a_4915_47217# a_10227_46804# 0.062269f
C7599 a_5934_30871# a_5742_30871# 16.7261f
C7600 a_20075_46420# VDD 0.347847f
C7601 a_n913_45002# a_2351_42308# 0.023646f
C7602 a_3090_45724# a_10729_43914# 0.135702f
C7603 a_n1613_43370# a_6655_43762# 0.013792f
C7604 a_10903_43370# a_n2661_43922# 0.039051f
C7605 a_11823_42460# a_11963_45334# 0.110904f
C7606 a_20202_43084# a_20512_43084# 0.130366f
C7607 a_n443_46116# a_765_45546# 0.297346f
C7608 a_n2438_43548# a_2443_46660# 0.237765f
C7609 a_n3565_38502# a_n3690_38528# 0.246863f
C7610 a_n4334_38528# a_n3420_38528# 0.015595f
C7611 a_n4209_38502# a_n2946_38778# 0.022704f
C7612 a_6123_31319# C0_N_btm 0.018968f
C7613 a_3905_42558# VDD 0.176395f
C7614 a_10341_43396# a_13678_32519# 0.011962f
C7615 a_n356_44636# a_6123_31319# 0.169259f
C7616 a_n2661_45010# a_n452_44636# 0.020671f
C7617 a_n913_45002# a_n2129_44697# 0.017685f
C7618 a_n2956_37592# a_n4318_40392# 2.71462f
C7619 a_14180_45002# a_14403_45348# 0.011458f
C7620 a_4883_46098# a_13259_45724# 0.011246f
C7621 a_17609_46634# a_765_45546# 0.256159f
C7622 a_4791_45118# a_n443_42852# 0.02747f
C7623 VDAC_N VREF_GND 0.203821f
C7624 C10_P_btm C5_P_btm 0.51798f
C7625 C9_P_btm C6_P_btm 0.165353f
C7626 C8_P_btm C7_P_btm 31.072699f
C7627 a_n3674_39768# a_n3565_39590# 0.128683f
C7628 a_4743_44484# VDD 0.266843f
C7629 a_19721_31679# VCM 0.03544f
C7630 a_13507_46334# a_18907_42674# 0.202065f
C7631 a_4223_44672# a_5891_43370# 0.020744f
C7632 a_526_44458# a_8387_43230# 0.032585f
C7633 a_5343_44458# a_6109_44484# 0.285594f
C7634 a_5518_44484# a_5826_44734# 0.017351f
C7635 a_18597_46090# a_19511_42282# 0.156698f
C7636 a_5111_44636# a_n2661_42282# 0.025961f
C7637 a_7499_43078# a_8791_43396# 0.04623f
C7638 a_17767_44458# a_18287_44626# 0.043567f
C7639 a_17970_44736# a_18248_44752# 0.117156f
C7640 a_1307_43914# a_2998_44172# 0.233292f
C7641 a_13259_45724# a_5649_42852# 1.92021f
C7642 a_13925_46122# a_14840_46494# 0.118759f
C7643 a_2804_46116# a_2981_46116# 0.134298f
C7644 a_13747_46662# a_19256_45572# 0.040187f
C7645 a_n1613_43370# a_2437_43646# 0.027497f
C7646 a_1138_42852# a_1337_46116# 0.039951f
C7647 a_5937_45572# a_6945_45028# 0.22046f
C7648 a_4190_30871# a_13258_32519# 0.039476f
C7649 a_n2017_45002# a_n2157_42858# 0.040763f
C7650 a_n2956_39304# a_n3674_38216# 0.023505f
C7651 a_n357_42282# a_20922_43172# 0.059485f
C7652 a_13661_43548# a_15004_44636# 0.012894f
C7653 a_n2293_45546# a_n755_45592# 0.061822f
C7654 a_n971_45724# a_n1331_43914# 0.015263f
C7655 a_3090_45724# a_1423_45028# 0.450367f
C7656 a_n2293_46098# a_2437_43646# 0.027185f
C7657 a_n2438_43548# a_949_44458# 1.62911f
C7658 a_4883_46098# a_n2661_43922# 0.022558f
C7659 a_21076_30879# a_19963_31679# 0.055082f
C7660 a_n2497_47436# a_453_43940# 0.09742f
C7661 a_n452_45724# a_n1099_45572# 0.053931f
C7662 a_n863_45724# a_310_45028# 0.033427f
C7663 a_17364_32525# VIN_N 0.03818f
C7664 a_n785_47204# a_327_47204# 0.237391f
C7665 a_n971_45724# a_2124_47436# 0.352461f
C7666 a_n237_47217# a_1239_47204# 0.203126f
C7667 a_n1741_47186# a_2905_45572# 0.012244f
C7668 a_n2109_47186# a_n1151_42308# 0.235661f
C7669 a_n1736_43218# VDD 0.082445f
C7670 a_14209_32519# VREF_GND 0.034351f
C7671 a_15493_43940# a_18533_43940# 0.052096f
C7672 a_2479_44172# a_2813_43396# 0.115852f
C7673 a_10193_42453# a_11633_42558# 0.017236f
C7674 a_21076_30879# VDD 1.23089f
C7675 a_8199_44636# a_8701_44490# 0.25266f
C7676 a_3483_46348# a_14539_43914# 1.24006f
C7677 a_15599_45572# a_16115_45572# 0.105995f
C7678 a_n2312_40392# a_n4318_39304# 0.025248f
C7679 a_6151_47436# a_9863_46634# 0.0481f
C7680 a_n2497_47436# a_3090_45724# 0.16041f
C7681 a_n1613_43370# a_n2661_46634# 0.279652f
C7682 a_768_44030# a_13661_43548# 0.175469f
C7683 a_12549_44172# a_13747_46662# 0.072812f
C7684 a_n4064_40160# a_n4209_39590# 0.059936f
C7685 a_n2302_40160# a_n2216_40160# 0.011479f
C7686 a_n4315_30879# a_n3565_39590# 0.027163f
C7687 a_n4334_40480# a_n4334_39616# 0.050585f
C7688 a_9145_43396# a_13667_43396# 0.074541f
C7689 a_n2956_37592# a_n4209_38502# 0.090878f
C7690 a_20202_43084# a_21381_43940# 0.108097f
C7691 a_19431_45546# a_19778_44110# 0.010264f
C7692 a_6171_45002# a_13777_45326# 0.010994f
C7693 a_10193_42453# a_n356_44636# 2.49128f
C7694 a_n2472_46634# a_n2472_46090# 0.026152f
C7695 a_10227_46804# a_10809_44734# 0.17883f
C7696 a_6755_46942# a_15368_46634# 0.033754f
C7697 a_18479_47436# a_6945_45028# 0.348097f
C7698 a_4883_46098# a_18189_46348# 0.012818f
C7699 a_768_44030# a_4185_45028# 0.022613f
C7700 a_n4334_38304# VDD 0.385989f
C7701 a_n4209_38502# VREF 0.059621f
C7702 a_n3565_38502# VIN_P 0.028513f
C7703 a_8605_42826# a_8387_43230# 0.209641f
C7704 a_8037_42858# a_9127_43156# 0.042737f
C7705 a_n2661_44458# a_n2129_44697# 0.035428f
C7706 a_n2017_45002# a_n1761_44111# 0.02974f
C7707 a_n443_42852# a_1209_43370# 0.010053f
C7708 a_n357_42282# a_2982_43646# 0.04908f
C7709 a_n2293_45010# a_n1331_43914# 0.02919f
C7710 a_n2293_42834# a_5891_43370# 0.669411f
C7711 a_13259_45724# a_8685_43396# 0.031693f
C7712 a_16327_47482# a_18479_45785# 0.841261f
C7713 a_1823_45246# a_3483_46348# 0.070929f
C7714 a_n971_45724# a_n967_45348# 0.581053f
C7715 a_12465_44636# a_8696_44636# 0.038471f
C7716 a_11599_46634# a_19256_45572# 0.051691f
C7717 a_2521_46116# a_2698_46116# 0.159555f
C7718 a_15368_46634# a_8049_45260# 0.032468f
C7719 a_5342_30871# a_13291_42460# 0.031084f
C7720 a_19237_31679# VIN_N 0.028884f
C7721 a_17730_32519# VREF_GND 0.241027f
C7722 a_4361_42308# a_5379_42460# 0.045451f
C7723 a_1414_42308# VDD 0.657887f
C7724 a_n3674_39304# a_n3674_37592# 0.024803f
C7725 a_743_42282# a_4921_42308# 0.015669f
C7726 a_1307_43914# a_1568_43370# 0.182552f
C7727 a_5111_44636# a_7112_43396# 0.041581f
C7728 a_17517_44484# a_19615_44636# 0.018532f
C7729 a_3381_47502# VDD 0.197761f
C7730 a_n2312_39304# a_n4318_40392# 0.023465f
C7731 a_12281_43396# VDD 0.341026f
C7732 a_9672_43914# a_9895_44260# 0.011458f
C7733 a_15009_46634# VDD 0.205396f
C7734 a_7281_43914# a_7499_43940# 0.08213f
C7735 a_13163_45724# a_13527_45546# 0.124682f
C7736 a_10053_45546# a_10210_45822# 0.18824f
C7737 a_13507_46334# a_11341_43940# 0.162723f
C7738 a_11823_42460# a_13249_42308# 0.360411f
C7739 a_2711_45572# a_8696_44636# 0.02621f
C7740 a_16327_47482# a_14021_43940# 0.061511f
C7741 a_8016_46348# a_n2661_43370# 0.028709f
C7742 a_2905_45572# a_n743_46660# 0.03492f
C7743 a_11599_46634# a_12549_44172# 0.075725f
C7744 a_n1151_42308# a_n1925_46634# 0.105874f
C7745 a_10227_46804# a_n881_46662# 0.146883f
C7746 a_4791_45118# a_n2661_46634# 0.026643f
C7747 a_3499_42826# a_3681_42891# 0.033957f
C7748 a_n2293_42834# a_n3674_37592# 0.025586f
C7749 a_20447_31679# a_413_45260# 0.226658f
C7750 a_n2293_45010# a_n967_45348# 0.018659f
C7751 a_n2109_45247# en_comp 0.108653f
C7752 a_3357_43084# a_2382_45260# 0.219664f
C7753 a_7499_43078# a_11827_44484# 0.104754f
C7754 a_n357_42282# a_14539_43914# 0.028064f
C7755 a_4646_46812# a_6547_43396# 0.03374f
C7756 a_n1151_42308# a_10355_46116# 0.043227f
C7757 a_4883_46098# a_20202_43084# 0.135688f
C7758 a_5907_46634# a_5257_43370# 0.070316f
C7759 a_n1613_43370# a_765_45546# 0.205521f
C7760 a_2063_45854# a_10903_43370# 0.277624f
C7761 a_4791_45118# a_8199_44636# 0.14611f
C7762 a_n3565_38216# a_n4064_37440# 0.032797f
C7763 a_n3420_37984# a_n3420_37440# 0.132162f
C7764 a_n4064_37984# a_n3565_37414# 0.029309f
C7765 a_1414_42308# a_n784_42308# 0.017857f
C7766 a_413_45260# START 0.035622f
C7767 a_1667_45002# VDD 0.315476f
C7768 a_526_44458# a_3539_42460# 0.213772f
C7769 a_n1925_42282# a_3626_43646# 0.031012f
C7770 a_n2661_45010# a_n2661_42834# 0.01412f
C7771 a_9482_43914# a_13076_44458# 0.103066f
C7772 a_1307_43914# a_5883_43914# 0.289388f
C7773 a_20202_43084# a_5649_42852# 0.011671f
C7774 a_1423_45028# a_4743_44484# 0.022983f
C7775 a_20273_46660# a_12741_44636# 0.540506f
C7776 a_765_45546# a_n2293_46098# 0.054689f
C7777 a_12861_44030# a_11823_42460# 1.2465f
C7778 a_743_42282# a_13291_42460# 0.068071f
C7779 a_n2017_45002# a_n2267_43396# 0.033995f
C7780 a_16979_44734# a_17325_44484# 0.013377f
C7781 a_5205_44484# a_6671_43940# 0.049504f
C7782 a_n357_42282# a_7871_42858# 0.035744f
C7783 a_14537_43396# a_14021_43940# 0.048774f
C7784 a_9313_44734# a_9159_44484# 0.056359f
C7785 a_13259_45724# a_17333_42852# 0.077331f
C7786 a_14275_46494# a_14371_46494# 0.013793f
C7787 a_4419_46090# a_n2661_45546# 0.019708f
C7788 a_n2293_46634# a_2382_45260# 0.046113f
C7789 a_12891_46348# a_9482_43914# 0.314487f
C7790 a_1823_45246# a_n357_42282# 0.031648f
C7791 a_1138_42852# a_n755_45592# 0.062548f
C7792 a_1176_45822# a_997_45618# 0.140567f
C7793 a_17538_32519# VREF_GND 0.117023f
C7794 a_3080_42308# C0_N_btm 0.018211f
C7795 a_n4318_38680# a_n4064_39072# 0.050323f
C7796 a_n356_44636# a_3080_42308# 0.072716f
C7797 a_2959_46660# VDD 0.19762f
C7798 a_4185_45028# a_22485_38105# 0.065539f
C7799 a_n2438_43548# a_n2293_43922# 0.575621f
C7800 a_2711_45572# a_7227_45028# 0.014767f
C7801 a_15227_44166# a_11827_44484# 0.084637f
C7802 a_6945_45028# a_2437_43646# 2.26888f
C7803 a_5907_45546# a_6472_45840# 0.041762f
C7804 a_12549_44172# a_19615_44636# 0.157395f
C7805 a_13661_43548# a_17517_44484# 0.01824f
C7806 a_2063_45854# a_4883_46098# 0.116597f
C7807 a_13381_47204# a_n1435_47204# 0.050056f
C7808 COMP_P a_13258_32519# 0.01028f
C7809 a_14955_43940# a_14955_43396# 0.012141f
C7810 a_19335_46494# VDD 0.198512f
C7811 a_n913_45002# a_2123_42473# 0.029944f
C7812 a_3090_45724# a_10405_44172# 0.126512f
C7813 a_n971_45724# a_n1853_43023# 0.02483f
C7814 a_10903_43370# a_n2661_42834# 0.269313f
C7815 a_11823_42460# a_11787_45002# 0.217891f
C7816 a_13507_46334# a_10341_43396# 0.030637f
C7817 a_4791_45118# a_765_45546# 0.052444f
C7818 a_16327_47482# a_19692_46634# 0.023298f
C7819 a_2107_46812# a_1983_46706# 0.212212f
C7820 a_768_44030# a_5257_43370# 0.028882f
C7821 a_n2438_43548# a_n2661_46098# 0.391488f
C7822 a_5932_42308# C4_N_btm 0.032349f
C7823 a_1169_39043# a_1107_38525# 0.031327f
C7824 a_n4209_38502# a_n3420_38528# 0.230544f
C7825 a_n3565_39304# a_n3420_37984# 0.028129f
C7826 a_n4064_39072# a_n4209_38216# 0.03057f
C7827 a_n3420_39072# a_n3565_38216# 0.030682f
C7828 a_5934_30871# C0_P_btm 0.015126f
C7829 a_1606_42308# VIN_N 0.014401f
C7830 a_n4209_39304# a_n4064_37984# 0.029462f
C7831 a_1666_39587# a_2113_38308# 0.100592f
C7832 a_18783_43370# a_15743_43084# 0.303966f
C7833 a_10341_43396# a_21855_43396# 0.011519f
C7834 a_n2293_43922# a_n1794_35082# 0.019388f
C7835 a_n97_42460# a_18083_42858# 0.010531f
C7836 a_3357_43084# a_5343_44458# 0.02588f
C7837 a_n2017_45002# a_n2267_44484# 0.034473f
C7838 a_n1059_45260# a_n2129_44697# 0.032443f
C7839 a_n2661_45010# a_n1352_44484# 0.051998f
C7840 a_n2810_45028# a_n4318_40392# 0.026026f
C7841 a_14180_45002# a_14309_45348# 0.010132f
C7842 a_n2661_46634# a_6945_45028# 0.03015f
C7843 a_4955_46873# a_5068_46348# 0.081759f
C7844 a_n881_46662# a_8034_45724# 0.020183f
C7845 a_17609_46634# a_17339_46660# 0.010277f
C7846 C10_P_btm C6_P_btm 0.895671f
C7847 C9_P_btm C7_P_btm 0.22201f
C7848 VDAC_P VIN_P 0.255243f
C7849 a_n3674_39768# a_n4334_39616# 0.05081f
C7850 a_n97_42460# a_n1794_35082# 0.035802f
C7851 a_18114_32519# VCM 0.121302f
C7852 a_n699_43396# VDD 0.922998f
C7853 a_13507_46334# a_18727_42674# 0.093566f
C7854 a_n1059_45260# a_15493_43396# 0.044794f
C7855 a_526_44458# a_8605_42826# 0.021896f
C7856 a_7499_43078# a_8147_43396# 0.227361f
C7857 a_3232_43370# a_3499_42826# 0.339727f
C7858 a_1307_43914# a_2889_44172# 0.02756f
C7859 a_13259_45724# a_13678_32519# 0.013938f
C7860 a_17767_44458# a_18248_44752# 0.041822f
C7861 a_13925_46122# a_15015_46420# 0.042415f
C7862 a_13759_46122# a_14840_46494# 0.102325f
C7863 a_14493_46090# a_14275_46494# 0.209641f
C7864 a_13747_46662# a_19431_45546# 0.02276f
C7865 a_n443_46116# a_1307_43914# 0.442637f
C7866 a_1176_45822# a_1337_46116# 0.026848f
C7867 a_n971_45724# a_2809_45028# 0.037351f
C7868 a_22959_43948# VDD 0.297936f
C7869 a_13887_32519# a_4958_30871# 0.030919f
C7870 a_4361_42308# a_18907_42674# 0.010379f
C7871 a_21195_42852# a_21671_42860# 0.177876f
C7872 a_2382_45260# a_743_42282# 0.023665f
C7873 SMPL_ON_N VIN_N 0.525208f
C7874 a_n2956_38680# a_n4318_38216# 0.023189f
C7875 a_n357_42282# a_19987_42826# 0.016903f
C7876 a_13661_43548# a_13720_44458# 0.122691f
C7877 a_n2293_45546# a_n357_42282# 0.032623f
C7878 a_13059_46348# a_6171_45002# 0.070496f
C7879 a_n971_45724# a_n1899_43946# 0.021838f
C7880 a_20820_30879# a_20447_31679# 0.053904f
C7881 a_n2438_43548# a_742_44458# 0.171623f
C7882 a_4883_46098# a_n2661_42834# 0.019268f
C7883 a_n2293_46634# a_5343_44458# 0.026475f
C7884 a_8034_45724# a_8162_45546# 0.14162f
C7885 a_n863_45724# a_n1099_45572# 0.172847f
C7886 a_n971_45724# a_1431_47204# 0.030942f
C7887 a_n237_47217# a_1209_47178# 0.206644f
C7888 a_n1741_47186# a_2952_47436# 0.010669f
C7889 a_n2109_47186# a_3160_47472# 0.054333f
C7890 a_n23_47502# a_327_47204# 0.140943f
C7891 a_1755_42282# a_2123_42473# 0.014573f
C7892 a_14635_42282# a_14113_42308# 0.052122f
C7893 a_1606_42308# a_2351_42308# 0.191324f
C7894 a_13887_32519# VCM 0.011087f
C7895 a_n4318_38680# VDD 0.417422f
C7896 a_22959_46660# VDD 0.299681f
C7897 a_15493_43940# a_19319_43548# 0.36082f
C7898 a_n913_45002# a_8495_42852# 0.030544f
C7899 a_10193_42453# a_11551_42558# 0.228057f
C7900 a_n2956_38216# a_n3565_39590# 0.021271f
C7901 a_13059_46348# a_14673_44172# 0.108306f
C7902 a_n443_42852# a_3065_45002# 0.022494f
C7903 a_5937_45572# a_6298_44484# 0.036004f
C7904 a_8199_44636# a_8103_44636# 0.256009f
C7905 a_15599_45572# a_16333_45814# 0.053479f
C7906 a_15903_45785# a_15765_45572# 0.205788f
C7907 a_6151_47436# a_8492_46660# 0.302615f
C7908 a_768_44030# a_5807_45002# 0.025167f
C7909 a_12549_44172# a_13661_43548# 0.149087f
C7910 COMP_P a_22629_37990# 0.010153f
C7911 a_n2840_43370# a_n2840_42826# 0.026152f
C7912 a_9145_43396# a_10695_43548# 0.053202f
C7913 a_8685_43396# a_14955_43396# 0.111211f
C7914 a_n2810_45028# a_n4209_38502# 0.022376f
C7915 a_n2312_38680# a_n4318_38680# 0.023332f
C7916 a_3537_45260# a_1307_43914# 0.290878f
C7917 a_6171_45002# a_13556_45296# 0.017156f
C7918 a_13249_42308# a_14539_43914# 0.032256f
C7919 a_18143_47464# a_6945_45028# 0.023139f
C7920 a_n881_46662# a_8016_46348# 0.024184f
C7921 a_18597_46090# a_19900_46494# 0.039688f
C7922 a_4883_46098# a_17715_44484# 0.024632f
C7923 a_6755_46942# a_14976_45028# 0.029836f
C7924 a_n4209_38216# VDD 0.839151f
C7925 VDAC_P a_11206_38545# 0.101449f
C7926 a_8912_37509# CAL_N 0.017398f
C7927 a_8037_42858# a_8387_43230# 0.225358f
C7928 a_7871_42858# a_8952_43230# 0.102355f
C7929 a_n2017_45002# a_n2065_43946# 0.045593f
C7930 a_n2293_45010# a_n1899_43946# 0.18948f
C7931 a_n443_42852# a_458_43396# 0.023429f
C7932 a_n2661_44458# a_n2433_44484# 0.039874f
C7933 a_2437_43646# a_895_43940# 0.025092f
C7934 a_13556_45296# a_14673_44172# 0.137701f
C7935 a_16327_47482# a_18175_45572# 0.346603f
C7936 a_14976_45028# a_8049_45260# 0.025611f
C7937 a_n2109_47186# a_413_45260# 0.027314f
C7938 a_584_46384# a_n2661_45010# 0.017317f
C7939 a_11599_46634# a_19431_45546# 0.056971f
C7940 a_167_45260# a_2698_46116# 0.019127f
C7941 a_765_45546# a_6945_45028# 4.99804f
C7942 a_1467_44172# VDD 0.391994f
C7943 a_5534_30871# a_14635_42282# 0.020227f
C7944 a_17517_44484# a_11967_42832# 0.342031f
C7945 a_5111_44636# a_7287_43370# 0.104641f
C7946 a_375_42282# a_458_43396# 0.014454f
C7947 a_10193_42453# a_10341_42308# 0.061874f
C7948 a_n1151_42308# VDD 2.57238f
C7949 a_12861_44030# a_14539_43914# 0.02276f
C7950 a_n2312_40392# a_n4318_40392# 0.025284f
C7951 a_3090_45724# a_3357_43084# 0.546562f
C7952 a_5534_30871# a_n3420_37984# 0.043974f
C7953 a_9672_43914# a_9801_44260# 0.010132f
C7954 a_5343_44458# a_743_42282# 0.010119f
C7955 a_14084_46812# VDD 0.087769f
C7956 a_13059_46348# a_12607_44458# 0.033056f
C7957 a_11823_42460# a_13904_45546# 0.067334f
C7958 a_11599_46634# a_12891_46348# 0.150715f
C7959 a_11453_44696# a_22959_47212# 0.182671f
C7960 a_3160_47472# a_n1925_46634# 0.026425f
C7961 a_14311_47204# a_768_44030# 0.033509f
C7962 a_n1435_47204# a_13675_47204# 0.012767f
C7963 a_n4318_37592# a_n4064_37984# 0.050508f
C7964 a_3626_43646# a_3539_42460# 0.017877f
C7965 a_19240_46482# VDD 0.077608f
C7966 a_10193_42453# a_18494_42460# 0.074751f
C7967 a_22959_45572# a_413_45260# 0.021231f
C7968 a_n2293_45010# en_comp 0.066194f
C7969 a_n1059_45260# a_n745_45366# 0.0613f
C7970 a_4646_46812# a_6765_43638# 0.043651f
C7971 a_n1151_42308# a_9823_46155# 0.061688f
C7972 a_n2293_46634# a_3090_45724# 1.2853f
C7973 a_2063_45854# a_11387_46155# 0.079443f
C7974 a_13507_46334# a_11415_45002# 0.160889f
C7975 a_n971_45724# a_2324_44458# 0.021839f
C7976 a_18214_42558# VDD 0.295211f
C7977 a_3754_39466# a_3754_39134# 0.296258f
C7978 a_n3420_37984# a_n3690_37440# 0.017537f
C7979 a_413_45260# RST_Z 0.199496f
C7980 a_327_44734# VDD 0.667364f
C7981 a_20202_43084# a_13678_32519# 0.027425f
C7982 a_526_44458# a_3626_43646# 0.022127f
C7983 a_20820_30879# a_13467_32519# 0.053319f
C7984 a_13556_45296# a_12607_44458# 0.01896f
C7985 a_n1151_42308# a_n784_42308# 0.154055f
C7986 a_11813_46116# a_12005_46116# 0.038046f
C7987 a_768_44030# a_n755_45592# 0.202175f
C7988 a_20411_46873# a_12741_44636# 0.095741f
C7989 a_21363_46634# a_20202_43084# 0.048242f
C7990 a_14401_32519# a_4958_30871# 0.079459f
C7991 a_13857_44734# VDD 0.18416f
C7992 a_n2017_45002# a_n2129_43609# 0.024338f
C7993 w_10694_33990# CAL_P 0.03776f
C7994 a_n357_42282# a_7227_42852# 0.185359f
C7995 a_18989_43940# a_17517_44484# 0.021791f
C7996 a_1176_45822# a_n755_45592# 0.091892f
C7997 a_1138_42852# a_n357_42282# 0.325445f
C7998 a_14275_46494# a_14180_46482# 0.049827f
C7999 a_4185_45028# a_n2661_45546# 0.047991f
C8000 a_n2293_46634# a_2274_45254# 0.018017f
C8001 a_n1613_43370# a_1307_43914# 0.056988f
C8002 a_n2497_47436# a_n699_43396# 0.355158f
C8003 a_2981_46116# a_526_44458# 0.077706f
C8004 a_12891_46348# a_13348_45260# 0.097519f
C8005 a_768_44030# a_13017_45260# 0.031385f
C8006 a_n1925_46634# a_413_45260# 0.02974f
C8007 a_n1809_43762# VDD 0.142403f
C8008 a_4190_30871# a_n3420_37984# 0.032285f
C8009 a_n3674_39304# a_n4064_39072# 0.539144f
C8010 a_3422_30871# a_15493_43940# 0.014587f
C8011 a_22315_44484# a_22223_43948# 0.012307f
C8012 a_18494_42460# a_16137_43396# 0.115144f
C8013 a_3177_46902# VDD 0.200982f
C8014 a_n2438_43548# a_n2661_43922# 0.06887f
C8015 a_2711_45572# a_6598_45938# 0.011792f
C8016 a_3483_46348# a_7229_43940# 0.03702f
C8017 a_n2293_46098# a_1307_43914# 0.107603f
C8018 a_5907_45546# a_6194_45824# 0.233657f
C8019 a_12549_44172# a_11967_42832# 0.193926f
C8020 a_n2293_46634# a_14815_43914# 0.057388f
C8021 a_6123_31319# a_5742_30871# 0.106954f
C8022 a_8791_42308# a_9223_42460# 0.014257f
C8023 a_n2840_43370# a_n2433_43396# 0.039807f
C8024 a_19553_46090# VDD 0.204238f
C8025 a_n913_45002# a_1755_42282# 0.169955f
C8026 a_17591_47464# a_17609_46634# 0.014668f
C8027 a_383_46660# a_491_47026# 0.057222f
C8028 a_16327_47482# a_19466_46812# 0.203994f
C8029 a_n2438_43548# a_1799_45572# 0.137623f
C8030 a_n743_46660# a_n2661_46098# 0.414618f
C8031 a_5932_42308# C3_N_btm 0.121156f
C8032 a_1606_42308# VIN_P 0.014401f
C8033 a_5742_30871# EN_VIN_BSTR_P 0.644551f
C8034 a_n4209_38502# a_n3690_38528# 0.045251f
C8035 a_5934_30871# C1_P_btm 0.011025f
C8036 a_18525_43370# a_15743_43084# 0.058072f
C8037 a_10341_43396# a_4361_42308# 0.027045f
C8038 a_16759_43396# a_16867_43762# 0.057222f
C8039 a_n2017_45002# a_n2129_44697# 0.033299f
C8040 a_n2661_45010# a_n1177_44458# 0.052759f
C8041 a_n443_42852# a_2479_44172# 0.035023f
C8042 a_15227_44166# a_16823_43084# 0.022136f
C8043 a_5257_43370# a_5111_42852# 0.013892f
C8044 a_n913_45002# a_n2661_44458# 0.024357f
C8045 a_13507_46334# a_13259_45724# 0.023413f
C8046 a_4955_46873# a_4704_46090# 0.109136f
C8047 a_22537_39537# VDD 0.313136f
C8048 C10_P_btm C7_P_btm 1.39624f
C8049 C9_P_btm C8_P_btm 39.4538f
C8050 EN_VIN_BSTR_P C0_dummy_P_btm 0.026355f
C8051 VDAC_N VIN_N 0.256435f
C8052 a_19721_31679# VREF 0.057702f
C8053 a_n4318_39768# a_n4334_39616# 0.084616f
C8054 a_n3674_39768# a_n4209_39590# 0.044895f
C8055 a_4223_44672# VDD 2.99073f
C8056 a_18114_32519# VREF_GND 0.493553f
C8057 a_526_44458# a_8037_42858# 0.01672f
C8058 a_626_44172# a_453_43940# 0.163589f
C8059 a_7499_43078# a_7112_43396# 0.012965f
C8060 a_1307_43914# a_2675_43914# 0.453622f
C8061 a_17767_44458# a_17970_44736# 0.233657f
C8062 a_13759_46122# a_15015_46420# 0.043475f
C8063 a_13925_46122# a_14275_46494# 0.20669f
C8064 a_18285_46348# a_18051_46116# 0.028958f
C8065 a_13747_46662# a_18691_45572# 0.030666f
C8066 a_5807_45002# a_19256_45572# 0.015716f
C8067 a_4791_45118# a_1307_43914# 0.027544f
C8068 a_1208_46090# a_1337_46116# 0.062574f
C8069 a_15493_43940# VDD 1.4617f
C8070 a_5649_42852# a_17303_42282# 0.060649f
C8071 a_21356_42826# a_21671_42860# 0.084365f
C8072 a_9313_44734# a_19862_44208# 0.024263f
C8073 a_n2956_39304# a_n4318_38216# 0.023331f
C8074 a_n357_42282# a_19164_43230# 0.011328f
C8075 a_n2497_47436# a_1467_44172# 0.046456f
C8076 a_n971_45724# a_n1761_44111# 0.084835f
C8077 a_n1079_45724# a_n1099_45572# 0.15766f
C8078 a_n2293_45546# a_310_45028# 0.113595f
C8079 a_15227_44166# a_15415_45028# 0.222342f
C8080 a_2107_46812# a_n2661_44458# 0.02628f
C8081 a_10903_43370# a_8696_44636# 0.031601f
C8082 a_12549_44172# a_18989_43940# 0.016062f
C8083 a_n2497_47436# a_n1151_42308# 0.156942f
C8084 a_n23_47502# a_n785_47204# 0.031198f
C8085 a_n237_47217# a_327_47204# 0.027301f
C8086 a_n971_45724# a_1239_47204# 0.022077f
C8087 a_n1741_47186# a_2553_47502# 0.010566f
C8088 a_n2109_47186# a_2905_45572# 0.124881f
C8089 a_14209_32519# VIN_N 0.043539f
C8090 a_1606_42308# a_2123_42473# 0.011716f
C8091 a_13291_42460# a_14113_42308# 0.025652f
C8092 a_13887_32519# VREF_GND 0.047292f
C8093 a_n3674_39304# VDD 0.587205f
C8094 a_12741_44636# VDD 0.988199f
C8095 a_1414_42308# a_3457_43396# 0.094207f
C8096 a_20820_30879# RST_Z 0.048737f
C8097 a_n2293_43922# a_4361_42308# 0.035634f
C8098 a_19862_44208# a_20974_43370# 0.026213f
C8099 a_10193_42453# a_5742_30871# 0.303452f
C8100 a_2277_45546# a_2274_45254# 0.011988f
C8101 a_19692_46634# a_20679_44626# 0.010957f
C8102 a_10809_44734# a_11827_44484# 0.029958f
C8103 a_15599_45572# a_15765_45572# 0.576512f
C8104 a_6151_47436# a_8667_46634# 0.357581f
C8105 a_n1741_47186# a_12251_46660# 0.011505f
C8106 a_12549_44172# a_5807_45002# 0.675558f
C8107 a_11136_42852# VDD 0.132515f
C8108 a_n4315_30879# a_n4209_39590# 4.31257f
C8109 a_9145_43396# a_9803_43646# 0.055143f
C8110 a_8685_43396# a_15095_43370# 0.064911f
C8111 a_n97_42460# a_4361_42308# 0.15989f
C8112 a_9290_44172# a_11341_43940# 0.040892f
C8113 a_n2312_38680# a_n3674_39304# 0.023501f
C8114 a_6171_45002# a_9482_43914# 0.016128f
C8115 a_18479_47436# a_20708_46348# 0.04299f
C8116 a_10227_46804# a_6945_45028# 0.220094f
C8117 a_n881_46662# a_7920_46348# 0.025724f
C8118 a_12465_44636# a_2324_44458# 0.070016f
C8119 a_18597_46090# a_20075_46420# 0.073857f
C8120 a_4883_46098# a_17583_46090# 0.012469f
C8121 a_6755_46942# a_3090_45724# 0.050558f
C8122 a_768_44030# a_3483_46348# 0.281593f
C8123 a_n743_46660# a_11415_45002# 0.038831f
C8124 a_8912_37509# a_11206_38545# 1.26605f
C8125 a_n4209_38502# VIN_P 0.028427f
C8126 a_n2293_42834# VDD 0.853754f
C8127 a_n2661_42282# a_5932_42308# 0.070536f
C8128 a_8037_42858# a_8605_42826# 0.178024f
C8129 a_7871_42858# a_9127_43156# 0.043633f
C8130 a_n2293_45010# a_n1761_44111# 0.148418f
C8131 a_n2293_42834# a_7640_43914# 0.040893f
C8132 a_4185_45028# a_4520_42826# 0.012305f
C8133 a_9482_43914# a_14673_44172# 0.42967f
C8134 a_4883_46098# a_8696_44636# 0.023202f
C8135 a_16327_47482# a_16147_45260# 0.017922f
C8136 a_3090_45724# a_8049_45260# 1.23904f
C8137 a_167_45260# a_2521_46116# 0.328009f
C8138 a_11599_46634# a_18691_45572# 0.034093f
C8139 a_4361_42308# a_3823_42558# 0.114877f
C8140 a_1115_44172# VDD 0.165092f
C8141 a_5534_30871# a_13291_42460# 0.045073f
C8142 a_14543_43071# a_14635_42282# 0.075815f
C8143 a_17730_32519# VIN_N 0.047591f
C8144 a_17517_44484# a_19006_44850# 0.016181f
C8145 a_5111_44636# a_6547_43396# 0.035842f
C8146 a_3537_45260# a_8791_43396# 0.071369f
C8147 a_18494_42460# a_14021_43940# 0.026241f
C8148 a_3160_47472# VDD 0.256092f
C8149 a_11453_44696# a_n2661_44458# 0.174607f
C8150 a_5257_43370# a_5205_44484# 0.021038f
C8151 a_2324_44458# a_2711_45572# 0.804101f
C8152 a_526_44458# a_n863_45724# 0.801581f
C8153 a_3483_46348# a_11652_45724# 0.035818f
C8154 a_10807_43548# a_11341_43940# 0.049779f
C8155 a_5891_43370# a_10341_43396# 0.087957f
C8156 a_9313_44734# a_14579_43548# 0.038528f
C8157 a_n2840_43914# a_n2840_43370# 0.025171f
C8158 a_6453_43914# a_6671_43940# 0.08213f
C8159 a_13607_46688# VDD 0.209568f
C8160 a_11823_42460# a_13527_45546# 0.027805f
C8161 a_n2293_46634# a_1414_42308# 0.260739f
C8162 a_n746_45260# a_288_46660# 0.010226f
C8163 a_2063_45854# a_n2438_43548# 0.033724f
C8164 a_2905_45572# a_n1925_46634# 0.029452f
C8165 a_13487_47204# a_768_44030# 0.371206f
C8166 a_n1435_47204# a_13569_47204# 0.011393f
C8167 a_16375_45002# VDD 1.14948f
C8168 a_10193_42453# a_18184_42460# 0.216199f
C8169 a_n2472_45002# en_comp 0.117861f
C8170 a_19963_31679# a_413_45260# 0.0432f
C8171 a_n2661_45010# a_n967_45348# 0.019427f
C8172 a_10907_45822# a_n2661_43370# 0.057449f
C8173 a_n1059_45260# a_n913_45002# 1.19505f
C8174 a_4646_46812# a_6197_43396# 0.601282f
C8175 a_20916_46384# a_15227_44166# 0.681561f
C8176 a_2063_45854# a_11133_46155# 0.026232f
C8177 a_n1151_42308# a_9569_46155# 0.05766f
C8178 a_13507_46334# a_20202_43084# 0.205796f
C8179 a_19594_46812# a_19692_46634# 0.134424f
C8180 a_19332_42282# VDD 0.227361f
C8181 a_n4064_39616# EN_VIN_BSTR_P 0.073198f
C8182 a_n4209_38216# a_n4064_37440# 0.028219f
C8183 a_n3565_38216# a_n3420_37440# 0.038559f
C8184 a_n4064_37984# a_n4209_37414# 0.027993f
C8185 a_n3420_37984# a_n3565_37414# 0.032929f
C8186 a_n3690_38304# a_n3690_37440# 0.050585f
C8187 a_413_45260# VDD 1.203f
C8188 a_9290_44172# a_10341_43396# 0.157042f
C8189 a_n1925_42282# a_2982_43646# 0.036209f
C8190 a_1423_45028# a_4223_44672# 0.013079f
C8191 a_9482_43914# a_12607_44458# 0.151452f
C8192 a_3090_45724# a_8953_45546# 0.032771f
C8193 a_4646_46812# a_5066_45546# 0.020397f
C8194 a_768_44030# a_n357_42282# 0.175577f
C8195 a_20107_46660# a_12741_44636# 0.527863f
C8196 a_n743_46660# a_13259_45724# 0.025444f
C8197 a_12861_44030# a_11962_45724# 0.184706f
C8198 a_3080_42308# a_5742_30871# 0.097222f
C8199 a_n97_42460# a_15890_42674# 0.022679f
C8200 a_n357_42282# a_5755_42852# 0.179701f
C8201 a_n2017_45002# a_n2433_43396# 0.035979f
C8202 a_18374_44850# a_17517_44484# 0.019155f
C8203 a_13259_45724# a_17701_42308# 0.137488f
C8204 a_n2497_47436# a_4223_44672# 0.047068f
C8205 a_12891_46348# a_13159_45002# 0.031652f
C8206 a_n746_45260# a_n2129_44697# 0.17701f
C8207 a_n2012_43396# VDD 0.08228f
C8208 a_17538_32519# VIN_N 0.040191f
C8209 a_14401_32519# VREF_GND 0.066097f
C8210 a_n4318_38680# a_n3420_39072# 0.310238f
C8211 a_5891_43370# a_n97_42460# 0.957548f
C8212 a_3422_30871# a_22223_43948# 0.011616f
C8213 a_18184_42460# a_16137_43396# 0.029846f
C8214 a_2609_46660# VDD 0.312974f
C8215 a_n2438_43548# a_n2661_42834# 0.057776f
C8216 a_2711_45572# a_6667_45809# 0.010894f
C8217 a_5164_46348# a_4927_45028# 0.09665f
C8218 a_13661_43548# a_16241_44734# 0.047309f
C8219 a_8685_42308# a_9223_42460# 0.166964f
C8220 a_n2840_43370# a_n4318_39304# 0.158695f
C8221 a_18985_46122# VDD 0.253642f
C8222 a_n913_45002# a_1606_42308# 0.025848f
C8223 a_19237_31679# a_17364_32525# 0.053938f
C8224 a_10807_43548# a_10341_43396# 0.042318f
C8225 a_9290_44172# a_n2293_43922# 0.369185f
C8226 a_4883_46098# a_11813_46116# 0.019696f
C8227 a_601_46902# a_491_47026# 0.097745f
C8228 a_383_46660# a_288_46660# 0.049827f
C8229 a_n743_46660# a_1799_45572# 0.034264f
C8230 a_n1925_46634# a_2443_46660# 0.054751f
C8231 a_5932_42308# C2_N_btm 0.011289f
C8232 a_5742_30871# a_n1057_35014# 0.171668f
C8233 a_n4209_38502# a_n3565_38502# 6.84323f
C8234 a_n3565_39304# a_n3565_38216# 0.02823f
C8235 a_n3420_39072# a_n4209_38216# 0.030577f
C8236 a_5934_30871# C2_P_btm 0.011047f
C8237 a_n4209_39304# a_n3420_37984# 0.029539f
C8238 a_5379_42460# VDD 0.213136f
C8239 a_6123_31319# C0_P_btm 0.018968f
C8240 a_18525_43370# a_18783_43370# 0.22264f
C8241 a_18429_43548# a_15743_43084# 0.053516f
C8242 a_16759_43396# a_16664_43396# 0.049827f
C8243 a_12281_43396# a_743_42282# 0.036414f
C8244 a_16977_43638# a_16867_43762# 0.097745f
C8245 a_n2293_43922# a_n3674_37592# 0.062473f
C8246 a_n2293_45010# a_n2267_44484# 0.0118f
C8247 a_n2661_45010# a_n1917_44484# 0.015623f
C8248 a_1423_45028# a_n2293_42834# 0.033636f
C8249 a_9290_44172# a_n97_42460# 0.351467f
C8250 a_n1059_45260# a_n2661_44458# 0.028647f
C8251 a_n2017_45002# a_n2433_44484# 0.039498f
C8252 a_21588_30879# a_10809_44734# 0.110956f
C8253 a_4651_46660# a_4704_46090# 0.013135f
C8254 a_22889_38993# VDD 0.495671f
C8255 C10_P_btm C8_P_btm 2.07867f
C8256 EN_VIN_BSTR_P C0_P_btm 0.12803f
C8257 a_n4318_39768# a_n4209_39590# 0.105246f
C8258 a_19721_31679# VIN_N 0.028583f
C8259 a_2779_44458# VDD 0.38604f
C8260 a_n97_42460# a_n3674_37592# 0.012074f
C8261 a_11691_44458# a_15433_44458# 0.110923f
C8262 a_526_44458# a_7765_42852# 0.023934f
C8263 a_11827_44484# a_11541_44484# 0.0442f
C8264 a_7499_43078# a_7287_43370# 0.057949f
C8265 a_1307_43914# a_895_43940# 0.754684f
C8266 a_13259_45724# a_4361_42308# 0.054653f
C8267 a_16327_47482# a_21335_42336# 0.081786f
C8268 a_13759_46122# a_14275_46494# 0.105995f
C8269 a_13925_46122# a_14493_46090# 0.17072f
C8270 a_19321_45002# a_18479_45785# 0.114441f
C8271 a_13661_43548# a_18691_45572# 0.020905f
C8272 a_5807_45002# a_19431_45546# 0.01527f
C8273 a_13747_46662# a_18909_45814# 0.025022f
C8274 a_1823_45246# a_n1925_42282# 0.099018f
C8275 a_n2497_47436# a_n2293_42834# 0.010004f
C8276 a_22223_43948# VDD 0.254313f
C8277 a_21356_42826# a_21195_42852# 0.03853f
C8278 a_5649_42852# a_4958_30871# 0.293366f
C8279 a_n2956_38680# a_n3674_38680# 0.023107f
C8280 a_4185_45028# a_5934_30871# 0.060401f
C8281 a_16922_45042# a_2982_43646# 0.010868f
C8282 a_n4318_40392# a_n4318_39304# 0.024428f
C8283 a_n863_45724# a_n452_45724# 0.046903f
C8284 a_n971_45724# a_n2065_43946# 0.016306f
C8285 a_n2497_47436# a_1115_44172# 0.069778f
C8286 a_15227_44166# a_14797_45144# 0.011685f
C8287 a_20820_30879# a_19963_31679# 0.057032f
C8288 a_21076_30879# a_19479_31679# 0.054875f
C8289 a_n2293_46634# a_n699_43396# 0.016884f
C8290 a_n2661_45546# a_n755_45592# 0.14317f
C8291 a_n237_47217# a_n785_47204# 0.018044f
C8292 a_n971_45724# a_1209_47178# 0.034982f
C8293 a_n1741_47186# a_2063_45854# 0.037801f
C8294 a_n2109_47186# a_2952_47436# 0.050821f
C8295 a_n746_45260# a_327_47204# 0.022743f
C8296 a_n13_43084# VDD 0.260551f
C8297 a_1606_42308# a_1755_42282# 0.278431f
C8298 a_13291_42460# a_13657_42558# 0.026223f
C8299 a_11341_43940# a_19319_43548# 0.042701f
C8300 a_20820_30879# VDD 0.744652f
C8301 a_n2956_38216# a_n4209_39590# 0.021267f
C8302 a_10193_42453# a_11323_42473# 0.034215f
C8303 a_3483_46348# a_13720_44458# 0.010665f
C8304 a_1609_45822# a_2274_45254# 0.11737f
C8305 a_n443_42852# a_2382_45260# 0.020006f
C8306 a_5937_45572# a_5343_44458# 0.024374f
C8307 a_15599_45572# a_15903_45785# 0.161702f
C8308 a_6151_47436# a_7927_46660# 0.182356f
C8309 a_7227_47204# a_7411_46660# 0.011806f
C8310 a_2063_45854# a_7832_46660# 0.011867f
C8311 a_12891_46348# a_5807_45002# 0.044188f
C8312 a_n4064_40160# a_n2302_40160# 0.249627f
C8313 a_8685_43396# a_14205_43396# 0.011249f
C8314 a_2982_43646# a_15743_43084# 0.023587f
C8315 en_comp comp_n 0.026386f
C8316 a_413_45260# a_1423_45028# 0.194002f
C8317 a_2324_44458# a_15682_43940# 0.321744f
C8318 a_8270_45546# a_9803_43646# 0.066865f
C8319 a_3065_45002# a_1307_43914# 0.033168f
C8320 a_3232_43370# a_9482_43914# 0.129525f
C8321 a_4883_46098# a_15682_46116# 0.06363f
C8322 a_2063_45854# a_10586_45546# 0.056181f
C8323 a_17591_47464# a_6945_45028# 0.025004f
C8324 a_n881_46662# a_6419_46155# 0.019005f
C8325 a_18597_46090# a_19335_46494# 0.036056f
C8326 a_6545_47178# a_5066_45546# 0.021464f
C8327 a_6755_46942# a_15009_46634# 0.012747f
C8328 a_12549_44172# a_3483_46348# 0.185475f
C8329 VDAC_N a_11206_38545# 0.15219f
C8330 a_8912_37509# VDAC_P 3.15325f
C8331 a_7871_42858# a_8387_43230# 0.106107f
C8332 a_n2661_42282# a_6171_42473# 0.013039f
C8333 a_1568_43370# a_1793_42852# 0.011559f
C8334 a_n2293_45010# a_n2065_43946# 0.023134f
C8335 a_n2840_44458# a_n2433_44484# 0.039807f
C8336 a_n4318_40392# a_n2661_44458# 0.026979f
C8337 a_2437_43646# a_2127_44172# 0.017247f
C8338 a_n1151_42308# a_3357_43084# 0.028306f
C8339 a_3815_47204# a_2437_43646# 0.012198f
C8340 a_768_44030# a_13249_42308# 0.012496f
C8341 a_n2497_47436# a_413_45260# 0.028795f
C8342 a_n746_45260# a_n745_45366# 0.119822f
C8343 a_11415_45002# a_9290_44172# 0.031886f
C8344 a_11599_46634# a_18909_45814# 0.042943f
C8345 a_644_44056# VDD 0.147321f
C8346 a_14543_43071# a_13291_42460# 0.107887f
C8347 a_17517_44484# a_18588_44850# 0.026595f
C8348 a_5111_44636# a_6765_43638# 0.022146f
C8349 a_n1059_45260# a_9145_43396# 0.016142f
C8350 a_5883_43914# a_n2661_42282# 0.107496f
C8351 a_3537_45260# a_8147_43396# 0.088185f
C8352 a_18184_42460# a_14021_43940# 0.029776f
C8353 a_5343_44458# a_8333_44056# 0.092296f
C8354 a_1431_47204# DATA[1] 0.334099f
C8355 a_2905_45572# VDD 1.22598f
C8356 a_19466_46812# a_20528_45572# 0.157758f
C8357 a_10949_43914# a_11341_43940# 0.0383f
C8358 a_14539_43914# a_15743_43084# 0.024623f
C8359 a_18326_43940# a_18451_43940# 0.145292f
C8360 a_12816_46660# VDD 0.293798f
C8361 a_10193_42453# a_20753_42852# 0.082713f
C8362 a_11823_42460# a_13163_45724# 0.038493f
C8363 a_5937_45572# a_8560_45348# 0.045711f
C8364 a_n971_45724# a_n2129_43609# 0.173854f
C8365 a_584_46384# a_n2438_43548# 0.099362f
C8366 a_2063_45854# a_n743_46660# 1.58762f
C8367 SMPL_ON_N a_11453_44696# 0.147722f
C8368 a_22731_47423# a_22959_47212# 0.08444f
C8369 a_n237_47217# a_2107_46812# 0.086093f
C8370 a_13487_47204# a_12549_44172# 0.036506f
C8371 a_12861_44030# a_768_44030# 0.260776f
C8372 a_n1151_42308# a_n2293_46634# 0.02925f
C8373 a_n4318_37592# a_n3420_37984# 0.404896f
C8374 a_n3674_38216# a_n4064_37984# 0.65176f
C8375 a_n1557_42282# a_648_43396# 0.048175f
C8376 a_19319_43548# a_10341_43396# 0.027205f
C8377 a_3540_43646# a_3626_43646# 0.100706f
C8378 a_2982_43646# a_3539_42460# 0.01563f
C8379 a_13059_46348# a_14021_43940# 0.082427f
C8380 a_n2472_45002# a_n2956_37592# 0.152938f
C8381 a_n2661_45010# en_comp 0.10363f
C8382 a_n2017_45002# a_n913_45002# 0.275686f
C8383 SMPL_ON_N a_17364_32525# 0.029237f
C8384 a_n443_42852# a_5343_44458# 0.057128f
C8385 a_4646_46812# a_6293_42852# 0.030189f
C8386 a_2107_46812# a_8270_45546# 0.047835f
C8387 a_2063_45854# a_11189_46129# 0.294233f
C8388 a_5167_46660# a_5263_46660# 0.013793f
C8389 a_n1151_42308# a_9625_46129# 0.046431f
C8390 a_13507_46334# a_22365_46825# 0.033904f
C8391 a_19594_46812# a_19466_46812# 0.100902f
C8392 a_19321_45002# a_19692_46634# 0.040279f
C8393 a_18907_42674# VDD 0.148872f
C8394 a_7754_39632# a_7754_39300# 0.296258f
C8395 a_22959_43396# a_17364_32525# 0.156288f
C8396 a_n37_45144# VDD 0.138f
C8397 a_13017_45260# a_13076_44458# 0.011055f
C8398 a_20202_43084# a_4361_42308# 0.472299f
C8399 a_1423_45028# a_2779_44458# 0.246285f
C8400 a_9482_43914# a_8975_43940# 0.186623f
C8401 a_526_44458# a_2982_43646# 0.048644f
C8402 a_626_44172# a_n699_43396# 0.042617f
C8403 a_11813_46116# a_11387_46155# 0.080527f
C8404 a_2063_45854# a_11136_45572# 0.054713f
C8405 DATA[5] CLK 0.059607f
C8406 a_13213_44734# VDD 0.184239f
C8407 a_5891_43370# a_n2661_43922# 0.042536f
C8408 a_n357_42282# a_5111_42852# 0.011577f
C8409 a_n2840_44458# a_n2840_43914# 0.026152f
C8410 a_18443_44721# a_17517_44484# 0.029904f
C8411 a_13259_45724# a_17595_43084# 0.118887f
C8412 a_22612_30879# a_13258_32519# 0.065697f
C8413 a_n971_45724# a_n2129_44697# 0.017407f
C8414 a_167_45260# a_n863_45724# 0.424358f
C8415 a_5807_45002# a_6431_45366# 0.018543f
C8416 a_13661_43548# a_6171_45002# 0.032575f
C8417 a_n2293_46634# a_327_44734# 0.024588f
C8418 a_13925_46122# a_14180_46482# 0.056391f
C8419 a_3483_46348# a_n2661_45546# 0.163728f
C8420 a_12891_46348# a_13017_45260# 0.210934f
C8421 a_9290_44172# a_13259_45724# 0.272297f
C8422 a_n2497_47436# a_2779_44458# 0.034441f
C8423 a_104_43370# VDD 0.252393f
C8424 a_17701_42308# a_17531_42308# 0.109201f
C8425 a_n3674_39304# a_n3420_39072# 0.065079f
C8426 a_3080_42308# C0_P_btm 0.018211f
C8427 a_2443_46660# VDD 0.413663f
C8428 a_3422_30871# a_11341_43940# 0.030182f
C8429 a_20512_43084# a_19862_44208# 0.023947f
C8430 SMPL_ON_N a_19237_31679# 0.029331f
C8431 a_8270_45546# a_n2661_44458# 0.019483f
C8432 a_2711_45572# a_6511_45714# 0.04109f
C8433 a_5164_46348# a_5111_44636# 0.024532f
C8434 a_3483_46348# a_5205_44484# 0.065176f
C8435 a_3090_45724# a_11691_44458# 0.245063f
C8436 a_13661_43548# a_14673_44172# 0.36897f
C8437 a_22400_42852# a_22485_38105# 0.198011f
C8438 a_8685_42308# a_8791_42308# 0.147376f
C8439 a_19319_43548# a_n97_42460# 0.029676f
C8440 a_18819_46122# VDD 0.453432f
C8441 a_n2017_45002# a_1755_42282# 0.012188f
C8442 a_9290_44172# a_n2661_43922# 0.029391f
C8443 a_11652_45724# a_11787_45002# 0.077604f
C8444 a_10193_42453# a_9482_43914# 0.029531f
C8445 a_33_46660# a_491_47026# 0.027606f
C8446 a_n1925_46634# a_n2661_46098# 0.059432f
C8447 a_n2661_46634# a_3524_46660# 0.0105f
C8448 a_8128_46384# a_8145_46902# 0.012246f
C8449 a_16327_47482# a_15227_44166# 0.239667f
C8450 a_5932_42308# C1_N_btm 0.011049f
C8451 a_n4209_38502# a_n4334_38528# 0.25243f
C8452 a_5934_30871# C3_P_btm 0.011274f
C8453 a_5267_42460# VDD 0.170631f
C8454 a_6123_31319# C1_P_btm 0.011005f
C8455 a_17324_43396# a_15743_43084# 0.050725f
C8456 a_16223_45938# VDD 0.132317f
C8457 a_16409_43396# a_16867_43762# 0.027606f
C8458 a_n97_42460# a_16795_42852# 0.126591f
C8459 a_1823_45246# a_3539_42460# 0.678673f
C8460 a_3357_43084# a_4223_44672# 0.029613f
C8461 a_n2293_45010# a_n2129_44697# 0.021404f
C8462 a_n2661_45010# a_n1699_44726# 0.04137f
C8463 a_n2017_45002# a_n2661_44458# 0.034362f
C8464 a_20916_46384# a_10809_44734# 0.038071f
C8465 a_4646_46812# a_4704_46090# 0.01107f
C8466 a_18597_46090# a_19240_46482# 0.025784f
C8467 a_n743_46660# a_17715_44484# 0.01357f
C8468 a_8128_46384# a_5066_45546# 0.032968f
C8469 a_22613_38993# VDD 0.533489f
C8470 C10_P_btm C9_P_btm 53.3168f
C8471 EN_VIN_BSTR_P C1_P_btm 0.110046f
C8472 a_18114_32519# VIN_N 0.062517f
C8473 a_949_44458# VDD 1.2275f
C8474 a_n97_42460# a_n327_42558# 0.020924f
C8475 a_19700_43370# a_19339_43156# 0.012115f
C8476 a_11691_44458# a_14815_43914# 0.018499f
C8477 a_16979_44734# a_17767_44458# 0.011457f
C8478 a_526_44458# a_7871_42858# 0.031818f
C8479 a_375_42282# a_453_43940# 0.021162f
C8480 a_11823_42460# a_3626_43646# 0.011402f
C8481 a_1307_43914# a_2479_44172# 0.300587f
C8482 a_3537_45260# a_n2661_42282# 0.105917f
C8483 a_13259_45724# a_13467_32519# 0.030863f
C8484 a_13507_46334# a_17303_42282# 1.68549f
C8485 a_13759_46122# a_14493_46090# 0.053479f
C8486 a_3090_45724# a_n443_42852# 0.269331f
C8487 a_19321_45002# a_18175_45572# 0.01259f
C8488 a_19123_46287# a_19240_46482# 0.157972f
C8489 a_13747_46662# a_18341_45572# 0.554429f
C8490 a_1823_45246# a_526_44458# 1.93329f
C8491 a_10903_43370# a_2324_44458# 0.038342f
C8492 a_11341_43940# VDD 1.23655f
C8493 a_20922_43172# a_21195_42852# 0.119168f
C8494 a_13678_32519# a_4958_30871# 0.031033f
C8495 a_n2956_39304# a_n3674_38680# 0.023226f
C8496 a_22959_44484# a_19237_31679# 0.155744f
C8497 SMPL_ON_N EN_OFFSET_CAL 0.066251f
C8498 a_12861_44030# a_17517_44484# 0.069119f
C8499 a_n2497_47436# a_644_44056# 0.016428f
C8500 a_12741_44636# a_3357_43084# 0.036536f
C8501 a_15227_44166# a_14537_43396# 0.105881f
C8502 a_n2661_45546# a_n357_42282# 0.044767f
C8503 a_13887_32519# VIN_N 0.059416f
C8504 a_n237_47217# a_n23_47502# 0.056864f
C8505 a_n746_45260# a_n785_47204# 0.198992f
C8506 a_n971_45724# a_327_47204# 0.075444f
C8507 a_n1741_47186# a_584_46384# 0.021978f
C8508 a_n2109_47186# a_2553_47502# 0.04572f
C8509 a_13678_32519# VCM 0.014539f
C8510 a_n1076_43230# VDD 0.292942f
C8511 a_3422_30871# a_10341_43396# 0.029183f
C8512 a_11967_42832# a_16547_43609# 0.176385f
C8513 a_19862_44208# a_21381_43940# 0.113704f
C8514 a_22591_46660# VDD 0.251892f
C8515 a_10193_42453# a_10723_42308# 0.046812f
C8516 a_21076_30879# C8_N_btm 0.384801f
C8517 a_n2810_45572# a_n3565_39590# 0.020853f
C8518 a_n1741_47186# a_11901_46660# 0.034005f
C8519 a_n1151_42308# a_6755_46942# 0.142929f
C8520 a_6151_47436# a_8145_46902# 0.178565f
C8521 a_11309_47204# a_5807_45002# 0.032739f
C8522 a_14097_32519# EN_VIN_BSTR_N 0.031989f
C8523 COMP_P CAL_P 0.037539f
C8524 a_327_44734# a_626_44172# 0.120093f
C8525 a_2324_44458# a_14955_43940# 0.029449f
C8526 a_3357_43084# a_n2293_42834# 0.045124f
C8527 a_8270_45546# a_9145_43396# 0.02247f
C8528 a_n2442_46660# a_n4318_38680# 0.023781f
C8529 a_6171_45002# a_13159_45002# 0.012283f
C8530 a_4883_46098# a_2324_44458# 0.074521f
C8531 a_18479_47436# a_20075_46420# 0.061108f
C8532 a_n2840_46634# a_n2840_46090# 0.026152f
C8533 a_16588_47582# a_6945_45028# 0.011591f
C8534 a_n1613_43370# a_6419_46155# 0.013016f
C8535 a_n1151_42308# a_8049_45260# 0.075767f
C8536 a_18597_46090# a_19553_46090# 0.021441f
C8537 a_6151_47436# a_5066_45546# 0.019067f
C8538 a_6755_46942# a_14084_46812# 0.052304f
C8539 a_12891_46348# a_3483_46348# 0.053153f
C8540 a_2684_37794# VDD 0.286899f
C8541 VDAC_N VDAC_P 4.74149f
C8542 a_7765_42852# a_8037_42858# 0.309282f
C8543 a_7871_42858# a_8605_42826# 0.06628f
C8544 a_2982_43646# a_21195_42852# 0.034024f
C8545 a_1568_43370# a_1709_42852# 0.015873f
C8546 a_n755_45592# a_n1557_42282# 0.199254f
C8547 a_n2840_44458# a_n2661_44458# 0.179135f
C8548 a_2202_46116# a_167_45260# 0.159883f
C8549 a_3785_47178# a_2437_43646# 0.015875f
C8550 a_12549_44172# a_13249_42308# 0.066967f
C8551 a_n746_45260# a_n913_45002# 0.051081f
C8552 a_11599_46634# a_18341_45572# 0.588263f
C8553 a_175_44278# VDD 0.20887f
C8554 a_5111_44636# a_6197_43396# 0.025934f
C8555 a_3537_45260# a_7112_43396# 0.046531f
C8556 a_10193_42453# a_10796_42968# 0.015009f
C8557 a_1239_47204# DATA[1] 0.01925f
C8558 a_2952_47436# VDD 0.089131f
C8559 a_3483_46348# a_11322_45546# 0.554731f
C8560 a_n2293_46634# a_n2293_42834# 0.027042f
C8561 a_n746_45260# a_556_44484# 0.045671f
C8562 a_10341_43396# VDD 0.401264f
C8563 a_10729_43914# a_11341_43940# 0.243062f
C8564 a_12991_46634# VDD 0.357655f
C8565 a_n755_45592# a_5934_30871# 0.040823f
C8566 a_5663_43940# a_5829_43940# 0.143754f
C8567 a_7499_43078# a_8697_45822# 0.038073f
C8568 a_18597_46090# a_15493_43940# 0.024181f
C8569 a_8199_44636# a_8560_45348# 0.03862f
C8570 a_n1613_43370# a_n2661_42282# 0.017743f
C8571 a_11823_42460# a_12791_45546# 0.030093f
C8572 a_584_46384# a_n743_46660# 0.42078f
C8573 a_22731_47423# a_11453_44696# 0.048111f
C8574 a_13717_47436# a_768_44030# 0.029731f
C8575 a_12861_44030# a_12549_44172# 1.20253f
C8576 a_2982_43646# a_3626_43646# 6.553431f
C8577 a_n2293_46098# a_n2661_42282# 0.182071f
C8578 a_3357_43084# a_413_45260# 7.24598f
C8579 a_n2661_45010# a_n2956_37592# 0.163638f
C8580 a_n2017_45002# a_n1059_45260# 6.27837f
C8581 a_2437_43646# a_2274_45254# 0.01398f
C8582 a_4646_46812# a_6031_43396# 0.849684f
C8583 a_19594_46812# a_19333_46634# 0.060858f
C8584 a_768_44030# a_14035_46660# 0.270355f
C8585 a_12549_44172# a_14180_46812# 0.023435f
C8586 a_2063_45854# a_9290_44172# 0.655982f
C8587 a_n1151_42308# a_8953_45546# 0.120628f
C8588 a_4791_45118# a_6419_46155# 0.371259f
C8589 a_18597_46090# a_12741_44636# 0.267775f
C8590 a_19321_45002# a_19466_46812# 0.130025f
C8591 a_4646_46812# a_7715_46873# 0.058457f
C8592 a_18727_42674# VDD 0.181095f
C8593 a_7174_31319# C0_N_btm 0.050478f
C8594 a_n4064_40160# C10_P_btm 0.460005f
C8595 a_n3420_39616# EN_VIN_BSTR_P 0.068222f
C8596 a_n4209_38216# a_n3420_37440# 0.035706f
C8597 a_2113_38308# VDAC_Ni 0.318652f
C8598 a_n3420_37984# a_n4209_37414# 0.03f
C8599 a_n3565_38216# a_n3565_37414# 0.046412f
C8600 VDAC_Pi a_3754_39134# 0.012307f
C8601 a_14209_32519# a_17364_32525# 0.056697f
C8602 a_n143_45144# VDD 0.092f
C8603 a_12281_43396# a_5534_30871# 0.012136f
C8604 a_20202_43084# a_13467_32519# 0.333168f
C8605 a_1423_45028# a_949_44458# 0.06121f
C8606 a_9482_43914# a_10057_43914# 0.401746f
C8607 a_1307_43914# a_5518_44484# 0.01058f
C8608 a_2711_45572# a_15493_43396# 0.054674f
C8609 a_n1151_42308# a_n961_42308# 0.109068f
C8610 a_3090_45724# a_8199_44636# 0.030057f
C8611 a_11599_46634# a_10193_42453# 0.100544f
C8612 a_n2293_43922# VDD 0.735266f
C8613 a_5891_43370# a_n2661_42834# 0.091553f
C8614 a_18287_44626# a_17517_44484# 0.031756f
C8615 a_21588_30879# a_13258_32519# 0.062822f
C8616 a_10903_43370# a_12839_46116# 0.115226f
C8617 a_5807_45002# a_6171_45002# 0.193427f
C8618 a_n2293_46634# a_413_45260# 0.497204f
C8619 a_13759_46122# a_14180_46482# 0.086708f
C8620 a_n746_45260# a_n2661_44458# 0.079054f
C8621 a_n2497_47436# a_949_44458# 0.127971f
C8622 a_n1853_46287# a_n356_45724# 0.011459f
C8623 a_n97_42460# VDD 3.61113f
C8624 a_19987_42826# a_20256_43172# 0.043356f
C8625 a_17701_42308# a_17303_42282# 0.049097f
C8626 a_14401_32519# VIN_N 0.030351f
C8627 a_n3674_39304# a_n3690_39392# 0.071784f
C8628 a_3080_42308# C1_P_btm 0.011373f
C8629 a_n357_42282# a_16877_42852# 0.016936f
C8630 a_n2661_46098# VDD 0.979859f
C8631 a_4185_45028# a_3232_43370# 0.018743f
C8632 a_2711_45572# a_6472_45840# 0.049759f
C8633 a_5164_46348# a_5147_45002# 0.060833f
C8634 a_3090_45724# a_19113_45348# 0.128103f
C8635 a_2063_45854# a_10807_43548# 0.094631f
C8636 a_n2109_47186# a_2747_46873# 0.087441f
C8637 a_9313_45822# a_11459_47204# 0.210847f
C8638 a_8325_42308# a_8791_42308# 0.173196f
C8639 a_n1794_35082# a_4958_30871# 0.036823f
C8640 a_19237_31679# a_14209_32519# 0.052426f
C8641 a_17730_32519# a_17364_32525# 0.054843f
C8642 a_17957_46116# VDD 0.138777f
C8643 a_n967_45348# a_n1794_35082# 0.03295f
C8644 a_n2017_45002# a_1606_42308# 0.04498f
C8645 a_11322_45546# a_11963_45334# 0.028732f
C8646 a_16375_45002# a_16237_45028# 0.035582f
C8647 a_9290_44172# a_n2661_42834# 0.046011f
C8648 a_n1613_43370# a_7112_43396# 0.245085f
C8649 a_33_46660# a_288_46660# 0.056391f
C8650 a_n1925_46634# a_1799_45572# 0.035794f
C8651 a_8128_46384# a_7577_46660# 0.023306f
C8652 a_10227_46804# a_14976_45028# 0.536884f
C8653 a_1123_46634# a_948_46660# 0.234322f
C8654 a_5932_42308# C0_N_btm 0.015561f
C8655 a_n3565_39304# a_n4209_38216# 0.02863f
C8656 a_5934_30871# C4_P_btm 0.030578f
C8657 a_3823_42558# VDD 0.170296f
C8658 a_n4209_39304# a_n3565_38216# 0.02945f
C8659 a_6123_31319# C2_P_btm 0.01106f
C8660 a_18429_43548# a_18525_43370# 0.419086f
C8661 a_17499_43370# a_15743_43084# 0.049383f
C8662 a_16020_45572# VDD 0.077625f
C8663 a_10341_43396# a_21487_43396# 0.010314f
C8664 a_n2293_43922# a_n784_42308# 1.67292f
C8665 a_n356_44636# a_5932_42308# 0.040714f
C8666 a_16409_43396# a_16664_43396# 0.056391f
C8667 a_n97_42460# a_16414_43172# 0.044625f
C8668 a_1823_45246# a_3626_43646# 0.033967f
C8669 a_n2661_45010# a_n2267_44484# 0.260289f
C8670 a_4185_45028# a_4905_42826# 0.039846f
C8671 a_n443_42852# a_1414_42308# 0.193113f
C8672 a_n2293_45010# a_n2433_44484# 0.016908f
C8673 a_768_44030# a_n1925_42282# 0.145535f
C8674 a_18597_46090# a_16375_45002# 0.105669f
C8675 a_6755_46942# a_12741_44636# 0.131965f
C8676 a_n443_46116# a_n23_45546# 0.118272f
C8677 a_22581_37893# VDD 0.902719f
C8678 EN_VIN_BSTR_P C2_P_btm 0.118072f
C8679 a_15743_43084# a_19164_43230# 0.0353f
C8680 a_742_44458# VDD 1.3845f
C8681 a_526_44458# a_7227_42852# 0.062474f
C8682 a_16327_47482# a_20712_42282# 0.030215f
C8683 a_n443_42852# a_12281_43396# 0.030395f
C8684 a_1307_43914# a_2127_44172# 0.127867f
C8685 a_13759_46122# a_13925_46122# 0.576786f
C8686 a_13661_43548# a_18341_45572# 0.037017f
C8687 a_13747_46662# a_18479_45785# 0.020713f
C8688 a_n743_46660# a_8696_44636# 0.032893f
C8689 a_17339_46660# a_18051_46116# 0.040259f
C8690 a_1138_42852# a_526_44458# 0.039045f
C8691 a_12741_44636# a_8049_45260# 0.037594f
C8692 a_21115_43940# VDD 0.145936f
C8693 a_4361_42308# a_17303_42282# 0.050893f
C8694 a_20922_43172# a_21356_42826# 0.017093f
C8695 a_17730_32519# a_19237_31679# 0.0582f
C8696 a_4185_45028# a_6123_31319# 0.068372f
C8697 a_11415_45002# a_19963_31679# 0.033926f
C8698 a_n2661_45546# a_310_45028# 0.035423f
C8699 a_n2497_47436# a_175_44278# 0.05097f
C8700 a_n1079_45724# a_n863_45724# 0.091159f
C8701 a_n971_45724# a_n785_47204# 0.385455f
C8702 a_n746_45260# a_n23_47502# 0.148631f
C8703 a_n2109_47186# a_2063_45854# 0.045645f
C8704 a_14635_42282# a_14456_42282# 0.172313f
C8705 a_13678_32519# VREF_GND 0.047887f
C8706 a_n901_43156# VDD 0.475947f
C8707 a_11415_45002# VDD 1.84504f
C8708 a_19862_44208# a_19741_43940# 0.038152f
C8709 a_11967_42832# a_16243_43396# 0.269605f
C8710 a_10193_42453# a_10533_42308# 0.101629f
C8711 a_8049_45260# a_n2293_42834# 0.224469f
C8712 a_5257_43370# a_5663_43940# 0.014098f
C8713 a_768_44030# a_3737_43940# 0.038628f
C8714 a_n237_47217# a_8270_45546# 0.552109f
C8715 a_n1151_42308# a_10249_46116# 0.060327f
C8716 a_6151_47436# a_7577_46660# 0.578207f
C8717 a_n4334_40480# a_n4064_40160# 0.43652f
C8718 a_n4315_30879# a_n2302_40160# 0.407166f
C8719 a_12800_43218# VDD 0.078978f
C8720 a_1606_42308# VDAC_N 0.010938f
C8721 a_17538_32519# a_17364_32525# 9.64512f
C8722 a_8685_43396# a_14579_43548# 0.03481f
C8723 a_20974_43370# a_20749_43396# 0.0837f
C8724 a_413_45260# a_626_44172# 0.032584f
C8725 a_13259_45724# a_3422_30871# 0.587088f
C8726 a_6171_45002# a_13017_45260# 0.045098f
C8727 a_2382_45260# a_1307_43914# 0.53878f
C8728 a_n2442_46660# a_n3674_39304# 0.024039f
C8729 a_16327_47482# a_10809_44734# 0.036039f
C8730 a_16763_47508# a_6945_45028# 0.01658f
C8731 a_13507_46334# a_15682_46116# 0.022078f
C8732 a_6755_46942# a_13607_46688# 0.129798f
C8733 a_18597_46090# a_18985_46122# 0.027318f
C8734 a_1107_38525# VDD 0.374783f
C8735 VDAC_N a_8912_37509# 3.43288f
C8736 a_6886_37412# VDAC_P 0.062773f
C8737 a_7871_42858# a_8037_42858# 0.772842f
C8738 a_2437_43646# a_1414_42308# 0.023872f
C8739 a_n357_42282# a_n1557_42282# 0.384406f
C8740 a_n2840_44458# a_n4318_40392# 0.161548f
C8741 a_1823_45246# a_167_45260# 0.155648f
C8742 SMPL_ON_P en_comp 0.034192f
C8743 a_12891_46348# a_13249_42308# 0.166217f
C8744 a_19123_46287# a_18985_46122# 0.215692f
C8745 a_n971_45724# a_n913_45002# 0.101346f
C8746 a_n746_45260# a_n1059_45260# 0.138039f
C8747 a_13661_43548# a_10193_42453# 0.211481f
C8748 a_11599_46634# a_18479_45785# 0.028968f
C8749 a_743_42282# a_5379_42460# 0.013947f
C8750 a_n984_44318# VDD 0.281427f
C8751 a_5111_44636# a_6293_42852# 0.072755f
C8752 a_7499_43078# a_10341_42308# 0.42152f
C8753 a_20193_45348# a_15493_43940# 0.10893f
C8754 a_3537_45260# a_7287_43370# 0.400907f
C8755 a_10193_42453# a_10835_43094# 0.041273f
C8756 a_1209_47178# DATA[1] 0.076054f
C8757 a_9290_44172# a_11554_42852# 0.031758f
C8758 a_2553_47502# VDD 0.150286f
C8759 a_12861_44030# a_13076_44458# 0.01178f
C8760 a_4185_45028# a_10193_42453# 3.16135f
C8761 a_3483_46348# a_10490_45724# 0.207668f
C8762 a_5257_43370# a_3232_43370# 0.022872f
C8763 a_8049_45260# a_16375_45002# 0.026933f
C8764 a_9885_43646# VDD 0.190473f
C8765 a_12251_46660# VDD 0.195617f
C8766 a_19721_31679# a_17364_32525# 0.053872f
C8767 a_19237_31679# a_17538_32519# 0.059552f
C8768 a_5663_43940# a_5745_43940# 0.096132f
C8769 a_18079_43940# a_18326_43940# 0.152347f
C8770 a_12741_44636# a_20193_45348# 0.012699f
C8771 a_11962_45724# a_13163_45724# 0.113317f
C8772 a_8568_45546# a_8697_45822# 0.062574f
C8773 a_n2497_47436# a_n97_42460# 0.026966f
C8774 a_8049_45260# a_413_45260# 0.140877f
C8775 a_12427_45724# a_12791_45546# 0.124682f
C8776 a_n2497_47436# a_n2661_46098# 0.026032f
C8777 a_22731_47423# SMPL_ON_N 0.194951f
C8778 a_n971_45724# a_2107_46812# 0.06261f
C8779 a_2063_45854# a_n1925_46634# 0.064288f
C8780 a_16327_47482# a_n881_46662# 0.195459f
C8781 a_12861_44030# a_12891_46348# 0.053595f
C8782 a_22223_47212# a_11453_44696# 0.057984f
C8783 a_n4318_38216# a_n4064_37984# 0.017009f
C8784 a_n3674_38216# a_n3420_37984# 0.064303f
C8785 a_13259_45724# VDD 2.41738f
C8786 a_5257_43370# a_4905_42826# 0.254437f
C8787 a_19479_31679# a_413_45260# 0.055869f
C8788 a_n2840_45002# a_n2956_37592# 0.035532f
C8789 a_n2293_45010# a_n913_45002# 0.015951f
C8790 SMPL_ON_N a_14209_32519# 0.02932f
C8791 a_n443_42852# a_n699_43396# 0.333516f
C8792 a_4646_46812# a_7411_46660# 0.266058f
C8793 a_19594_46812# a_15227_44166# 0.073663f
C8794 a_12549_44172# a_14035_46660# 0.026143f
C8795 a_768_44030# a_13885_46660# 0.029614f
C8796 a_n1151_42308# a_5937_45572# 0.11638f
C8797 a_4791_45118# a_6165_46155# 0.291653f
C8798 a_11453_44696# a_20731_47026# 0.026307f
C8799 a_18057_42282# VDD 0.130308f
C8800 a_7174_31319# C0_dummy_N_btm 0.029132f
C8801 a_14209_32519# a_22959_43396# 0.015679f
C8802 a_n467_45028# VDD 0.385804f
C8803 a_n913_45002# a_9313_44734# 0.055701f
C8804 a_1423_45028# a_742_44458# 0.019572f
C8805 a_1307_43914# a_5343_44458# 0.02568f
C8806 a_375_42282# a_n699_43396# 0.127058f
C8807 a_2711_45572# a_19328_44172# 0.010017f
C8808 a_n1151_42308# a_n1329_42308# 0.167748f
C8809 a_10227_46804# a_13003_42852# 0.012229f
C8810 a_20623_46660# a_20719_46660# 0.013793f
C8811 a_3681_42891# a_n2293_42282# 0.012859f
C8812 a_n97_42460# a_15764_42576# 0.174403f
C8813 a_n2661_43922# VDD 0.611934f
C8814 a_16112_44458# a_16335_44484# 0.011458f
C8815 a_19721_31679# a_19237_31679# 0.071506f
C8816 a_7640_43914# a_n2661_43922# 0.019048f
C8817 a_18248_44752# a_17517_44484# 0.561898f
C8818 a_5807_45002# a_3232_43370# 0.091049f
C8819 a_n2438_43548# en_comp 0.915368f
C8820 a_1823_45246# a_n863_45724# 0.207189f
C8821 a_n971_45724# a_n2661_44458# 0.051008f
C8822 a_n2497_47436# a_742_44458# 0.153038f
C8823 a_167_45260# a_n2293_45546# 0.681309f
C8824 a_n447_43370# VDD 0.204801f
C8825 a_n3674_39304# a_n3565_39304# 0.128699f
C8826 a_3080_42308# C2_P_btm 0.108823f
C8827 a_3600_43914# a_3499_42826# 0.125876f
C8828 a_1799_45572# VDD 0.381212f
C8829 a_4185_45028# a_22775_42308# 0.023674f
C8830 a_3483_46348# a_6171_45002# 0.153232f
C8831 a_19466_46812# a_19778_44110# 0.116901f
C8832 a_2711_45572# a_6194_45824# 0.013872f
C8833 SMPL_ON_N a_17730_32519# 0.029186f
C8834 a_2107_46812# a_9313_44734# 0.023852f
C8835 a_2063_45854# a_10949_43914# 0.129837f
C8836 a_8325_42308# a_8685_42308# 0.141819f
C8837 a_18189_46348# VDD 0.211855f
C8838 en_comp a_n1794_35082# 2.31448f
C8839 a_3483_46348# a_14673_44172# 0.026455f
C8840 a_11322_45546# a_11787_45002# 0.035999f
C8841 a_20202_43084# a_3422_30871# 0.527141f
C8842 a_n1613_43370# a_7287_43370# 0.337957f
C8843 a_11599_46634# a_19692_46634# 0.069066f
C8844 a_171_46873# a_288_46660# 0.159893f
C8845 a_10227_46804# a_3090_45724# 0.320681f
C8846 a_5934_30871# C5_P_btm 0.139996f
C8847 a_3318_42354# VDD 0.203036f
C8848 a_6123_31319# C3_P_btm 0.011333f
C8849 a_n97_42460# a_15567_42826# 0.040819f
C8850 a_16759_43396# a_15743_43084# 0.033478f
C8851 a_16547_43609# a_16664_43396# 0.161376f
C8852 a_17478_45572# VDD 0.411207f
C8853 a_18494_42460# a_7174_31319# 0.023968f
C8854 a_n2661_45010# a_n2129_44697# 0.18531f
C8855 a_4185_45028# a_3080_42308# 0.030391f
C8856 a_2437_43646# a_n699_43396# 0.037149f
C8857 a_8696_44636# a_5891_43370# 0.084594f
C8858 a_n2293_45010# a_n2661_44458# 0.031066f
C8859 a_10193_42453# a_11967_42832# 0.752992f
C8860 a_3090_45724# a_17339_46660# 0.019979f
C8861 a_14976_45028# a_15312_46660# 0.01024f
C8862 a_20916_46384# a_6945_45028# 0.036695f
C8863 a_768_44030# a_526_44458# 0.341438f
C8864 a_15227_44166# a_16388_46812# 0.02839f
C8865 a_n743_46660# a_15682_46116# 0.051046f
C8866 a_16327_47482# a_19443_46116# 0.012553f
C8867 a_n443_46116# a_n356_45724# 0.113738f
C8868 EN_VIN_BSTR_P C3_P_btm 0.100325f
C8869 a_15743_43084# a_19339_43156# 0.128224f
C8870 a_n452_44636# VDD 0.112149f
C8871 a_n3674_39768# a_n4064_40160# 0.139482f
C8872 a_11691_44458# a_13857_44734# 0.049356f
C8873 a_526_44458# a_5755_42852# 0.054788f
C8874 a_16922_45042# a_17517_44484# 0.020096f
C8875 a_14539_43914# a_16979_44734# 0.132799f
C8876 a_1307_43914# a_453_43940# 0.05952f
C8877 a_626_44172# a_644_44056# 0.126386f
C8878 a_13661_43548# a_18479_45785# 0.087389f
C8879 a_13747_46662# a_18175_45572# 0.03273f
C8880 a_n743_46660# a_16680_45572# 0.011176f
C8881 a_20935_43940# VDD 0.184334f
C8882 a_4361_42308# a_4958_30871# 0.087697f
C8883 a_13467_32519# a_17303_42282# 0.040387f
C8884 a_4190_30871# a_18214_42558# 0.078091f
C8885 a_5883_43914# a_9165_43940# 0.019684f
C8886 a_17730_32519# a_22959_44484# 0.015145f
C8887 a_n2661_42834# a_10949_43914# 0.037251f
C8888 a_12465_44636# CLK 0.795478f
C8889 a_2747_46873# VDD 0.626468f
C8890 a_22223_47212# EN_OFFSET_CAL 0.011048f
C8891 a_3090_45724# a_1307_43914# 2.66267f
C8892 a_n2661_45546# a_n1099_45572# 0.068604f
C8893 a_20820_30879# a_19479_31679# 0.052973f
C8894 a_9290_44172# a_8696_44636# 0.032264f
C8895 a_n2293_45546# a_n863_45724# 0.17075f
C8896 a_11415_45002# a_22591_45572# 0.02488f
C8897 a_n746_45260# a_n237_47217# 0.285294f
C8898 a_n971_45724# a_n23_47502# 0.225828f
C8899 a_n452_47436# a_n785_47204# 0.03755f
C8900 a_n1741_47186# a_1431_47204# 0.014137f
C8901 a_n2109_47186# a_584_46384# 0.352889f
C8902 a_1184_42692# a_2123_42473# 0.107417f
C8903 a_13291_42460# a_14456_42282# 0.015899f
C8904 a_n1641_43230# VDD 0.203991f
C8905 a_7499_43078# a_5742_30871# 0.019993f
C8906 a_n2810_45572# a_n4209_39590# 0.020489f
C8907 a_20202_43084# VDD 0.987622f
C8908 a_11967_42832# a_16137_43396# 0.300696f
C8909 a_2253_43940# a_2455_43940# 0.092725f
C8910 SMPL_ON_N a_17538_32519# 0.029166f
C8911 a_n2293_46634# a_11341_43940# 0.487839f
C8912 a_3090_45724# a_18579_44172# 0.16932f
C8913 a_13661_43548# a_14021_43940# 0.103152f
C8914 a_5937_45572# a_4223_44672# 0.016442f
C8915 a_n1741_47186# a_11735_46660# 0.029236f
C8916 a_6151_47436# a_7715_46873# 0.025823f
C8917 a_6491_46660# a_5257_43370# 0.1719f
C8918 a_n4315_30879# a_n4064_40160# 0.363059f
C8919 a_2711_45572# CLK 0.032985f
C8920 a_327_44734# a_375_42282# 0.067169f
C8921 a_4185_45028# a_14021_43940# 0.038946f
C8922 a_n2438_43548# a_n2157_42858# 0.266513f
C8923 a_4883_46098# a_15015_46420# 0.010147f
C8924 a_13507_46334# a_2324_44458# 0.033576f
C8925 a_n881_46662# a_5204_45822# 0.089827f
C8926 a_6755_46942# a_12816_46660# 0.061031f
C8927 a_18597_46090# a_18819_46122# 0.230891f
C8928 a_6886_37412# a_8912_37509# 0.339465f
C8929 a_5700_37509# VDAC_P 0.081094f
C8930 a_4338_37500# CAL_N 0.052373f
C8931 a_7871_42858# a_7765_42852# 0.379881f
C8932 a_5837_45028# VDD 0.191549f
C8933 a_1423_45028# a_n2661_43922# 0.099477f
C8934 a_2107_46812# a_2711_45572# 0.034922f
C8935 SMPL_ON_P a_n2956_37592# 0.039523f
C8936 a_n1151_42308# a_2437_43646# 0.036608f
C8937 a_12549_44172# a_13527_45546# 0.09647f
C8938 a_19123_46287# a_18819_46122# 0.172712f
C8939 a_1138_42852# a_167_45260# 0.250282f
C8940 a_1823_45246# a_2202_46116# 0.25354f
C8941 a_n971_45724# a_n1059_45260# 0.322275f
C8942 a_11599_46634# a_18175_45572# 0.844188f
C8943 a_743_42282# a_5267_42460# 0.010719f
C8944 a_n809_44244# VDD 0.47719f
C8945 a_5111_44636# a_6031_43396# 0.207345f
C8946 a_20193_45348# a_22223_43948# 0.041425f
C8947 a_3537_45260# a_6547_43396# 0.03331f
C8948 a_4223_44672# a_8333_44056# 0.122173f
C8949 a_2063_45854# VDD 3.60498f
C8950 a_12861_44030# a_12883_44458# 0.041056f
C8951 a_12549_44172# a_16922_45042# 0.803336f
C8952 a_12379_46436# a_12638_46436# 0.093752f
C8953 a_n2497_47436# a_n2661_43922# 0.095407f
C8954 a_3483_46348# a_8746_45002# 0.605995f
C8955 SMPL_ON_N a_19721_31679# 0.029197f
C8956 a_n1925_42282# a_n2661_45546# 0.181908f
C8957 a_14955_43396# VDD 0.401358f
C8958 a_18114_32519# a_17364_32525# 0.053739f
C8959 a_9313_44734# a_9145_43396# 0.021257f
C8960 a_5495_43940# a_5745_43940# 0.014406f
C8961 a_12469_46902# VDD 0.203316f
C8962 a_n755_45592# a_6123_31319# 0.199766f
C8963 a_5164_46348# a_n2661_43370# 0.010428f
C8964 a_5937_45572# a_n2293_42834# 0.097247f
C8965 a_18479_47436# a_15493_43940# 0.05409f
C8966 a_12741_44636# a_11691_44458# 0.81445f
C8967 a_18597_46090# a_11341_43940# 0.033543f
C8968 a_n2497_47436# a_n447_43370# 0.192476f
C8969 a_2711_45572# a_15903_45785# 0.028735f
C8970 a_12427_45724# a_11823_42460# 0.17307f
C8971 a_11962_45724# a_12791_45546# 0.124167f
C8972 a_584_46384# a_n1925_46634# 0.047378f
C8973 a_n1151_42308# a_n2661_46634# 0.832521f
C8974 a_6491_46660# a_5807_45002# 0.01567f
C8975 a_n1435_47204# a_12549_44172# 0.072753f
C8976 a_12465_44636# a_11453_44696# 0.084038f
C8977 a_15890_42674# a_4958_30871# 0.017137f
C8978 a_n3674_38216# a_n3690_38304# 0.071735f
C8979 a_5742_30871# a_7174_31319# 0.34728f
C8980 a_14383_46116# VDD 0.132317f
C8981 a_12549_44172# a_15743_43084# 0.021095f
C8982 a_n2109_45247# a_n2017_45002# 0.193269f
C8983 a_n2840_45002# a_n2810_45028# 0.161831f
C8984 a_n2293_45010# a_n1059_45260# 0.020223f
C8985 a_n2293_46634# a_10341_43396# 2.04894f
C8986 a_18479_47436# a_12741_44636# 0.020666f
C8987 a_4646_46812# a_5257_43370# 0.024804f
C8988 a_19321_45002# a_15227_44166# 0.145462f
C8989 a_12549_44172# a_13885_46660# 0.036345f
C8990 a_n1151_42308# a_8199_44636# 0.161616f
C8991 a_4791_45118# a_5497_46414# 0.056648f
C8992 a_n443_46116# a_5204_45822# 0.020803f
C8993 a_11453_44696# a_20528_46660# 0.016145f
C8994 a_13747_46662# a_19466_46812# 0.869986f
C8995 a_13661_43548# a_19692_46634# 0.093373f
C8996 a_7174_31319# C0_dummy_P_btm 0.029132f
C8997 a_n4315_30879# C10_P_btm 1.5848f
C8998 a_n4209_38216# a_n3565_37414# 0.031622f
C8999 a_n3565_38216# a_n4209_37414# 5.88577f
C9000 a_n4334_38304# a_n4334_37440# 0.050585f
C9001 a_17531_42308# VDD 0.262303f
C9002 a_13887_32519# a_17364_32525# 0.050078f
C9003 a_20447_31679# VCM 0.035344f
C9004 a_n1761_44111# a_n1794_35082# 0.060838f
C9005 a_20202_43084# a_21487_43396# 0.019942f
C9006 a_n443_42852# a_15493_43940# 0.301211f
C9007 a_n1059_45260# a_9313_44734# 0.089245f
C9008 a_9482_43914# a_10334_44484# 0.015932f
C9009 a_18479_45785# a_11967_42832# 0.038105f
C9010 a_1307_43914# a_4743_44484# 0.011512f
C9011 a_9290_44172# a_14205_43396# 0.010382f
C9012 a_10903_43370# a_10695_43548# 0.041719f
C9013 a_2711_45572# a_18451_43940# 0.010207f
C9014 a_n1151_42308# COMP_P 0.034f
C9015 a_3090_45724# a_8016_46348# 0.0122f
C9016 a_11453_44696# a_2711_45572# 0.033654f
C9017 a_n97_42460# a_15486_42560# 0.055334f
C9018 a_n2661_42834# VDD 1.00348f
C9019 a_16112_44458# a_16241_44484# 0.010132f
C9020 a_3357_43084# a_n97_42460# 0.113127f
C9021 a_18114_32519# a_19237_31679# 8.86269f
C9022 a_6109_44484# a_n2661_43922# 0.021636f
C9023 a_7640_43914# a_n2661_42834# 0.030156f
C9024 a_17970_44736# a_17517_44484# 0.075165f
C9025 a_n2293_46098# a_n356_45724# 0.022803f
C9026 a_5807_45002# a_5691_45260# 0.19412f
C9027 a_1138_42852# a_n863_45724# 0.135594f
C9028 a_2324_44458# a_10586_45546# 0.436403f
C9029 a_n1352_43396# VDD 0.288329f
C9030 a_16795_42852# a_17303_42282# 0.010298f
C9031 a_n3674_39304# a_n4334_39392# 0.060327f
C9032 a_3080_42308# C3_P_btm 0.027071f
C9033 a_2998_44172# a_3499_42826# 0.027036f
C9034 a_11967_42832# a_14021_43940# 0.030676f
C9035 a_n356_44636# a_1049_43396# 0.042597f
C9036 a_4185_45028# a_21613_42308# 0.028903f
C9037 a_n2293_46634# a_n2293_43922# 0.02819f
C9038 a_3483_46348# a_3232_43370# 0.220803f
C9039 a_2711_45572# a_5907_45546# 0.01826f
C9040 a_11031_47542# a_9313_45822# 0.063846f
C9041 SMPL_ON_P a_n2312_39304# 0.040801f
C9042 a_5932_42308# a_5742_30871# 1.14154f
C9043 a_17730_32519# a_14209_32519# 0.054558f
C9044 a_15493_43396# a_8685_43396# 0.011009f
C9045 a_17715_44484# VDD 0.526119f
C9046 a_n1059_45260# a_961_42354# 0.07089f
C9047 a_n913_45002# a_1184_42692# 0.031137f
C9048 a_19237_31679# a_13887_32519# 0.052352f
C9049 a_3316_45546# a_n2661_43370# 0.022024f
C9050 a_n443_42852# a_n2293_42834# 1.60683f
C9051 a_18597_46090# a_10341_43396# 0.027979f
C9052 a_n2293_46634# a_n97_42460# 0.108602f
C9053 a_n1613_43370# a_6547_43396# 0.154311f
C9054 a_18691_45572# a_18787_45572# 0.013793f
C9055 a_13249_42308# a_6171_45002# 0.026329f
C9056 a_n2438_43548# a_n2267_43396# 0.120634f
C9057 a_11599_46634# a_19466_46812# 0.453656f
C9058 a_5807_45002# a_4646_46812# 0.032485f
C9059 a_n881_46662# a_7927_46660# 0.017621f
C9060 a_n1151_42308# a_765_45546# 1.7705f
C9061 a_10227_46804# a_15009_46634# 0.02057f
C9062 a_601_46902# a_948_46660# 0.051162f
C9063 a_n2293_46634# a_n2661_46098# 0.022053f
C9064 a_16327_47482# a_16292_46812# 0.027563f
C9065 a_n133_46660# a_288_46660# 0.086708f
C9066 a_8128_46384# a_7411_46660# 0.019875f
C9067 a_n4209_39304# a_n4209_38216# 0.029694f
C9068 a_n2302_39072# a_n2302_38778# 0.050477f
C9069 a_2903_42308# VDD 0.22017f
C9070 a_6123_31319# C4_P_btm 0.132906f
C9071 a_n97_42460# a_5342_30871# 0.068562f
C9072 a_16977_43638# a_15743_43084# 0.042866f
C9073 a_10341_43396# a_743_42282# 0.017833f
C9074 a_16243_43396# a_16664_43396# 0.090164f
C9075 a_15861_45028# VDD 0.690795f
C9076 a_375_42282# a_n2293_42834# 0.027465f
C9077 a_4185_45028# a_4699_43561# 0.010947f
C9078 a_1823_45246# a_2982_43646# 0.022597f
C9079 a_13249_42308# a_14673_44172# 0.026424f
C9080 a_n2661_45010# a_n2433_44484# 0.217176f
C9081 a_20916_46384# a_21137_46414# 0.118131f
C9082 a_19594_46812# a_10809_44734# 0.042242f
C9083 a_3877_44458# a_4185_45028# 0.338483f
C9084 a_n743_46660# a_2324_44458# 0.036195f
C9085 a_22527_39145# VDD 0.626886f
C9086 EN_VIN_BSTR_P C4_P_btm 0.116925f
C9087 a_n1352_44484# VDD 0.276725f
C9088 a_n4318_39768# a_n4064_40160# 0.293052f
C9089 a_n97_42460# a_n473_42460# 0.096579f
C9090 a_1307_43914# a_1414_42308# 0.147738f
C9091 a_526_44458# a_5111_42852# 0.265994f
C9092 a_626_44172# a_175_44278# 0.017096f
C9093 a_16327_47482# a_13258_32519# 0.019817f
C9094 a_12861_44030# a_6171_45002# 0.05507f
C9095 a_13661_43548# a_18175_45572# 0.029369f
C9096 a_5807_45002# a_18479_45785# 0.174313f
C9097 a_13747_46662# a_16147_45260# 0.027471f
C9098 a_13351_46090# a_13759_46122# 0.043782f
C9099 a_20623_43914# VDD 0.258478f
C9100 a_13467_32519# a_4958_30871# 0.031235f
C9101 a_4190_30871# a_19332_42282# 0.154377f
C9102 a_n2661_42834# a_10729_43914# 0.01161f
C9103 a_15227_44166# a_13556_45296# 0.047404f
C9104 a_12861_44030# a_14673_44172# 0.015418f
C9105 a_5066_45546# a_8568_45546# 0.04527f
C9106 a_n2661_45546# a_380_45546# 0.012814f
C9107 a_n2497_47436# a_n809_44244# 0.029871f
C9108 a_n2438_43548# a_n2267_44484# 0.120608f
C9109 a_12741_44636# a_2437_43646# 0.023858f
C9110 a_11415_45002# a_3357_43084# 0.053912f
C9111 a_13678_32519# VIN_N 0.067554f
C9112 a_n815_47178# a_n785_47204# 0.123817f
C9113 a_n971_45724# a_n237_47217# 0.134971f
C9114 a_n1741_47186# a_1239_47204# 0.022889f
C9115 a_n2109_47186# a_2124_47436# 0.037038f
C9116 a_13467_32519# VCM 0.020152f
C9117 a_n1423_42826# VDD 0.211036f
C9118 a_1184_42692# a_1755_42282# 0.016329f
C9119 a_13291_42460# a_13575_42558# 0.074792f
C9120 a_n2293_43922# a_743_42282# 0.034167f
C9121 a_22365_46825# VDD 0.193587f
C9122 a_3483_46348# a_8975_43940# 0.016137f
C9123 a_19692_46634# a_11967_42832# 0.032909f
C9124 a_n2312_39304# a_n2438_43548# 0.052323f
C9125 a_n971_45724# a_8270_45546# 0.251101f
C9126 a_9804_47204# a_5807_45002# 0.039093f
C9127 a_6151_47436# a_7411_46660# 0.330209f
C9128 COMP_P a_22537_39537# 0.03695f
C9129 a_11554_42852# VDD 0.078978f
C9130 a_n4315_30879# a_n4334_40480# 0.253307f
C9131 a_3775_45552# VDD 0.089667f
C9132 a_n97_42460# a_743_42282# 0.107736f
C9133 a_17538_32519# a_14209_32519# 0.051332f
C9134 a_14401_32519# a_17364_32525# 7.49646f
C9135 a_n2956_39768# a_n4318_38680# 0.023624f
C9136 a_6709_45028# a_7705_45326# 0.099282f
C9137 a_413_45260# a_375_42282# 0.112554f
C9138 a_n2438_43548# a_n2472_42826# 0.026866f
C9139 a_6171_45002# a_11787_45002# 0.01986f
C9140 a_n1741_47186# a_12839_46116# 0.113988f
C9141 a_16327_47482# a_6945_45028# 0.111399f
C9142 a_n881_46662# a_5164_46348# 0.03104f
C9143 a_768_44030# a_167_45260# 0.014856f
C9144 a_6755_46942# a_12991_46634# 0.077634f
C9145 a_18597_46090# a_17957_46116# 0.018356f
C9146 a_12465_44636# a_13925_46122# 0.018086f
C9147 a_5088_37509# VDAC_P 1.15441f
C9148 a_5700_37509# a_8912_37509# 15.051701f
C9149 a_8530_39574# CAL_P 0.037066f
C9150 a_6886_37412# VDAC_N 0.067053f
C9151 a_4338_37500# a_11206_38545# 0.072616f
C9152 a_3726_37500# CAL_N 0.036205f
C9153 a_7227_42852# a_7765_42852# 0.118623f
C9154 a_3080_42308# a_n2293_42282# 0.122474f
C9155 a_5093_45028# VDD 0.168437f
C9156 a_3422_30871# a_17303_42282# 0.063198f
C9157 a_n2661_45546# a_3539_42460# 0.091495f
C9158 a_n357_42282# a_4905_42826# 0.026713f
C9159 a_n755_45592# a_3080_42308# 0.237742f
C9160 a_12549_44172# a_13163_45724# 0.172293f
C9161 a_16388_46812# a_10809_44734# 0.013923f
C9162 a_1176_45822# a_167_45260# 0.091673f
C9163 a_11599_46634# a_16147_45260# 0.065926f
C9164 SMPL_ON_P a_n2810_45028# 0.039575f
C9165 a_n971_45724# a_n2017_45002# 0.048447f
C9166 a_n4318_38680# a_n4318_37592# 0.027855f
C9167 a_743_42282# a_3823_42558# 0.015894f
C9168 a_n1549_44318# VDD 0.200608f
C9169 a_12895_43230# a_13003_42852# 0.057222f
C9170 a_n237_47217# DATA[3] 0.0265f
C9171 a_327_47204# DATA[0] 0.353891f
C9172 a_20193_45348# a_11341_43940# 0.21261f
C9173 a_3537_45260# a_6765_43638# 0.025724f
C9174 a_584_46384# VDD 2.50905f
C9175 a_12861_44030# a_12607_44458# 0.020604f
C9176 a_n2497_47436# a_n2661_42834# 0.099608f
C9177 a_3483_46348# a_10193_42453# 0.359034f
C9178 SMPL_ON_N a_18114_32519# 0.02927f
C9179 a_526_44458# a_n2661_45546# 0.071855f
C9180 a_15095_43370# VDD 0.169652f
C9181 a_17730_32519# a_17538_32519# 9.37324f
C9182 a_19237_31679# a_14401_32519# 0.055111f
C9183 a_19721_31679# a_14209_32519# 0.051313f
C9184 a_17973_43940# a_18079_43940# 0.419086f
C9185 a_11901_46660# VDD 0.57548f
C9186 a_8199_44636# a_n2293_42834# 0.048304f
C9187 a_n2438_43548# a_n2065_43946# 0.265458f
C9188 a_18597_46090# a_21115_43940# 0.015966f
C9189 a_n2497_47436# a_n1352_43396# 0.061218f
C9190 a_2711_45572# a_15599_45572# 0.045207f
C9191 a_11962_45724# a_11823_42460# 0.177935f
C9192 a_n746_45260# a_383_46660# 0.011439f
C9193 a_3160_47472# a_n2661_46634# 0.026361f
C9194 a_6545_47178# a_5807_45002# 0.030195f
C9195 a_13381_47204# a_12549_44172# 0.135267f
C9196 a_22223_47212# a_22731_47423# 0.011229f
C9197 a_n3674_37592# a_n4064_38528# 0.019942f
C9198 a_15959_42545# a_4958_30871# 0.043235f
C9199 a_n3674_38216# a_n3565_38216# 0.128699f
C9200 a_2896_43646# a_2982_43646# 0.100706f
C9201 a_3090_45724# a_10651_43940# 0.014051f
C9202 a_2437_43646# a_413_45260# 0.20387f
C9203 SMPL_ON_N a_13887_32519# 0.029238f
C9204 a_n2293_45010# a_n2017_45002# 0.076023f
C9205 a_n2661_45010# a_n913_45002# 0.019536f
C9206 a_18597_46090# a_11415_45002# 0.061694f
C9207 a_3877_44458# a_5257_43370# 0.142219f
C9208 a_13747_46662# a_19333_46634# 0.011849f
C9209 a_5167_46660# a_5275_47026# 0.057222f
C9210 a_n1151_42308# a_8349_46414# 0.095055f
C9211 a_4791_45118# a_5204_45822# 0.053732f
C9212 a_13661_43548# a_19466_46812# 0.011727f
C9213 a_4958_30871# RST_Z 0.087554f
C9214 a_7174_31319# C0_P_btm 0.050478f
C9215 a_13258_32519# C0_N_btm 0.033333f
C9216 a_17303_42282# VDD 0.37938f
C9217 a_22591_43396# a_14209_32519# 0.158752f
C9218 a_3357_43084# a_n2661_43922# 0.031253f
C9219 a_626_44172# a_742_44458# 0.022141f
C9220 a_9482_43914# a_10157_44484# 0.321004f
C9221 a_n1925_42282# a_n1557_42282# 0.013245f
C9222 a_526_44458# a_1427_43646# 0.028942f
C9223 a_1307_43914# a_n699_43396# 0.094953f
C9224 a_n2661_45010# a_556_44484# 0.038106f
C9225 a_768_44030# a_n863_45724# 0.020071f
C9226 a_n2293_46634# a_13259_45724# 0.032341f
C9227 a_n743_46660# a_12839_46116# 0.011568f
C9228 a_n97_42460# a_15051_42282# 0.049661f
C9229 a_17767_44458# a_17517_44484# 0.055175f
C9230 a_n357_42282# a_2905_42968# 0.011153f
C9231 a_6109_44484# a_n2661_42834# 0.026239f
C9232 a_18114_32519# a_22959_44484# 0.016108f
C9233 a_19721_31679# a_17730_32519# 0.051334f
C9234 a_n443_42852# a_n13_43084# 0.13203f
C9235 a_n2293_46098# a_3503_45724# 0.01404f
C9236 a_1823_45246# a_n2293_45546# 0.234971f
C9237 a_n2661_46634# a_413_45260# 0.029743f
C9238 a_6755_46942# a_16020_45572# 0.010518f
C9239 a_12594_46348# a_12638_46436# 0.049443f
C9240 a_n1177_43370# VDD 0.354704f
C9241 a_n3674_39304# a_n4209_39304# 0.059449f
C9242 a_20193_45348# a_10341_43396# 0.086741f
C9243 a_5343_44458# a_8147_43396# 0.014327f
C9244 a_n356_44636# a_1209_43370# 0.025313f
C9245 a_n2293_46634# a_n2661_43922# 0.023539f
C9246 a_12741_44636# a_16751_45260# 0.01378f
C9247 a_2711_45572# a_5263_45724# 0.013854f
C9248 a_n357_42282# a_10193_42453# 0.634772f
C9249 a_3090_45724# a_11827_44484# 0.066595f
C9250 a_10903_43370# a_n913_45002# 0.021559f
C9251 a_9863_47436# a_9313_45822# 0.049145f
C9252 a_n1151_42308# a_10227_46804# 0.458569f
C9253 SMPL_ON_P a_n2312_40392# 4.89949f
C9254 a_6151_47436# a_14955_47212# 0.192081f
C9255 a_8337_42558# a_8325_42308# 0.01416f
C9256 a_17583_46090# VDD 0.23578f
C9257 a_10903_43370# CLK 0.018377f
C9258 a_n1059_45260# a_1184_42692# 0.019924f
C9259 en_comp a_n3674_37592# 0.050998f
C9260 a_7499_43078# a_9482_43914# 0.062333f
C9261 a_n1613_43370# a_6765_43638# 0.164755f
C9262 a_n2438_43548# a_n2129_43609# 0.068602f
C9263 a_n2438_43548# a_288_46660# 0.013776f
C9264 a_4915_47217# a_13059_46348# 0.021189f
C9265 a_n2661_46634# a_2609_46660# 0.045654f
C9266 a_5807_45002# a_3877_44458# 0.034811f
C9267 a_3160_47472# a_765_45546# 0.027219f
C9268 a_33_46660# a_948_46660# 0.117156f
C9269 a_2713_42308# VDD 0.208275f
C9270 a_5932_42308# C0_P_btm 0.015561f
C9271 a_n1794_35082# VIN_N 0.03907f
C9272 a_6123_31319# C5_P_btm 0.022099f
C9273 a_17499_43370# a_18429_43548# 0.012474f
C9274 a_16409_43396# a_15743_43084# 0.586918f
C9275 a_8696_44636# VDD 1.12228f
C9276 a_18494_42460# a_20107_42308# 0.035023f
C9277 a_8953_45546# a_n97_42460# 0.015611f
C9278 a_n2661_45010# a_n2661_44458# 0.090852f
C9279 a_6755_46942# a_11415_45002# 0.02226f
C9280 a_n881_46662# a_5066_45546# 0.801045f
C9281 a_n237_47217# a_2711_45572# 0.025745f
C9282 a_20916_46384# a_20708_46348# 0.189941f
C9283 a_19321_45002# a_10809_44734# 0.035502f
C9284 a_3877_44458# a_3699_46348# 0.084544f
C9285 a_4646_46812# a_3483_46348# 0.048267f
C9286 a_n743_46660# a_14840_46494# 0.010488f
C9287 a_22589_40055# VDD 1.08898f
C9288 EN_VIN_BSTR_P C5_P_btm 0.115337f
C9289 a_19998_34978# a_21753_35474# 0.150805f
C9290 a_n1177_44458# VDD 0.347966f
C9291 a_n357_42282# a_16137_43396# 1.09442f
C9292 a_11691_44458# a_13213_44734# 0.046347f
C9293 a_1307_43914# a_1467_44172# 0.228571f
C9294 a_n1925_42282# a_3935_42891# 0.010366f
C9295 a_526_44458# a_4520_42826# 0.247914f
C9296 a_13259_45724# a_743_42282# 0.066992f
C9297 a_11827_44484# a_14815_43914# 0.029578f
C9298 a_16112_44458# a_14539_43914# 0.13299f
C9299 a_11415_45002# a_8049_45260# 0.426371f
C9300 a_9290_44172# a_2324_44458# 0.026216f
C9301 a_n743_46660# a_16115_45572# 0.012735f
C9302 a_8270_45546# a_2711_45572# 0.063301f
C9303 a_4915_47217# a_13556_45296# 0.146395f
C9304 a_20365_43914# VDD 0.261299f
C9305 a_4190_30871# a_18907_42674# 0.040515f
C9306 a_4883_46098# CLK 0.032195f
C9307 a_19721_31679# a_17538_32519# 0.051191f
C9308 a_22591_44484# a_17730_32519# 0.156987f
C9309 a_n913_45002# a_5649_42852# 0.0586f
C9310 a_n2312_40392# CLK_DATA 0.213071f
C9311 a_15227_44166# a_9482_43914# 0.020073f
C9312 a_14976_45028# a_15415_45028# 0.027906f
C9313 a_5066_45546# a_8162_45546# 0.025437f
C9314 a_n2497_47436# a_n1549_44318# 0.018493f
C9315 a_n2438_43548# a_n2129_44697# 0.060059f
C9316 a_20202_43084# a_3357_43084# 0.029548f
C9317 a_11415_45002# a_19479_31679# 0.224531f
C9318 a_765_45546# a_413_45260# 0.031429f
C9319 a_n971_45724# a_n746_45260# 0.393354f
C9320 a_n452_47436# a_n237_47217# 0.061523f
C9321 a_n1741_47186# a_1209_47178# 0.046323f
C9322 a_n2109_47186# a_1431_47204# 0.050586f
C9323 a_n2497_47436# a_584_46384# 0.06459f
C9324 a_13467_32519# VREF_GND 0.048151f
C9325 a_n1991_42858# VDD 0.575656f
C9326 a_22959_42860# a_22775_42308# 0.019713f
C9327 a_1576_42282# a_1755_42282# 0.168925f
C9328 a_1184_42692# a_1606_42308# 0.125247f
C9329 a_13291_42460# a_13070_42354# 0.155164f
C9330 a_20269_44172# a_19319_43548# 0.12985f
C9331 a_19328_44172# a_19741_43940# 0.04732f
C9332 a_9313_44734# a_14209_32519# 0.068114f
C9333 a_7499_43078# a_10723_42308# 0.029878f
C9334 a_20820_30879# C7_N_btm 0.184297f
C9335 a_3316_45546# a_3537_45260# 0.078381f
C9336 a_n443_42852# a_n37_45144# 0.137227f
C9337 a_16375_45002# a_16751_45260# 0.047561f
C9338 a_2711_45572# a_n2017_45002# 0.02728f
C9339 SMPL_ON_N a_14401_32519# 0.029323f
C9340 a_n1151_42308# a_10467_46802# 0.031981f
C9341 a_8128_46384# a_5807_45002# 0.023925f
C9342 a_4883_46098# a_2107_46812# 2.95673f
C9343 a_7227_45028# VDD 0.501104f
C9344 a_14401_32519# a_22959_43396# 0.016242f
C9345 a_20974_43370# a_14209_32519# 0.049701f
C9346 a_n2956_39768# a_n3674_39304# 0.023853f
C9347 a_7229_43940# a_7705_45326# 0.203098f
C9348 a_3483_46348# a_14021_43940# 0.066924f
C9349 a_n443_46116# a_5066_45546# 0.130975f
C9350 a_11453_44696# a_10903_43370# 0.040346f
C9351 a_16241_47178# a_6945_45028# 0.011279f
C9352 a_15811_47375# a_10809_44734# 0.049971f
C9353 a_22612_30879# a_21076_30879# 0.056101f
C9354 a_n881_46662# a_5068_46348# 0.078135f
C9355 a_6755_46942# a_12251_46660# 0.033714f
C9356 a_12465_44636# a_13759_46122# 0.018063f
C9357 a_n1151_42308# a_8034_45724# 0.040415f
C9358 a_5700_37509# VDAC_N 1.09421f
C9359 a_4338_37500# VDAC_P 0.037246f
C9360 a_5088_37509# a_8912_37509# 16.1906f
C9361 a_n2302_38778# VDD 0.35162f
C9362 a_n4064_39072# VCM 0.035838f
C9363 a_3726_37500# a_11206_38545# 0.11542f
C9364 a_5009_45028# VDD 0.151712f
C9365 a_3422_30871# a_4958_30871# 0.101017f
C9366 a_626_44172# a_n2661_43922# 0.03074f
C9367 a_n2312_40392# a_n1794_35082# 0.033733f
C9368 a_n357_42282# a_3080_42308# 0.023702f
C9369 a_2063_45854# a_3357_43084# 0.023045f
C9370 a_12861_44030# a_18341_45572# 0.026945f
C9371 a_18285_46348# a_17957_46116# 0.12677f
C9372 a_768_44030# a_11823_42460# 0.066425f
C9373 a_12549_44172# a_12791_45546# 0.083854f
C9374 a_6755_46942# a_13259_45724# 0.021651f
C9375 a_4646_46812# a_n357_42282# 0.030404f
C9376 a_n746_45260# a_n2293_45010# 0.023201f
C9377 a_n3674_39304# a_n4318_37592# 0.023516f
C9378 a_743_42282# a_3318_42354# 0.01411f
C9379 a_3422_30871# VCM 1.12142f
C9380 a_5649_42852# a_1755_42282# 0.023826f
C9381 a_n1331_43914# VDD 0.203823f
C9382 a_13113_42826# a_13003_42852# 0.097745f
C9383 a_7499_43078# a_10796_42968# 0.030705f
C9384 a_20193_45348# a_21115_43940# 0.01963f
C9385 a_n356_44636# a_895_43940# 0.026898f
C9386 a_3537_45260# a_6197_43396# 0.337459f
C9387 a_n913_45002# a_8685_43396# 0.03156f
C9388 a_n2312_38680# a_n2302_38778# 0.161815f
C9389 a_n785_47204# DATA[0] 0.598846f
C9390 SMPL_ON_P VIN_P 0.525401f
C9391 a_2124_47436# VDD 0.086403f
C9392 a_8049_45260# a_13259_45724# 0.895805f
C9393 a_19466_46812# a_20273_45572# 0.328586f
C9394 a_5257_43370# a_5111_44636# 0.22597f
C9395 a_3483_46348# a_10180_45724# 0.047643f
C9396 a_4883_46098# a_n2661_44458# 0.019556f
C9397 a_14205_43396# VDD 0.311811f
C9398 a_11813_46116# VDD 0.434656f
C9399 a_18114_32519# a_14209_32519# 0.054602f
C9400 a_17730_32519# a_20974_43370# 0.016457f
C9401 a_n2497_47436# a_n1177_43370# 0.062743f
C9402 a_n2438_43548# a_n2472_43914# 0.032003f
C9403 a_11962_45724# a_12427_45724# 0.064229f
C9404 a_11652_45724# a_11823_42460# 0.035142f
C9405 a_4883_46098# a_11453_44696# 0.071224f
C9406 a_2905_45572# a_n2661_46634# 0.029475f
C9407 a_6151_47436# a_5807_45002# 0.099462f
C9408 a_15803_42450# a_4958_30871# 0.093396f
C9409 a_15959_42545# a_16269_42308# 0.013793f
C9410 a_n3674_38216# a_n4334_38304# 0.059852f
C9411 a_n2293_45010# a_n2109_45247# 0.068458f
C9412 a_n2661_45010# a_n1059_45260# 0.021417f
C9413 a_4185_45028# a_3905_42865# 0.09316f
C9414 a_8696_44636# a_1423_45028# 0.095059f
C9415 a_17339_46660# a_15493_43940# 0.020994f
C9416 a_18597_46090# a_20202_43084# 0.04177f
C9417 a_13661_43548# a_19333_46634# 0.011985f
C9418 a_13747_46662# a_15227_44166# 0.05203f
C9419 a_n881_46662# a_13059_46348# 0.642888f
C9420 a_10227_46804# a_12741_44636# 0.188309f
C9421 a_5385_46902# a_5275_47026# 0.097745f
C9422 a_5907_46634# a_6540_46812# 0.017547f
C9423 a_5167_46660# a_5072_46660# 0.049827f
C9424 a_n1151_42308# a_8016_46348# 0.580516f
C9425 a_4791_45118# a_5164_46348# 0.42219f
C9426 a_11453_44696# a_21188_46660# 0.047802f
C9427 a_5807_45002# a_19466_46812# 0.178376f
C9428 a_n4209_38216# a_n4209_37414# 0.041723f
C9429 VDAC_Pi a_3754_39466# 0.308867f
C9430 a_4958_30871# VDD 1.06745f
C9431 a_15095_43370# a_15567_42826# 0.167909f
C9432 a_13887_32519# a_14209_32519# 0.086073f
C9433 en_comp RST_Z 4.35406f
C9434 a_n967_45348# VDD 0.556063f
C9435 a_19963_31679# VCM 0.035453f
C9436 a_20447_31679# VREF 0.059621f
C9437 a_n443_42852# a_11341_43940# 0.51832f
C9438 a_3357_43084# a_n2661_42834# 0.081135f
C9439 a_10903_43370# a_9145_43396# 0.041756f
C9440 a_9482_43914# a_9838_44484# 0.175591f
C9441 a_526_44458# a_n1557_42282# 0.31675f
C9442 a_8953_45546# a_9885_43646# 0.011162f
C9443 a_1307_43914# a_4223_44672# 0.747516f
C9444 a_20202_43084# a_743_42282# 0.135735f
C9445 a_10227_46804# a_11136_42852# 0.012196f
C9446 a_17339_46660# a_12741_44636# 0.032832f
C9447 VDD VCM 1.50561f
C9448 a_n97_42460# a_14113_42308# 0.356407f
C9449 a_18114_32519# a_17730_32519# 9.15095f
C9450 a_16979_44734# a_17517_44484# 0.109784f
C9451 a_n755_45592# a_1847_42826# 0.053279f
C9452 a_1307_43914# a_15493_43940# 0.057588f
C9453 a_18189_46348# a_8049_45260# 0.030061f
C9454 a_167_45260# a_n2661_45546# 0.084316f
C9455 a_1138_42852# a_n2293_45546# 0.021487f
C9456 a_5807_45002# a_5111_44636# 0.204193f
C9457 a_12594_46348# a_12379_46436# 0.04209f
C9458 a_n1917_43396# VDD 0.204644f
C9459 a_18599_43230# a_18707_42852# 0.057222f
C9460 a_n4318_39768# a_n3674_39768# 3.06574f
C9461 a_18579_44172# a_15493_43940# 0.377126f
C9462 a_2675_43914# a_3499_42826# 0.010775f
C9463 a_n2017_45002# a_18817_42826# 0.018518f
C9464 a_20692_30879# a_14097_32519# 0.051423f
C9465 a_n2293_46634# a_n2661_42834# 0.025484f
C9466 a_8049_45260# a_17478_45572# 0.010438f
C9467 a_2711_45572# a_4099_45572# 0.176427f
C9468 a_10903_43370# a_n1059_45260# 0.028694f
C9469 a_3483_46348# a_4927_45028# 0.032156f
C9470 a_12741_44636# a_1307_43914# 0.05146f
C9471 a_9067_47204# a_9313_45822# 0.013659f
C9472 a_n1920_47178# a_n2312_39304# 0.157528f
C9473 a_6151_47436# a_14311_47204# 0.136645f
C9474 a_5934_30871# a_9223_42460# 0.051891f
C9475 a_n784_42308# a_4958_30871# 0.020733f
C9476 a_17730_32519# a_13887_32519# 0.053953f
C9477 a_n2293_43922# a_5534_30871# 0.271171f
C9478 a_15682_46116# VDD 1.25004f
C9479 a_n2017_45002# a_1184_42692# 0.040166f
C9480 a_n2956_37592# a_n3674_37592# 0.025613f
C9481 a_n2438_43548# a_n2433_43396# 0.415301f
C9482 a_4883_46098# a_9145_43396# 0.02956f
C9483 a_3090_45724# a_n2661_42282# 0.039366f
C9484 a_n1613_43370# a_6197_43396# 0.03252f
C9485 a_13259_45724# a_20193_45348# 0.014145f
C9486 a_8953_45546# a_n2661_43922# 0.024071f
C9487 a_10193_42453# a_11787_45002# 0.0195f
C9488 a_n743_46660# a_288_46660# 0.024827f
C9489 a_n2438_43548# a_1983_46706# 0.057412f
C9490 a_n2661_46634# a_2443_46660# 0.021792f
C9491 a_n881_46662# a_7577_46660# 0.028487f
C9492 a_2905_45572# a_765_45546# 0.039575f
C9493 a_10227_46804# a_13607_46688# 0.027032f
C9494 a_11599_46634# a_15227_44166# 0.101252f
C9495 a_601_46902# a_383_46660# 0.209641f
C9496 a_33_46660# a_1123_46634# 0.041798f
C9497 a_5932_42308# C1_P_btm 0.011049f
C9498 a_n4064_39072# a_n4064_38528# 0.05966f
C9499 a_n1794_35082# VIN_P 0.047209f
C9500 a_n784_42308# VCM 0.195503f
C9501 a_17499_43370# a_17324_43396# 0.234322f
C9502 a_16547_43609# a_15743_43084# 0.028834f
C9503 a_10341_43396# a_4190_30871# 0.090771f
C9504 a_16680_45572# VDD 0.275078f
C9505 a_n97_42460# a_5534_30871# 0.109695f
C9506 a_18494_42460# a_13258_32519# 0.298557f
C9507 a_18184_42460# a_20107_42308# 0.013525f
C9508 a_413_45260# a_22959_45036# 0.024709f
C9509 a_n2956_38216# a_n3674_39768# 0.031697f
C9510 a_2437_43646# a_949_44458# 0.038046f
C9511 a_1307_43914# a_n2293_42834# 0.089964f
C9512 a_n1613_43370# a_5066_45546# 0.015391f
C9513 a_19594_46812# a_6945_45028# 0.014072f
C9514 a_3877_44458# a_3483_46348# 0.083955f
C9515 a_16292_46812# a_16388_46812# 0.318472f
C9516 a_2063_45854# a_2277_45546# 0.057116f
C9517 EN_VIN_BSTR_P C6_P_btm 0.118916f
C9518 a_3422_30871# a_n4064_38528# 0.031148f
C9519 a_n1917_44484# VDD 0.186988f
C9520 a_16327_47482# a_19511_42282# 0.089559f
C9521 a_11691_44458# a_n2293_43922# 0.02314f
C9522 a_1307_43914# a_1115_44172# 0.115939f
C9523 a_526_44458# a_3935_42891# 0.012937f
C9524 a_375_42282# a_175_44278# 0.017991f
C9525 a_n443_42852# a_10341_43396# 0.23026f
C9526 a_1208_46090# a_1431_46436# 0.011458f
C9527 a_n2293_46098# a_5066_45546# 0.140248f
C9528 a_20202_43084# a_8049_45260# 0.042894f
C9529 a_n743_46660# a_16333_45814# 0.014466f
C9530 a_4915_47217# a_9482_43914# 0.269756f
C9531 a_17339_46660# a_16375_45002# 0.0296f
C9532 a_20269_44172# VDD 0.169009f
C9533 a_4190_30871# a_18727_42674# 0.035226f
C9534 a_18114_32519# a_17538_32519# 0.054232f
C9535 a_5883_43914# a_7499_43940# 0.04798f
C9536 a_22485_44484# a_17730_32519# 0.091577f
C9537 a_n913_45002# a_13678_32519# 0.023168f
C9538 a_n1059_45260# a_5649_42852# 0.030637f
C9539 a_14976_45028# a_14797_45144# 0.137651f
C9540 a_11415_45002# a_22223_45572# 0.021019f
C9541 a_n2438_43548# a_n2433_44484# 0.421822f
C9542 a_n2661_45546# a_n863_45724# 0.045552f
C9543 a_n452_47436# a_n746_45260# 0.187792f
C9544 a_n1741_47186# a_327_47204# 0.013765f
C9545 a_n2109_47186# a_1239_47204# 0.080115f
C9546 a_1576_42282# a_1606_42308# 0.176925f
C9547 a_n1853_43023# VDD 0.370563f
C9548 a_7499_43078# a_10533_42308# 0.225871f
C9549 a_n2956_38216# a_n4315_30879# 0.025091f
C9550 a_19862_44208# a_19319_43548# 0.049274f
C9551 a_n443_42852# a_n143_45144# 0.104427f
C9552 a_3090_45724# a_19279_43940# 0.046663f
C9553 a_3316_45546# a_3429_45260# 0.142842f
C9554 a_584_46384# a_3457_43396# 0.120485f
C9555 a_16375_45002# a_1307_43914# 0.101951f
C9556 a_5257_43370# a_3905_42865# 0.106385f
C9557 a_n1151_42308# a_10428_46928# 0.011222f
C9558 a_2063_45854# a_6755_46942# 0.131005f
C9559 a_20974_43370# a_22591_43396# 0.046632f
C9560 a_14401_32519# a_14209_32519# 10.7535f
C9561 a_8685_43396# a_9145_43396# 0.201058f
C9562 a_17538_32519# a_13887_32519# 0.051087f
C9563 a_n97_42460# a_4190_30871# 0.140814f
C9564 a_6598_45938# VDD 0.204705f
C9565 a_7229_43940# a_6709_45028# 0.136786f
C9566 a_15861_45028# a_16237_45028# 0.062212f
C9567 a_413_45260# a_1307_43914# 0.080885f
C9568 a_n443_42852# a_n2293_43922# 0.021367f
C9569 a_n881_46662# a_4704_46090# 0.049125f
C9570 a_4791_45118# a_5066_45546# 0.238282f
C9571 a_768_44030# a_1823_45246# 0.287407f
C9572 a_15673_47210# a_6945_45028# 0.056077f
C9573 a_21588_30879# a_21076_30879# 8.21286f
C9574 a_6755_46942# a_12469_46902# 0.042969f
C9575 a_2063_45854# a_8049_45260# 0.037406f
C9576 a_5700_37509# a_6886_37412# 0.13762f
C9577 a_5088_37509# VDAC_N 0.420254f
C9578 a_3726_37500# VDAC_P 0.059581f
C9579 a_4338_37500# a_8912_37509# 0.331796f
C9580 a_n4064_38528# VDD 1.69554f
C9581 a_n4064_39072# VREF_GND 0.048253f
C9582 a_2809_45028# VDD 0.189682f
C9583 a_1423_45028# a_9159_44484# 0.037664f
C9584 a_626_44172# a_n2661_42834# 0.032386f
C9585 a_n443_42852# a_n97_42460# 0.822111f
C9586 a_18114_32519# a_19721_31679# 0.051894f
C9587 en_comp a_3422_30871# 0.357746f
C9588 a_13249_42308# a_14021_43940# 0.07296f
C9589 a_n2312_39304# a_n3674_37592# 0.026622f
C9590 a_584_46384# a_3357_43084# 0.060446f
C9591 a_n2497_47436# a_n967_45348# 0.021003f
C9592 a_12861_44030# a_18479_45785# 0.058482f
C9593 a_1799_45572# a_1609_45822# 0.079527f
C9594 a_18285_46348# a_18189_46348# 0.118603f
C9595 a_12549_44172# a_11823_42460# 0.624462f
C9596 a_12891_46348# a_12791_45546# 0.012918f
C9597 a_n971_45724# a_n2293_45010# 0.549225f
C9598 a_743_42282# a_2903_42308# 0.010301f
C9599 a_3422_30871# VREF_GND 0.10463f
C9600 a_n4318_38680# a_n3674_38216# 0.023866f
C9601 a_12545_42858# a_13003_42852# 0.027606f
C9602 a_n1899_43946# VDD 0.475205f
C9603 a_7499_43078# a_10835_43094# 0.028158f
C9604 a_375_42282# a_n97_42460# 0.039466f
C9605 a_20193_45348# a_20935_43940# 0.016238f
C9606 a_3537_45260# a_6293_42852# 0.01772f
C9607 a_n1059_45260# a_8685_43396# 0.036086f
C9608 a_n2312_38680# a_n4064_38528# 0.22404f
C9609 a_n971_45724# DATA[3] 0.09508f
C9610 a_n23_47502# DATA[0] 0.022435f
C9611 a_n237_47217# DATA[1] 0.139838f
C9612 a_1431_47204# VDD 0.423871f
C9613 a_19466_46812# a_20107_45572# 0.283769f
C9614 a_5257_43370# a_5147_45002# 0.836149f
C9615 a_14358_43442# VDD 0.170277f
C9616 a_17737_43940# a_17973_43940# 0.22264f
C9617 a_n2956_38680# a_n3565_39590# 0.021577f
C9618 a_11735_46660# VDD 0.407307f
C9619 a_19721_31679# a_13887_32519# 0.051264f
C9620 a_17730_32519# a_14401_32519# 0.086728f
C9621 a_14539_43914# a_16759_43396# 0.012597f
C9622 a_5013_44260# a_5025_43940# 0.011829f
C9623 a_n2497_47436# a_n1917_43396# 0.012526f
C9624 SMPL_ON_P a_n4318_39304# 0.039268f
C9625 a_12861_44030# a_14021_43940# 0.035798f
C9626 a_n1925_42282# a_3232_43370# 0.021554f
C9627 a_20202_43084# a_20193_45348# 0.116706f
C9628 a_11415_45002# a_11691_44458# 0.047412f
C9629 a_584_46384# a_n2293_46634# 0.374996f
C9630 a_4915_47217# a_13747_46662# 0.710704f
C9631 a_12465_44636# a_22223_47212# 0.175138f
C9632 a_n746_45260# a_33_46660# 0.035747f
C9633 a_n3674_37592# a_n3420_38528# 0.020112f
C9634 a_15764_42576# a_4958_30871# 0.413236f
C9635 a_n3674_38216# a_n4209_38216# 0.059407f
C9636 a_21115_43940# a_4190_30871# 0.01145f
C9637 a_n2661_45010# a_n2017_45002# 0.087596f
C9638 a_n443_42852# a_742_44458# 0.168627f
C9639 a_10193_42453# a_17023_45118# 0.027968f
C9640 a_n443_46116# a_4704_46090# 0.017894f
C9641 a_13661_43548# a_15227_44166# 0.805606f
C9642 a_18479_47436# a_11415_45002# 0.033153f
C9643 a_5907_46634# a_5732_46660# 0.233657f
C9644 a_4817_46660# a_5275_47026# 0.031068f
C9645 a_n1151_42308# a_7920_46348# 0.085186f
C9646 a_11453_44696# a_21363_46634# 0.027075f
C9647 a_15095_43370# a_5342_30871# 0.238762f
C9648 a_13678_32519# a_17364_32525# 0.050075f
C9649 a_20447_31679# VIN_N 0.028298f
C9650 en_comp VDD 4.30454f
C9651 a_1307_43914# a_2779_44458# 0.332183f
C9652 a_2711_45572# a_17973_43940# 0.011171f
C9653 a_9290_44172# a_13667_43396# 0.136018f
C9654 VDD VREF_GND 0.482759f
C9655 a_3626_43646# a_5934_30871# 0.192998f
C9656 a_n97_42460# a_13657_42558# 0.011259f
C9657 a_10617_44484# VDD 0.141193f
C9658 a_18114_32519# a_22591_44484# 0.018563f
C9659 a_16979_44734# a_17061_44734# 0.171361f
C9660 a_13259_45724# a_5534_30871# 0.032063f
C9661 a_2437_43646# a_n97_42460# 0.201806f
C9662 a_n357_42282# a_1847_42826# 0.037548f
C9663 a_n443_42852# a_n901_43156# 0.367747f
C9664 a_n2312_39304# a_n2302_39072# 0.130454f
C9665 a_n2497_47436# a_n1917_44484# 0.011319f
C9666 a_17715_44484# a_8049_45260# 0.03139f
C9667 a_12005_46116# a_12379_46436# 0.038694f
C9668 a_n2661_46098# a_2437_43646# 0.025093f
C9669 a_6945_45028# a_5066_45546# 0.018752f
C9670 a_376_46348# a_380_45546# 0.011689f
C9671 a_6755_46942# a_15861_45028# 0.033041f
C9672 a_5807_45002# a_5147_45002# 0.035651f
C9673 a_n1699_43638# VDD 0.210236f
C9674 a_3422_30871# a_19862_44208# 0.030442f
C9675 a_n2017_45002# a_18249_42858# 0.545311f
C9676 a_n1059_45260# a_17333_42852# 0.270324f
C9677 a_20205_31679# a_14097_32519# 0.051224f
C9678 a_4185_45028# a_7174_31319# 0.027406f
C9679 a_n2438_43548# a_556_44484# 0.011144f
C9680 a_15227_44166# a_18587_45118# 0.040339f
C9681 a_4185_45028# a_4558_45348# 0.059418f
C9682 a_10903_43370# a_n2017_45002# 0.029479f
C9683 a_3483_46348# a_5111_44636# 0.340106f
C9684 a_6151_47436# a_13487_47204# 0.038134f
C9685 a_6575_47204# a_9313_45822# 0.017088f
C9686 a_n2109_47186# a_n2312_39304# 0.06316f
C9687 a_4915_47217# a_11599_46634# 0.015066f
C9688 a_n237_47217# a_4883_46098# 0.181672f
C9689 a_8515_42308# a_8685_42308# 0.108744f
C9690 a_5934_30871# a_8791_42308# 0.223675f
C9691 a_22400_42852# a_21613_42308# 0.02387f
C9692 a_14401_32519# a_17538_32519# 0.052152f
C9693 a_22485_44484# a_22591_43396# 0.025074f
C9694 a_19237_31679# a_13678_32519# 0.052466f
C9695 a_2324_44458# VDD 2.73366f
C9696 en_comp a_n784_42308# 0.025103f
C9697 a_n2810_45028# a_n3674_37592# 0.025732f
C9698 a_13259_45724# a_11691_44458# 0.337184f
C9699 a_8953_45546# a_n2661_42834# 0.019463f
C9700 a_5937_45572# a_n2661_43922# 0.048264f
C9701 a_4883_46098# a_8270_45546# 0.278829f
C9702 a_15811_47375# a_16292_46812# 0.080078f
C9703 a_n2438_43548# a_2107_46812# 0.111283f
C9704 a_n133_46660# a_948_46660# 0.102355f
C9705 a_n881_46662# a_7715_46873# 0.02091f
C9706 a_10227_46804# a_12816_46660# 0.253017f
C9707 a_11599_46634# a_18834_46812# 0.012948f
C9708 a_33_46660# a_383_46660# 0.20669f
C9709 a_12861_44030# a_19692_46634# 0.097215f
C9710 a_n2661_46634# a_n2661_46098# 0.066513f
C9711 a_5932_42308# C2_P_btm 0.011289f
C9712 a_n4064_39616# a_n4064_37984# 0.048968f
C9713 a_4958_30871# a_n4064_37440# 0.031235f
C9714 a_n784_42308# VREF_GND 0.068593f
C9715 a_16243_43396# a_15743_43084# 0.600668f
C9716 a_n2293_43922# COMP_P 0.151768f
C9717 a_16855_45546# VDD 0.339227f
C9718 a_11967_42832# a_18504_43218# 0.015494f
C9719 a_18494_42460# a_19647_42308# 0.030348f
C9720 a_18184_42460# a_13258_32519# 0.038977f
C9721 a_18479_45785# a_18287_44626# 0.024431f
C9722 a_n2956_38216# a_n4318_39768# 0.045702f
C9723 a_2437_43646# a_742_44458# 0.081793f
C9724 a_n971_45724# a_2711_45572# 0.214535f
C9725 a_19321_45002# a_6945_45028# 0.042647f
C9726 a_13747_46662# a_10809_44734# 0.045104f
C9727 a_n443_46116# a_2957_45546# 0.020365f
C9728 a_2063_45854# a_1609_45822# 0.035351f
C9729 a_22537_40625# VDD 0.534319f
C9730 a_n4064_37440# VCM 0.020152f
C9731 a_19250_34978# a_19998_34978# 0.08192f
C9732 EN_VIN_BSTR_P C7_P_btm 0.115875f
C9733 a_n1699_44726# VDD 0.198612f
C9734 a_11691_44458# a_n2661_43922# 0.038882f
C9735 a_13259_45724# a_4190_30871# 0.271537f
C9736 a_1208_46090# a_1337_46436# 0.010132f
C9737 a_n743_46660# a_15765_45572# 0.026376f
C9738 a_13507_46334# a_n913_45002# 0.023897f
C9739 a_584_46384# a_626_44172# 0.450256f
C9740 a_19862_44208# VDD 0.588967f
C9741 a_4190_30871# a_18057_42282# 0.02374f
C9742 a_743_42282# a_17303_42282# 0.034786f
C9743 a_19339_43156# a_19987_42826# 0.016188f
C9744 a_22485_44484# a_22591_44484# 0.15878f
C9745 a_5883_43914# a_6671_43940# 0.051304f
C9746 a_19721_31679# a_14401_32519# 0.053967f
C9747 a_n2017_45002# a_5649_42852# 0.03149f
C9748 a_4185_45028# a_5932_42308# 0.118319f
C9749 a_14976_45028# a_14537_43396# 0.087031f
C9750 a_11415_45002# a_2437_43646# 0.01065f
C9751 a_12549_44172# a_14539_43914# 0.110516f
C9752 a_13259_45724# a_n443_42852# 0.022577f
C9753 a_n2472_45546# a_n2293_45546# 0.171197f
C9754 a_n2497_47436# a_n1899_43946# 0.040963f
C9755 a_n2438_43548# a_n2661_44458# 0.136664f
C9756 a_n452_47436# a_n971_45724# 0.330438f
C9757 a_n1741_47186# a_n785_47204# 0.026399f
C9758 a_n2109_47186# a_1209_47178# 0.226908f
C9759 a_13467_32519# VIN_N 0.075801f
C9760 a_n2157_42858# VDD 0.424058f
C9761 a_1241_43940# a_1443_43940# 0.092725f
C9762 a_9313_44734# a_13887_32519# 0.191376f
C9763 a_10193_42453# a_9803_42558# 0.20198f
C9764 a_11967_42832# a_15781_43660# 0.026392f
C9765 a_15227_44166# a_11967_42832# 0.132673f
C9766 a_3316_45546# a_3065_45002# 0.141454f
C9767 a_n357_42282# a_5111_44636# 0.033023f
C9768 a_16375_45002# a_16019_45002# 0.032313f
C9769 a_n881_46662# a_13747_46662# 0.550574f
C9770 a_n2312_39304# a_n1925_46634# 0.071018f
C9771 a_2063_45854# a_10249_46116# 0.078073f
C9772 a_4958_30871# a_n3420_39072# 0.079459f
C9773 a_14401_32519# a_22591_43396# 0.01561f
C9774 a_20974_43370# a_13887_32519# 0.033282f
C9775 a_6667_45809# VDD 0.195842f
C9776 a_n2956_37592# a_n4064_39072# 0.010695f
C9777 a_7276_45260# a_6709_45028# 0.215102f
C9778 a_2711_45572# a_9313_44734# 0.036278f
C9779 a_n443_42852# a_n2661_43922# 0.045456f
C9780 a_16147_45260# a_17719_45144# 0.049848f
C9781 a_6171_45002# a_8953_45002# 0.034987f
C9782 a_6755_46942# a_11901_46660# 0.587021f
C9783 a_n881_46662# a_4419_46090# 0.045203f
C9784 a_4883_46098# a_13759_46122# 0.044004f
C9785 a_16327_47482# a_19900_46494# 0.216811f
C9786 a_n2661_46098# a_765_45546# 0.0407f
C9787 a_15811_47375# a_6945_45028# 0.037131f
C9788 a_n2661_46634# a_11415_45002# 0.494836f
C9789 a_768_44030# a_1138_42852# 0.021091f
C9790 a_11599_46634# a_10809_44734# 0.06157f
C9791 a_5088_37509# a_6886_37412# 0.136505f
C9792 a_4338_37500# VDAC_N 0.046178f
C9793 a_3726_37500# a_8912_37509# 0.267651f
C9794 a_n2946_38778# VDD 0.383009f
C9795 a_375_42282# a_n2661_43922# 0.024229f
C9796 a_n863_45724# a_n1557_42282# 0.034373f
C9797 a_14537_43396# a_15433_44458# 0.018743f
C9798 a_n2312_40392# a_n3674_37592# 0.035844f
C9799 a_1176_45822# a_1138_42852# 0.41217f
C9800 a_12861_44030# a_18175_45572# 0.031037f
C9801 a_n1925_46634# a_6511_45714# 0.028817f
C9802 a_12549_44172# a_12427_45724# 0.152925f
C9803 a_12891_46348# a_11823_42460# 0.033376f
C9804 a_765_45546# a_17957_46116# 0.133328f
C9805 a_n746_45260# a_n2661_45010# 0.400342f
C9806 a_743_42282# a_2713_42308# 0.024879f
C9807 a_n3674_39304# a_n3674_38216# 0.023464f
C9808 a_n1761_44111# VDD 0.620042f
C9809 a_18479_45785# a_19268_43646# 0.12682f
C9810 a_n2312_38680# a_n2946_38778# 0.024631f
C9811 a_n971_45724# DATA[2] 0.099284f
C9812 a_n1741_47186# CLK 0.028114f
C9813 a_7499_43078# a_10518_42984# 0.03265f
C9814 a_n237_47217# DATA[0] 0.040942f
C9815 a_20193_45348# a_20623_43914# 0.048456f
C9816 a_3537_45260# a_6031_43396# 0.034593f
C9817 a_1239_47204# VDD 0.278979f
C9818 a_11827_44484# a_15493_43940# 0.010315f
C9819 a_3483_46348# a_9049_44484# 0.117501f
C9820 a_14579_43548# VDD 0.278225f
C9821 a_18114_32519# a_13887_32519# 0.054996f
C9822 a_14539_43914# a_16977_43638# 0.013865f
C9823 a_22485_44484# a_20974_43370# 0.101193f
C9824 a_13259_45724# a_13657_42558# 0.023664f
C9825 a_n2956_39304# a_n3565_39590# 0.072956f
C9826 a_11186_47026# VDD 0.077608f
C9827 a_n2497_47436# a_n1699_43638# 0.038204f
C9828 a_5937_45572# a_5837_45028# 0.043505f
C9829 a_18479_47436# a_20935_43940# 0.207572f
C9830 a_11322_45546# a_11823_42460# 0.133185f
C9831 a_2324_44458# a_1423_45028# 0.154419f
C9832 a_4185_45028# a_n2661_43370# 0.053994f
C9833 a_10227_46804# a_11341_43940# 0.057378f
C9834 a_526_44458# a_3232_43370# 0.461444f
C9835 a_11415_45002# a_19113_45348# 0.012208f
C9836 a_12741_44636# a_11827_44484# 0.305294f
C9837 a_11459_47204# a_11309_47204# 0.183357f
C9838 a_11599_46634# a_n881_46662# 0.100714f
C9839 a_13507_46334# a_11453_44696# 0.060476f
C9840 a_21811_47423# a_22223_47212# 0.031065f
C9841 a_n746_45260# a_171_46873# 0.120194f
C9842 a_n4318_38216# a_n4334_38304# 0.081663f
C9843 a_10586_45546# CLK 0.125859f
C9844 a_12839_46116# VDD 0.347766f
C9845 SMPL_ON_N a_13678_32519# 0.029315f
C9846 a_n2472_45002# a_n2293_45010# 0.177252f
C9847 a_n2661_45010# a_n2109_45247# 0.025907f
C9848 a_10193_42453# a_16922_45042# 0.035103f
C9849 a_17339_46660# a_11341_43940# 0.023304f
C9850 a_n443_46116# a_4419_46090# 0.20069f
C9851 a_5807_45002# a_15227_44166# 0.042586f
C9852 a_13661_43548# a_18834_46812# 0.1407f
C9853 a_18479_47436# a_20202_43084# 0.040227f
C9854 a_4817_46660# a_5072_46660# 0.06121f
C9855 a_2063_45854# a_5937_45572# 0.012248f
C9856 a_n1151_42308# a_6419_46155# 0.028969f
C9857 a_n2497_47436# a_2324_44458# 0.796031f
C9858 a_11453_44696# a_20623_46660# 0.029618f
C9859 a_7754_39964# a_7754_39632# 0.296522f
C9860 a_n4064_38528# a_n4064_37440# 0.045121f
C9861 a_12281_43396# a_12545_42858# 0.029151f
C9862 a_19963_31679# VREF 0.055795f
C9863 a_n1761_44111# a_n784_42308# 0.034368f
C9864 a_15095_43370# a_15279_43071# 0.105784f
C9865 a_n2956_37592# VDD 1.25966f
C9866 a_1307_43914# a_949_44458# 0.028157f
C9867 a_2437_43646# a_n2661_43922# 0.033401f
C9868 a_9290_44172# a_10695_43548# 0.011352f
C9869 a_n1925_42282# a_3080_42308# 0.897997f
C9870 a_526_44458# a_4905_42826# 0.202895f
C9871 a_12465_44636# a_2711_45572# 0.027219f
C9872 VDD VREF 4.8299f
C9873 C10_N_btm VCM 10.5945f
C9874 a_15743_43084# a_15597_42852# 0.055955f
C9875 a_18114_32519# a_22485_44484# 0.020813f
C9876 a_14539_43914# a_17061_44734# 0.020462f
C9877 a_10193_42453# a_15743_43084# 0.027326f
C9878 a_1307_43914# a_11341_43940# 2.31482f
C9879 a_n2312_39304# a_n4064_39072# 0.094407f
C9880 a_n2497_47436# a_n1699_44726# 0.012807f
C9881 a_22612_30879# a_413_45260# 0.11791f
C9882 a_768_44030# a_7229_43940# 0.042486f
C9883 a_15227_44166# a_15143_45578# 0.010748f
C9884 a_n2312_38680# a_n2956_37592# 0.048307f
C9885 a_6755_46942# a_8696_44636# 0.04097f
C9886 a_1823_45246# a_n2661_45546# 0.181403f
C9887 SMPL_ON_P a_n4318_40392# 0.039594f
C9888 a_n2267_43396# VDD 0.570924f
C9889 a_5342_30871# a_4958_30871# 10.9366f
C9890 a_18579_44172# a_11341_43940# 0.030765f
C9891 a_n1059_45260# a_18083_42858# 0.021784f
C9892 a_n2017_45002# a_17333_42852# 0.314084f
C9893 a_n743_46660# CLK 0.028835f
C9894 a_491_47026# VDD 0.132552f
C9895 a_15227_44166# a_18315_45260# 0.272047f
C9896 a_3483_46348# a_5147_45002# 0.363215f
C9897 a_n755_45592# a_7499_43078# 0.157526f
C9898 a_6151_47436# a_12861_44030# 0.39397f
C9899 a_n2288_47178# a_n2312_39304# 0.01565f
C9900 a_8515_42308# a_8325_42308# 0.134955f
C9901 a_5934_30871# a_8685_42308# 0.186981f
C9902 a_5342_30871# VCM 0.325566f
C9903 a_n2017_45002# a_1067_42314# 0.01039f
C9904 a_10807_43548# a_10695_43548# 0.159782f
C9905 a_14840_46494# VDD 0.275785f
C9906 a_14401_32519# a_20974_43370# 0.118041f
C9907 a_10227_46804# a_10341_43396# 0.188948f
C9908 a_2324_44458# a_6109_44484# 0.101116f
C9909 a_8746_45002# a_8953_45002# 0.257529f
C9910 a_n1613_43370# a_6031_43396# 0.308901f
C9911 a_5937_45572# a_n2661_42834# 0.043505f
C9912 a_8199_44636# a_n2661_43922# 0.04879f
C9913 a_16327_47482# a_3090_45724# 1.00134f
C9914 a_15811_47375# a_15559_46634# 0.018669f
C9915 a_n743_46660# a_2107_46812# 0.72755f
C9916 a_n2438_43548# a_948_46660# 0.054839f
C9917 a_n133_46660# a_1123_46634# 0.043619f
C9918 a_10227_46804# a_12991_46634# 0.349162f
C9919 a_n881_46662# a_7411_46660# 0.025876f
C9920 a_33_46660# a_601_46902# 0.17072f
C9921 a_1273_38525# a_2684_37794# 0.224374f
C9922 a_5932_42308# C3_P_btm 0.121156f
C9923 a_n3420_39072# a_n4064_38528# 7.47287f
C9924 a_n2946_39072# a_n2946_38778# 0.050477f
C9925 a_1666_39043# a_2112_39137# 0.553829f
C9926 a_n4064_39072# a_n3420_38528# 0.048218f
C9927 a_16137_43396# a_15743_43084# 0.029757f
C9928 a_16977_43638# a_17324_43396# 0.051162f
C9929 a_20193_45348# a_17303_42282# 0.013391f
C9930 a_n2293_43922# a_n4318_37592# 0.019728f
C9931 a_16115_45572# VDD 0.194492f
C9932 a_n2956_37592# a_n2302_37690# 0.04217f
C9933 a_18184_42460# a_19647_42308# 0.034507f
C9934 a_18494_42460# a_19511_42282# 0.047119f
C9935 a_17339_46660# a_10341_43396# 0.023552f
C9936 a_n357_42282# a_3905_42865# 0.059842f
C9937 a_n2840_45002# a_n2840_44458# 0.025171f
C9938 a_13661_43548# a_10809_44734# 0.043589f
C9939 a_15559_46634# a_13059_46348# 0.167936f
C9940 a_11599_46634# a_19443_46116# 0.026712f
C9941 a_n443_46116# a_1848_45724# 0.041711f
C9942 a_22589_40599# VDD 0.821011f
C9943 CAL_N RST_Z 0.058301f
C9944 a_n4064_37440# VREF_GND 0.048151f
C9945 a_18194_34908# a_19998_34978# 0.04535f
C9946 EN_VIN_BSTR_P C8_P_btm 0.090252f
C9947 a_3422_30871# a_n3420_38528# 0.031237f
C9948 a_n2267_44484# VDD 0.289888f
C9949 a_n443_42852# a_14955_43396# 0.076467f
C9950 a_11691_44458# a_n2661_42834# 0.018854f
C9951 a_765_45546# a_13259_45724# 0.036082f
C9952 a_10903_43370# a_13351_46090# 0.181897f
C9953 a_12005_46116# a_12594_46348# 0.065075f
C9954 a_743_42282# a_4958_30871# 0.063224f
C9955 a_19339_43156# a_19164_43230# 0.233657f
C9956 a_19478_44306# VDD 0.127794f
C9957 a_n2312_39304# VDD 0.587668f
C9958 a_18114_32519# a_14401_32519# 0.087478f
C9959 a_n913_45002# a_4361_42308# 0.250497f
C9960 a_n1613_43370# a_n1809_44850# 0.012196f
C9961 a_3090_45724# a_14537_43396# 0.530123f
C9962 a_8953_45546# a_8696_44636# 0.022578f
C9963 a_20202_43084# a_2437_43646# 0.129143f
C9964 a_11415_45002# a_21513_45002# 0.050445f
C9965 a_5257_43370# a_n2661_43370# 0.027779f
C9966 a_n2472_45546# a_n2956_38216# 0.157892f
C9967 a_n2661_45546# a_n2293_45546# 0.077901f
C9968 a_n2497_47436# a_n1761_44111# 0.045728f
C9969 a_n815_47178# a_n971_45724# 0.013837f
C9970 a_n2109_47186# a_327_47204# 0.041762f
C9971 a_n2472_42826# VDD 0.229608f
C9972 a_22165_42308# a_21613_42308# 0.027246f
C9973 a_1184_42692# a_961_42354# 0.100246f
C9974 a_n1794_35082# a_1606_42308# 0.032246f
C9975 a_18579_44172# a_10341_43396# 0.023217f
C9976 a_15493_43396# a_19319_43548# 0.120111f
C9977 a_7499_43078# a_9885_42558# 0.020607f
C9978 a_n1613_43370# a_6671_43940# 0.03314f
C9979 a_3316_45546# a_2680_45002# 0.050127f
C9980 a_n443_46116# a_1512_43396# 0.010064f
C9981 a_17715_44484# a_11691_44458# 0.036149f
C9982 a_10227_46804# a_n97_42460# 0.18445f
C9983 a_2747_46873# a_n2661_46634# 0.019513f
C9984 a_n2312_39304# a_n2312_38680# 0.082563f
C9985 a_20974_43370# a_22223_43396# 0.04256f
C9986 a_14401_32519# a_13887_32519# 0.07508f
C9987 a_6511_45714# VDD 0.405279f
C9988 a_7276_45260# a_7229_43940# 0.322065f
C9989 a_5205_44484# a_6709_45028# 0.095031f
C9990 a_11823_42460# a_12883_44458# 0.026633f
C9991 a_18479_45785# a_16922_45042# 0.02321f
C9992 a_16147_45260# a_17613_45144# 0.028566f
C9993 a_n443_42852# a_n2661_42834# 0.076984f
C9994 a_3232_43370# a_8953_45002# 0.012103f
C9995 a_6171_45002# a_8191_45002# 0.024424f
C9996 a_6755_46942# a_11813_46116# 0.028837f
C9997 a_16327_47482# a_20075_46420# 0.270434f
C9998 a_1799_45572# a_765_45546# 0.225248f
C9999 a_22612_30879# a_20820_30879# 0.061094f
C10000 a_15507_47210# a_6945_45028# 0.04755f
C10001 a_4338_37500# a_6886_37412# 1.95816f
C10002 a_3726_37500# VDAC_N 0.06247f
C10003 a_n3420_38528# VDD 0.523642f
C10004 a_5088_37509# a_5700_37509# 1.48771f
C10005 a_n3420_39072# VREF_GND 0.066097f
C10006 a_375_42282# a_n2661_42834# 0.035547f
C10007 a_1823_45246# a_4520_42826# 0.053569f
C10008 a_14537_43396# a_14815_43914# 0.015948f
C10009 a_1307_43914# a_n2293_43922# 0.022859f
C10010 SMPL_ON_N a_n1794_35082# 0.150383f
C10011 w_10694_33990# a_4958_30871# 0.016533f
C10012 a_12549_44172# a_11962_45724# 0.034917f
C10013 a_17339_46660# a_17957_46116# 0.098952f
C10014 a_765_45546# a_18189_46348# 0.013467f
C10015 a_n2293_46098# a_4419_46090# 0.051687f
C10016 a_1208_46090# a_1138_42852# 0.043831f
C10017 a_2063_45854# a_2437_43646# 0.392331f
C10018 a_n971_45724# a_n2661_45010# 0.017233f
C10019 a_4361_42308# a_1755_42282# 0.015476f
C10020 a_12281_43396# a_12563_42308# 0.173003f
C10021 a_3422_30871# VIN_N 0.057975f
C10022 a_n4318_38680# a_n4318_38216# 0.055776f
C10023 a_n2065_43946# VDD 0.4213f
C10024 a_1307_43914# a_n97_42460# 0.23336f
C10025 a_4223_44672# a_n2661_42282# 0.064384f
C10026 a_3232_43370# a_3626_43646# 0.204337f
C10027 a_7499_43078# a_10083_42826# 0.375624f
C10028 a_n746_45260# DATA[0] 0.03466f
C10029 a_n971_45724# DATA[1] 0.050116f
C10030 a_20193_45348# a_20365_43914# 0.025746f
C10031 a_n356_44636# a_453_43940# 0.02089f
C10032 a_1209_47178# VDD 0.38145f
C10033 a_9313_44734# a_20512_43084# 0.028182f
C10034 a_16922_45042# a_14021_43940# 0.11663f
C10035 a_3483_46348# a_7499_43078# 0.207714f
C10036 a_5807_45002# a_n2661_43370# 0.018021f
C10037 a_5204_45822# a_4880_45572# 0.046074f
C10038 a_13667_43396# VDD 0.402378f
C10039 a_5342_30871# a_n4064_38528# 0.028644f
C10040 a_5891_43370# a_9803_43646# 0.011447f
C10041 a_14539_43914# a_16409_43396# 0.031761f
C10042 a_22485_44484# a_14401_32519# 0.01705f
C10043 a_20512_43084# a_20974_43370# 0.020132f
C10044 a_n755_45592# a_5932_42308# 0.040158f
C10045 a_10768_47026# VDD 0.132317f
C10046 a_n2956_38680# a_n4209_39590# 0.020934f
C10047 a_n2497_47436# a_n2267_43396# 0.222725f
C10048 a_18479_47436# a_20623_43914# 0.012705f
C10049 a_11525_45546# a_11962_45724# 0.095856f
C10050 a_11322_45546# a_12427_45724# 0.010517f
C10051 a_10490_45724# a_11823_42460# 0.022778f
C10052 a_2063_45854# a_n2661_46634# 1.75382f
C10053 a_4915_47217# a_5807_45002# 0.766023f
C10054 a_9313_45822# a_11309_47204# 0.027145f
C10055 a_n237_47217# a_n2438_43548# 0.02231f
C10056 a_n746_45260# a_n133_46660# 0.042075f
C10057 a_n4318_38216# a_n4209_38216# 0.135236f
C10058 a_14021_43940# a_15743_43084# 0.045789f
C10059 a_3080_42308# a_3539_42460# 0.037567f
C10060 a_n2661_45010# a_n2293_45010# 0.400159f
C10061 a_4955_46873# a_5072_46660# 0.17431f
C10062 a_5385_46902# a_5732_46660# 0.051162f
C10063 a_2747_46873# a_765_45546# 0.040029f
C10064 a_n1151_42308# a_6165_46155# 0.055317f
C10065 a_2063_45854# a_8199_44636# 0.037924f
C10066 a_10227_46804# a_11415_45002# 0.139042f
C10067 a_11453_44696# a_20841_46902# 0.0185f
C10068 a_4958_30871# C9_N_btm 0.209166f
C10069 a_12281_43396# a_12089_42308# 0.210903f
C10070 a_22223_43396# a_13887_32519# 0.154411f
C10071 a_13678_32519# a_14209_32519# 0.048492f
C10072 a_n2810_45028# VDD 0.526631f
C10073 a_19963_31679# VIN_N 0.02847f
C10074 a_19479_31679# VCM 0.03628f
C10075 a_1307_43914# a_742_44458# 0.355379f
C10076 a_10775_45002# a_10057_43914# 0.010331f
C10077 a_2711_45572# a_15682_43940# 0.038198f
C10078 a_n913_45002# a_5891_43370# 0.255618f
C10079 a_2437_43646# a_n2661_42834# 0.033942f
C10080 a_526_44458# a_3080_42308# 0.041925f
C10081 a_9290_44172# a_9803_43646# 0.010228f
C10082 a_15227_44166# a_3483_46348# 0.595533f
C10083 a_17339_46660# a_11415_45002# 0.025523f
C10084 a_6755_46942# a_15682_46116# 0.116442f
C10085 a_4646_46812# a_526_44458# 0.020719f
C10086 a_3877_44458# a_n1925_42282# 0.034241f
C10087 VDD VIN_N 1.51335f
C10088 C10_N_btm VREF_GND 10.3207f
C10089 C9_N_btm VCM 6.06251f
C10090 a_3422_30871# CAL_N 0.236929f
C10091 a_3626_43646# a_6123_31319# 0.109715f
C10092 a_2982_43646# a_5934_30871# 0.178f
C10093 a_9482_43914# a_11173_44260# 0.043729f
C10094 a_n2293_42834# a_n2661_42282# 0.026231f
C10095 a_13259_45724# a_13460_43230# 0.015281f
C10096 a_n2312_39304# a_n2946_39072# 0.020842f
C10097 a_n2497_47436# a_n2267_44484# 0.025633f
C10098 a_15682_46116# a_8049_45260# 0.015666f
C10099 a_1138_42852# a_n2661_45546# 0.023338f
C10100 a_21588_30879# a_413_45260# 0.041669f
C10101 a_n1853_46287# a_n755_45592# 0.021472f
C10102 a_n2438_43548# a_n2017_45002# 0.29197f
C10103 a_n2312_38680# a_n2810_45028# 0.044149f
C10104 a_n2129_43609# VDD 0.400674f
C10105 a_19279_43940# a_15493_43940# 0.019758f
C10106 a_9313_44734# a_21381_43940# 0.028978f
C10107 a_288_46660# VDD 0.079457f
C10108 en_comp a_5342_30871# 0.032532f
C10109 a_n1059_45260# a_17701_42308# 0.073596f
C10110 a_n2017_45002# a_18083_42858# 0.03192f
C10111 a_4185_45028# a_3537_45260# 1.06643f
C10112 a_19692_46634# a_16922_45042# 0.055961f
C10113 a_5257_43370# a_5883_43914# 0.019234f
C10114 a_2324_44458# a_3357_43084# 0.216574f
C10115 a_9290_44172# a_n913_45002# 0.632534f
C10116 a_3483_46348# a_4558_45348# 0.068916f
C10117 a_n357_42282# a_7499_43078# 0.259858f
C10118 a_15227_44166# a_17719_45144# 0.187414f
C10119 a_6151_47436# a_13717_47436# 0.17202f
C10120 a_n2288_47178# a_n2312_40392# 0.153632f
C10121 a_n2497_47436# a_n2312_39304# 0.061823f
C10122 a_n971_45724# a_4883_46098# 0.031452f
C10123 a_5934_30871# a_8325_42308# 0.173576f
C10124 a_5342_30871# VREF_GND 0.055227f
C10125 a_17730_32519# a_13678_32519# 0.054146f
C10126 a_21381_43940# a_20974_43370# 0.02221f
C10127 a_n2017_45002# a_n1794_35082# 0.111641f
C10128 a_9290_44172# CLK 0.151406f
C10129 a_15015_46420# VDD 0.337162f
C10130 a_n967_45348# a_n961_42308# 0.174237f
C10131 a_n1059_45260# a_564_42282# 0.043244f
C10132 a_n755_45592# a_n2661_43370# 0.036276f
C10133 a_10903_43370# a_9313_44734# 0.030402f
C10134 a_11823_42460# a_6171_45002# 0.123118f
C10135 a_10180_45724# a_10775_45002# 0.073185f
C10136 a_8199_44636# a_n2661_42834# 0.032396f
C10137 a_n743_46660# a_948_46660# 0.038448f
C10138 a_n2438_43548# a_1123_46634# 0.075317f
C10139 a_n133_46660# a_383_46660# 0.105995f
C10140 a_2063_45854# a_765_45546# 1.71006f
C10141 a_10227_46804# a_12251_46660# 0.188053f
C10142 a_15507_47210# a_15559_46634# 0.011624f
C10143 a_n881_46662# a_5257_43370# 0.447042f
C10144 a_2351_42308# VDD 0.188239f
C10145 a_1273_38525# a_1107_38525# 0.236832f
C10146 a_5932_42308# C4_P_btm 0.032349f
C10147 a_n4064_39616# a_n3420_37984# 0.050009f
C10148 a_n3420_39616# a_n4064_37984# 0.046151f
C10149 a_4958_30871# a_n3420_37440# 0.033151f
C10150 a_16409_43396# a_17324_43396# 0.118759f
C10151 a_16333_45814# VDD 0.201203f
C10152 a_n2956_37592# a_n4064_37440# 0.070596f
C10153 a_18184_42460# a_19511_42282# 0.058931f
C10154 a_n2810_45028# a_n2302_37690# 0.162246f
C10155 a_n2810_45572# a_n3674_39768# 0.023119f
C10156 a_n881_46662# a_1337_46116# 0.043447f
C10157 a_2107_46812# a_9290_44172# 0.091636f
C10158 a_5807_45002# a_10809_44734# 0.065594f
C10159 a_13747_46662# a_6945_45028# 0.035381f
C10160 a_n2293_46634# a_2324_44458# 0.021161f
C10161 a_15368_46634# a_13059_46348# 0.101997f
C10162 a_n443_46116# a_997_45618# 0.080297f
C10163 a_10227_46804# a_13259_45724# 0.335001f
C10164 a_584_46384# a_n443_42852# 1.36389f
C10165 a_n743_46660# a_13925_46122# 0.041274f
C10166 CAL_N VDD 26.0839f
C10167 a_11206_38545# RST_Z 0.382319f
C10168 a_n3420_37440# VCM 0.033198f
C10169 EN_VIN_BSTR_N a_19998_34978# 0.573018f
C10170 a_18194_34908# a_19250_34978# 0.559484f
C10171 EN_VIN_BSTR_P C9_P_btm 0.226529f
C10172 a_n2129_44697# VDD 1.4165f
C10173 a_n4318_39304# a_n3674_37592# 0.024848f
C10174 a_n913_45002# a_10807_43548# 0.023237f
C10175 a_7229_43940# a_7542_44172# 0.086946f
C10176 a_2382_45260# a_3499_42826# 0.040227f
C10177 a_n2661_44458# a_5891_43370# 0.013115f
C10178 a_526_44458# a_2075_43172# 0.227071f
C10179 a_10193_42453# a_3626_43646# 0.13905f
C10180 a_584_46384# a_375_42282# 0.480677f
C10181 a_n743_46660# a_15599_45572# 0.022482f
C10182 a_17339_46660# a_13259_45724# 0.038367f
C10183 a_10903_43370# a_12594_46348# 0.169312f
C10184 a_15227_44166# a_n357_42282# 0.023198f
C10185 a_4190_30871# a_17303_42282# 0.279034f
C10186 a_15493_43396# VDD 2.34659f
C10187 a_20447_31679# a_17364_32525# 0.054026f
C10188 a_n2312_40392# VDD 0.947797f
C10189 a_n913_45002# a_13467_32519# 0.024166f
C10190 a_n1059_45260# a_4361_42308# 0.033614f
C10191 a_5937_45572# a_8696_44636# 0.041815f
C10192 a_20202_43084# a_21513_45002# 0.13666f
C10193 a_4883_46098# a_9313_44734# 0.015767f
C10194 a_10227_46804# a_n2661_43922# 0.041913f
C10195 a_768_44030# a_13720_44458# 0.178939f
C10196 a_n2661_45546# a_n2956_38216# 0.15505f
C10197 a_n2497_47436# a_n2065_43946# 0.036632f
C10198 a_n815_47178# a_n452_47436# 0.107449f
C10199 a_n1741_47186# a_n237_47217# 0.083957f
C10200 a_n2109_47186# a_n785_47204# 0.43597f
C10201 a_n2840_42826# VDD 0.302305f
C10202 a_22165_42308# a_21887_42336# 0.110763f
C10203 a_9313_44734# a_5649_42852# 0.028023f
C10204 a_18451_43940# a_18533_43940# 0.171361f
C10205 a_19328_44172# a_19319_43548# 0.033025f
C10206 a_n2810_45572# a_n4315_30879# 0.024132f
C10207 a_13259_45724# a_1307_43914# 0.023098f
C10208 a_3316_45546# a_2382_45260# 0.052075f
C10209 a_n971_45724# a_8685_43396# 0.079658f
C10210 a_9290_44172# a_n2661_44458# 0.027487f
C10211 a_3483_46348# a_9838_44484# 0.014242f
C10212 a_12549_44172# a_768_44030# 0.490163f
C10213 a_n881_46662# a_5807_45002# 0.243322f
C10214 a_n2312_40392# a_n2312_38680# 0.052461f
C10215 a_n2312_39304# a_n2104_46634# 0.018871f
C10216 COMP_P a_22527_39145# 0.033008f
C10217 a_20974_43370# a_5649_42852# 0.186094f
C10218 a_6472_45840# VDD 0.257073f
C10219 a_17538_32519# a_13678_32519# 0.051187f
C10220 a_11823_42460# a_12607_44458# 0.01822f
C10221 a_n2293_46098# a_5829_43940# 0.05512f
C10222 a_8696_44636# a_11691_44458# 0.141053f
C10223 a_16147_45260# a_17023_45118# 0.040001f
C10224 a_3232_43370# a_8191_45002# 0.045343f
C10225 a_6431_45366# a_6709_45028# 0.112564f
C10226 a_6755_46942# a_11735_46660# 0.61229f
C10227 a_n881_46662# a_3699_46348# 0.203393f
C10228 a_n1741_47186# a_12638_46436# 0.016323f
C10229 a_16327_47482# a_19335_46494# 0.155998f
C10230 a_20916_46384# a_12741_44636# 0.023496f
C10231 a_21588_30879# a_20820_30879# 0.084472f
C10232 a_4883_46098# a_12594_46348# 0.022174f
C10233 a_11599_46634# a_6945_45028# 0.04727f
C10234 a_11453_44696# a_9290_44172# 0.064153f
C10235 a_3726_37500# a_6886_37412# 0.702909f
C10236 a_n3690_38528# VDD 0.363159f
C10237 a_4338_37500# a_5700_37509# 2.69237f
C10238 a_n3565_39304# VCM 0.035438f
C10239 a_n4064_39072# VIN_P 0.038211f
C10240 a_n2661_42282# a_5379_42460# 0.121051f
C10241 a_20447_31679# a_19237_31679# 0.051563f
C10242 a_1307_43914# a_n2661_43922# 0.023892f
C10243 a_17339_46660# a_18189_46348# 0.170772f
C10244 a_765_45546# a_17715_44484# 0.117636f
C10245 a_n2293_46098# a_4185_45028# 0.06423f
C10246 a_1208_46090# a_1176_45822# 0.141891f
C10247 a_n881_46662# a_15143_45578# 0.069805f
C10248 a_584_46384# a_2437_43646# 0.302508f
C10249 a_3422_30871# VIN_P 0.057975f
C10250 a_n3674_39304# a_n4318_38216# 0.043431f
C10251 a_12895_43230# a_12991_43230# 0.013793f
C10252 a_n2472_43914# VDD 0.236691f
C10253 a_7499_43078# a_8952_43230# 0.054554f
C10254 a_n356_44636# a_1414_42308# 0.179164f
C10255 a_11827_44484# a_11341_43940# 0.231114f
C10256 a_n971_45724# DATA[0] 0.213213f
C10257 a_n1741_47186# DATA[5] 0.069294f
C10258 a_327_47204# VDD 0.367528f
C10259 a_5937_45572# a_7227_45028# 0.064518f
C10260 a_n1151_42308# a_n23_44458# 0.101137f
C10261 a_10903_43370# a_2711_45572# 0.213719f
C10262 a_3483_46348# a_8568_45546# 0.137016f
C10263 a_10695_43548# VDD 0.201247f
C10264 a_19721_31679# a_13678_32519# 0.051384f
C10265 a_5891_43370# a_9145_43396# 0.049186f
C10266 a_9313_44734# a_8685_43396# 0.124273f
C10267 a_14539_43914# a_16547_43609# 0.01221f
C10268 a_n2956_39304# a_n4209_39590# 0.022939f
C10269 a_10490_45724# a_12427_45724# 0.108721f
C10270 a_n2497_47436# a_n2129_43609# 0.216536f
C10271 a_18597_46090# a_19862_44208# 0.536021f
C10272 a_11415_45002# a_22223_45036# 0.011148f
C10273 a_11322_45546# a_11962_45724# 0.270736f
C10274 a_11525_45546# a_11652_45724# 0.138143f
C10275 a_3483_46348# a_n2661_43370# 0.953959f
C10276 a_584_46384# a_n2661_46634# 0.034039f
C10277 a_11031_47542# a_11309_47204# 0.110775f
C10278 a_n746_45260# a_n2438_43548# 0.031949f
C10279 a_n237_47217# a_n743_46660# 0.192378f
C10280 a_n971_45724# a_n133_46660# 0.011188f
C10281 a_4883_46098# a_12465_44636# 0.024607f
C10282 a_n2109_47186# a_2107_46812# 0.032545f
C10283 a_14311_47204# a_n881_46662# 0.037789f
C10284 a_14113_42308# a_4958_30871# 0.058048f
C10285 a_4699_43561# a_3539_42460# 0.109444f
C10286 a_3080_42308# a_3626_43646# 0.092602f
C10287 a_n2661_45010# a_n2472_45002# 0.065751f
C10288 a_n2293_46634# a_14579_43548# 0.035629f
C10289 a_15861_45028# a_16751_45260# 0.044248f
C10290 a_4791_45118# a_4185_45028# 0.064362f
C10291 a_4651_46660# a_5072_46660# 0.083408f
C10292 a_4817_46660# a_5732_46660# 0.118759f
C10293 a_n2661_46634# a_11901_46660# 0.030789f
C10294 a_n743_46660# a_8270_45546# 0.274248f
C10295 a_10227_46804# a_20202_43084# 0.022898f
C10296 a_11453_44696# a_20273_46660# 0.545219f
C10297 a_n1151_42308# a_5497_46414# 0.089064f
C10298 a_n4064_40160# EN_VIN_BSTR_P 0.149623f
C10299 a_n4064_38528# a_n3420_37440# 0.050813f
C10300 a_n3420_38528# a_n4064_37440# 0.045626f
C10301 a_14579_43548# a_5342_30871# 0.041574f
C10302 a_12281_43396# a_12379_42858# 0.036584f
C10303 a_13467_32519# a_17364_32525# 0.050014f
C10304 a_n745_45366# VDD 0.20887f
C10305 a_n1761_44111# a_n473_42460# 0.110251f
C10306 a_327_44734# a_n23_44458# 0.141544f
C10307 a_n1925_42282# a_4235_43370# 0.199349f
C10308 a_n1059_45260# a_5891_43370# 0.186322f
C10309 a_9290_44172# a_9145_43396# 0.103991f
C10310 a_4883_46098# a_2711_45572# 0.041245f
C10311 a_768_44030# a_n2661_45546# 0.07332f
C10312 a_n881_46662# a_n755_45592# 0.077214f
C10313 a_6755_46942# a_2324_44458# 0.155169f
C10314 a_3877_44458# a_526_44458# 0.017621f
C10315 RST_Z CLK 0.064624f
C10316 C10_N_btm VREF 14.773f
C10317 C9_N_btm VREF_GND 5.18245f
C10318 C8_N_btm VCM 2.61094f
C10319 VDD VIN_P 1.52779f
C10320 a_n97_42460# a_14456_42282# 0.067807f
C10321 a_9482_43914# a_10555_44260# 0.088693f
C10322 a_n863_45724# a_2905_42968# 0.269475f
C10323 a_14539_43914# a_14673_44172# 0.205935f
C10324 a_16112_44458# a_16241_44734# 0.062574f
C10325 a_13259_45724# a_13635_43156# 0.017822f
C10326 a_n2497_47436# a_n2129_44697# 0.019202f
C10327 a_2324_44458# a_8049_45260# 0.054166f
C10328 a_768_44030# a_5205_44484# 0.033081f
C10329 a_n2442_46660# en_comp 0.02478f
C10330 a_5534_30871# a_4958_30871# 0.024536f
C10331 a_n2433_43396# VDD 0.416276f
C10332 a_1983_46706# VDD 0.119964f
C10333 a_4185_45028# a_13258_32519# 0.068774f
C10334 a_n1059_45260# a_17595_43084# 0.049f
C10335 a_n2017_45002# a_17701_42308# 0.132871f
C10336 a_7542_44172# a_7845_44172# 0.137004f
C10337 a_12549_44172# a_17517_44484# 0.019389f
C10338 a_3483_46348# a_4574_45260# 0.022358f
C10339 a_19466_46812# a_16922_45042# 0.030378f
C10340 a_9290_44172# a_n1059_45260# 0.092471f
C10341 a_15227_44166# a_17613_45144# 0.048772f
C10342 a_6151_47436# a_n1435_47204# 0.061966f
C10343 a_6575_47204# a_9067_47204# 0.210614f
C10344 a_4915_47217# a_13487_47204# 0.013601f
C10345 a_2063_45854# a_10227_46804# 0.186188f
C10346 a_n2497_47436# a_n2312_40392# 0.194574f
C10347 a_5534_30871# VCM 0.095752f
C10348 a_10807_43548# a_9145_43396# 0.290878f
C10349 a_9313_44734# a_17333_42852# 0.010555f
C10350 a_19237_31679# a_13467_32519# 0.052472f
C10351 a_n967_45348# a_n1329_42308# 0.033651f
C10352 a_14275_46494# VDD 0.196859f
C10353 a_n2017_45002# a_564_42282# 0.013024f
C10354 a_n357_42282# a_n2661_43370# 0.034578f
C10355 a_10227_46804# a_14955_43396# 0.035123f
C10356 a_10180_45724# a_8953_45002# 0.107499f
C10357 a_12861_44030# a_15781_43660# 0.025765f
C10358 a_18691_45572# a_18799_45938# 0.057222f
C10359 a_5937_45572# a_9159_44484# 0.040512f
C10360 a_8016_46348# a_n2661_43922# 0.02895f
C10361 a_12861_44030# a_15227_44166# 0.810382f
C10362 a_n743_46660# a_1123_46634# 0.054493f
C10363 a_n2438_43548# a_383_46660# 0.0336f
C10364 a_n133_46660# a_601_46902# 0.053479f
C10365 a_584_46384# a_765_45546# 0.086068f
C10366 a_n1613_43370# a_5257_43370# 0.025984f
C10367 a_n1925_46634# a_2107_46812# 1.12874f
C10368 a_171_46873# a_33_46660# 0.207108f
C10369 a_11599_46634# a_15559_46634# 0.028826f
C10370 a_10227_46804# a_12469_46902# 0.181535f
C10371 a_n3565_39304# a_n4064_38528# 0.029566f
C10372 a_n3420_39072# a_n3420_38528# 0.127439f
C10373 a_n4064_39072# a_n3565_38502# 0.030685f
C10374 a_2123_42473# VDD 0.1936f
C10375 a_16409_43396# a_17499_43370# 0.042737f
C10376 a_16977_43638# a_16759_43396# 0.209641f
C10377 a_n2956_37592# a_n2946_37690# 0.148852f
C10378 a_n2293_43922# a_n3674_38216# 0.032717f
C10379 a_15765_45572# VDD 0.249471f
C10380 a_n2810_45028# a_n4064_37440# 0.22413f
C10381 a_n2810_45572# a_n4318_39768# 0.023737f
C10382 a_5257_43370# a_n2293_46098# 0.049293f
C10383 a_13661_43548# a_6945_45028# 0.015293f
C10384 a_15368_46634# a_15227_46910# 0.050747f
C10385 a_n443_46116# a_n755_45592# 0.651643f
C10386 a_10227_46804# a_14383_46116# 0.01306f
C10387 a_14976_45028# a_13059_46348# 0.209989f
C10388 a_n743_46660# a_13759_46122# 0.01783f
C10389 a_n3420_37440# VREF_GND 0.033872f
C10390 a_11206_38545# VDD 8.87267f
C10391 a_10890_34112# a_19998_34978# 0.201872f
C10392 EN_VIN_BSTR_N a_19250_34978# 0.651142f
C10393 VDAC_P RST_Z 0.158793f
C10394 EN_VIN_BSTR_P C10_P_btm 0.320569f
C10395 a_18249_42858# a_18817_42826# 0.16939f
C10396 a_n2433_44484# VDD 0.40658f
C10397 a_n699_43396# a_n356_44636# 0.044884f
C10398 a_n1059_45260# a_10807_43548# 0.031771f
C10399 a_n443_42852# a_14205_43396# 0.118229f
C10400 a_7229_43940# a_7281_43914# 0.164835f
C10401 a_11827_44484# a_n2293_43922# 0.028646f
C10402 a_526_44458# a_1847_42826# 0.154735f
C10403 a_8953_45546# a_2324_44458# 0.047906f
C10404 a_3483_46348# a_10809_44734# 0.02965f
C10405 a_3090_45724# a_3316_45546# 0.04556f
C10406 SMPL_ON_N a_20447_31679# 0.029368f
C10407 a_10903_43370# a_12005_46116# 0.277468f
C10408 a_4190_30871# a_4958_30871# 11.510201f
C10409 a_19328_44172# VDD 0.263964f
C10410 a_22959_47212# VDD 0.245964f
C10411 a_n2661_45546# a_n2472_45546# 0.040937f
C10412 a_8199_44636# a_8696_44636# 0.265919f
C10413 a_10227_46804# a_n2661_42834# 0.024624f
C10414 a_768_44030# a_13076_44458# 0.132449f
C10415 a_5066_45546# a_4880_45572# 0.04794f
C10416 a_10903_43370# a_14033_45822# 0.040019f
C10417 a_n2810_45572# a_n2956_38216# 6.20057f
C10418 a_17364_32525# RST_Z 0.050609f
C10419 a_n1741_47186# a_n746_45260# 0.032595f
C10420 a_n2109_47186# a_n23_47502# 0.043455f
C10421 a_4190_30871# VCM 1.23535f
C10422 a_1576_42282# a_1184_42692# 0.033078f
C10423 a_n784_42308# a_2123_42473# 0.216332f
C10424 a_1067_42314# a_961_42354# 0.13675f
C10425 a_n473_42460# a_n327_42308# 0.013377f
C10426 a_9313_44734# a_13678_32519# 0.097255f
C10427 a_n357_42282# a_20712_42282# 0.173926f
C10428 a_n755_45592# a_3537_45260# 0.025346f
C10429 a_12891_46348# a_768_44030# 0.193145f
C10430 a_n1613_43370# a_5807_45002# 0.086053f
C10431 a_2063_45854# a_10467_46802# 0.036614f
C10432 a_4791_45118# a_5257_43370# 0.36404f
C10433 a_n2312_39304# a_n2293_46634# 0.021162f
C10434 a_8495_42852# VDD 0.132018f
C10435 a_20974_43370# a_13678_32519# 0.020999f
C10436 a_6194_45824# VDD 0.274689f
C10437 a_n4318_40392# a_n3674_37592# 0.032206f
C10438 a_3090_45724# a_6197_43396# 0.010809f
C10439 a_10193_42453# a_16979_44734# 0.016398f
C10440 a_n2293_46098# a_5745_43940# 0.019006f
C10441 a_n1925_42282# a_3905_42865# 0.023709f
C10442 a_16147_45260# a_16922_45042# 0.016249f
C10443 a_3232_43370# a_7705_45326# 0.02181f
C10444 a_6171_45002# a_6709_45028# 0.021915f
C10445 a_6755_46942# a_11186_47026# 0.014167f
C10446 a_n881_46662# a_3483_46348# 0.5947f
C10447 a_n1741_47186# a_12379_46436# 0.067348f
C10448 a_16327_47482# a_19553_46090# 0.172776f
C10449 a_14955_47212# a_6945_45028# 0.013254f
C10450 a_13507_46334# a_13351_46090# 0.214666f
C10451 a_4883_46098# a_12005_46116# 0.012933f
C10452 a_2063_45854# a_8034_45724# 0.034258f
C10453 a_n3565_38502# VDD 0.774466f
C10454 a_4338_37500# a_5088_37509# 0.896828f
C10455 a_3726_37500# a_5700_37509# 0.574743f
C10456 a_n3565_39304# VREF_GND 0.010456f
C10457 a_n4064_37984# C3_P_btm 0.030933f
C10458 a_13556_45296# a_15433_44458# 0.1084f
C10459 a_n913_45002# a_3422_30871# 0.145467f
C10460 a_n357_42282# a_1568_43370# 0.036942f
C10461 a_1307_43914# a_n2661_42834# 3.43601f
C10462 a_17339_46660# a_17715_44484# 0.018672f
C10463 a_765_45546# a_17583_46090# 0.067337f
C10464 a_472_46348# a_1138_42852# 0.028956f
C10465 a_805_46414# a_1176_45822# 0.024739f
C10466 a_2124_47436# a_2437_43646# 0.025048f
C10467 a_n881_46662# a_14495_45572# 0.170589f
C10468 a_n2840_43914# VDD 0.304745f
C10469 a_n4318_38680# a_n3674_38680# 3.04229f
C10470 a_19237_31679# RST_Z 0.050685f
C10471 a_12895_43230# a_12800_43218# 0.049827f
C10472 a_n4318_39304# a_n4064_39072# 0.017224f
C10473 a_3232_43370# a_2982_43646# 0.416054f
C10474 a_7499_43078# a_9127_43156# 0.08498f
C10475 a_n356_44636# a_1467_44172# 0.061333f
C10476 a_20193_45348# a_19862_44208# 0.041264f
C10477 a_n1741_47186# DATA[4] 0.020035f
C10478 a_n2312_38680# a_n3565_38502# 0.134976f
C10479 a_n452_47436# DATA[0] 0.039965f
C10480 a_n785_47204# VDD 0.452945f
C10481 a_n1151_42308# a_n356_44636# 0.093166f
C10482 a_5342_30871# a_n3420_38528# 0.028503f
C10483 a_9803_43646# VDD 0.261557f
C10484 a_5534_30871# a_n4064_38528# 0.057361f
C10485 a_14539_43914# a_16243_43396# 0.029808f
C10486 a_20512_43084# a_21381_43940# 0.019564f
C10487 a_n357_42282# a_6171_42473# 0.010166f
C10488 a_18114_32519# a_13678_32519# 0.055126f
C10489 a_3600_43914# a_3992_43940# 0.016359f
C10490 a_10490_45724# a_11962_45724# 0.114064f
C10491 a_10193_42453# a_11823_42460# 0.235429f
C10492 a_16327_47482# a_15493_43940# 0.04211f
C10493 a_11415_45002# a_11827_44484# 0.169126f
C10494 a_11322_45546# a_11652_45724# 0.26844f
C10495 a_526_44458# a_5111_44636# 0.338508f
C10496 a_n2497_47436# a_n2433_43396# 0.173242f
C10497 a_8270_45546# a_5891_43370# 0.052984f
C10498 a_4883_46098# a_21811_47423# 0.054014f
C10499 a_4791_45118# a_5807_45002# 0.129041f
C10500 a_13487_47204# a_n881_46662# 0.108977f
C10501 a_n746_45260# a_n743_46660# 0.068305f
C10502 a_n971_45724# a_n2438_43548# 0.038673f
C10503 a_15890_42674# a_16104_42674# 0.097745f
C10504 a_15959_42545# a_16522_42674# 0.049827f
C10505 a_15861_45028# a_1307_43914# 0.067929f
C10506 SMPL_ON_N a_13467_32519# 0.029246f
C10507 a_13507_46334# a_22591_43396# 0.011335f
C10508 a_n2293_46634# a_13667_43396# 0.011502f
C10509 a_8696_44636# a_16751_45260# 0.265287f
C10510 a_16327_47482# a_12741_44636# 0.074082f
C10511 a_4646_46812# a_5072_46660# 0.013764f
C10512 a_13747_46662# a_15368_46634# 0.110984f
C10513 a_5807_45002# a_16292_46812# 0.202526f
C10514 a_n881_46662# a_14513_46634# 0.017832f
C10515 a_5385_46902# a_5167_46660# 0.209641f
C10516 a_4817_46660# a_5907_46634# 0.042415f
C10517 a_n2661_46634# a_11813_46116# 0.162517f
C10518 a_19321_45002# a_3090_45724# 0.163821f
C10519 a_11453_44696# a_20411_46873# 0.020751f
C10520 a_n1151_42308# a_5204_45822# 0.487224f
C10521 a_17124_42282# VDD 0.28176f
C10522 a_n913_45002# VDD 9.190901f
C10523 a_14579_43548# a_15279_43071# 0.108607f
C10524 a_5649_42852# a_22223_43396# 0.165664f
C10525 a_13678_32519# a_13887_32519# 10.751599f
C10526 a_19479_31679# VREF 0.056254f
C10527 a_327_44734# a_n356_44636# 0.085841f
C10528 a_526_44458# a_4235_43370# 0.032501f
C10529 a_n1925_42282# a_4093_43548# 0.018682f
C10530 a_n2017_45002# a_5891_43370# 0.065487f
C10531 a_n971_45724# a_n1794_35082# 0.028303f
C10532 a_20623_46660# a_20731_47026# 0.057222f
C10533 a_n1613_43370# a_n755_45592# 0.052236f
C10534 a_6755_46942# a_14840_46494# 0.021842f
C10535 a_8270_45546# a_9290_44172# 0.433963f
C10536 a_4915_47217# a_13249_42308# 0.161597f
C10537 C9_N_btm VREF 7.369471f
C10538 C10_N_btm VIN_N 3.66034f
C10539 VDD CLK 0.49309f
C10540 C8_N_btm VREF_GND 2.58605f
C10541 C7_N_btm VCM 1.58335f
C10542 RST_Z EN_OFFSET_CAL 0.044122f
C10543 a_n97_42460# a_13575_42558# 0.179828f
C10544 a_3422_30871# VDAC_P 0.476125f
C10545 a_2982_43646# a_6123_31319# 0.163265f
C10546 a_n443_42852# a_n1853_43023# 0.141267f
C10547 a_16112_44458# a_14673_44172# 0.077293f
C10548 a_n2438_43548# a_n2293_45010# 0.033143f
C10549 a_n2293_46098# a_n755_45592# 0.086057f
C10550 a_n2442_46660# a_n2956_37592# 0.049818f
C10551 a_n2497_47436# a_n2433_44484# 0.027254f
C10552 a_4190_30871# a_n4064_38528# 0.031783f
C10553 a_n4318_39304# VDD 0.643395f
C10554 en_comp a_5534_30871# 0.021896f
C10555 a_2127_44172# a_2253_44260# 0.013015f
C10556 a_1414_42308# a_3499_42826# 0.023314f
C10557 a_n2017_45002# a_17595_43084# 0.016123f
C10558 a_n1059_45260# a_16795_42852# 0.182174f
C10559 a_2107_46812# VDD 0.350275f
C10560 a_10193_42453# a_20922_43172# 0.059157f
C10561 a_3483_46348# a_3537_45260# 0.605469f
C10562 a_1823_45246# a_3232_43370# 0.344002f
C10563 a_4185_45028# a_3065_45002# 0.060303f
C10564 a_9290_44172# a_n2017_45002# 0.089856f
C10565 a_12741_44636# a_14537_43396# 0.094691f
C10566 a_4915_47217# a_12861_44030# 0.025257f
C10567 a_6151_47436# a_13381_47204# 0.014822f
C10568 a_n2833_47464# a_n2312_40392# 0.064992f
C10569 a_5534_30871# VREF_GND 0.060532f
C10570 COMP_P a_4958_30871# 0.02709f
C10571 a_20512_43084# a_5649_42852# 0.141324f
C10572 a_9313_44734# a_18083_42858# 0.05022f
C10573 a_14493_46090# VDD 0.203567f
C10574 a_n2017_45002# a_n3674_37592# 0.241068f
C10575 a_13259_45724# a_11827_44484# 0.062801f
C10576 a_310_45028# a_n2661_43370# 0.027265f
C10577 a_10227_46804# a_15095_43370# 0.264777f
C10578 a_n2312_38680# a_n4318_39304# 0.023234f
C10579 a_19431_45546# a_19256_45572# 0.233657f
C10580 a_18909_45814# a_18799_45938# 0.097745f
C10581 a_18691_45572# a_18596_45572# 0.049827f
C10582 a_8016_46348# a_n2661_42834# 0.041785f
C10583 a_12861_44030# a_15681_43442# 0.137136f
C10584 a_4915_47217# a_14180_46812# 0.017902f
C10585 a_n743_46660# a_383_46660# 0.035839f
C10586 a_n2438_43548# a_601_46902# 0.043115f
C10587 a_n133_46660# a_33_46660# 0.580914f
C10588 a_11599_46634# a_15368_46634# 0.320705f
C10589 a_10227_46804# a_11901_46660# 0.055248f
C10590 a_1606_42308# RST_Z 1.44945f
C10591 a_1666_39587# a_2684_37794# 0.565516f
C10592 a_n3420_39072# a_n3690_38528# 0.017537f
C10593 a_n4064_39616# a_n3565_38216# 0.028071f
C10594 a_n3420_39616# a_n3420_37984# 0.047086f
C10595 a_n3565_39590# a_n4064_37984# 0.031327f
C10596 a_1755_42282# VDD 0.215277f
C10597 a_16243_43396# a_17324_43396# 0.102355f
C10598 a_16409_43396# a_16759_43396# 0.20669f
C10599 a_10341_43396# a_16823_43084# 0.044262f
C10600 a_n2956_37592# a_n3420_37440# 0.233174f
C10601 a_15903_45785# VDD 0.291109f
C10602 a_n2810_45028# a_n2946_37690# 0.024678f
C10603 a_4646_46812# a_7765_42852# 0.122773f
C10604 a_1823_45246# a_4905_42826# 0.110836f
C10605 a_16327_47482# a_16375_45002# 0.032962f
C10606 a_5807_45002# a_6945_45028# 0.057813f
C10607 a_n443_46116# a_n357_42282# 0.153614f
C10608 a_3090_45724# a_13059_46348# 0.167043f
C10609 a_14976_45028# a_15227_46910# 0.060892f
C10610 a_n3565_37414# VCM 0.03748f
C10611 a_n4064_37440# VIN_P 0.075801f
C10612 VDAC_P VDD 5.18919f
C10613 a_10890_34112# a_19250_34978# 0.481434f
C10614 EN_VIN_BSTR_N a_18194_34908# 0.335951f
C10615 a_8912_37509# RST_Z 0.082942f
C10616 a_n2661_44458# VDD 1.06317f
C10617 a_n2017_45002# a_10807_43548# 0.0319f
C10618 a_n443_42852# a_14358_43442# 0.037176f
C10619 a_10193_42453# a_2982_43646# 0.231527f
C10620 a_11827_44484# a_n2661_43922# 0.32722f
C10621 a_5937_45572# a_2324_44458# 0.407894f
C10622 a_3090_45724# a_3218_45724# 0.100752f
C10623 a_584_46384# a_1307_43914# 0.314947f
C10624 a_18451_43940# VDD 0.172318f
C10625 a_7871_42858# a_6123_31319# 0.010286f
C10626 a_n2293_43922# a_n2661_42282# 0.133253f
C10627 a_20447_31679# a_14209_32519# 0.051502f
C10628 en_comp a_4190_30871# 0.086973f
C10629 a_19963_31679# a_17364_32525# 0.053794f
C10630 a_11453_44696# VDD 3.75355f
C10631 SMPL_ON_N RST_Z 2.43362f
C10632 a_n2840_45546# a_n2956_38216# 0.019918f
C10633 a_3090_45724# a_13556_45296# 0.032207f
C10634 a_13507_46334# a_9313_44734# 0.145766f
C10635 a_n1741_47186# a_n971_45724# 0.157081f
C10636 a_n2109_47186# a_n237_47217# 0.730469f
C10637 a_n784_42308# a_1755_42282# 0.073102f
C10638 a_1067_42314# a_1184_42692# 0.147283f
C10639 a_17364_32525# VDD 0.511917f
C10640 a_4190_30871# VREF_GND 0.105109f
C10641 a_3905_42865# a_3539_42460# 0.022817f
C10642 a_7499_43078# a_9803_42558# 0.158876f
C10643 a_n2661_42282# a_n97_42460# 0.025699f
C10644 a_2324_44458# a_11691_44458# 0.045025f
C10645 a_13507_46334# a_20974_43370# 0.017855f
C10646 a_n357_42282# a_3537_45260# 0.200175f
C10647 a_12891_46348# a_12549_44172# 0.309821f
C10648 a_n971_45724# a_7832_46660# 0.013782f
C10649 a_2063_45854# a_10428_46928# 0.04306f
C10650 a_6491_46660# a_6540_46812# 0.079263f
C10651 a_n2312_39304# a_n2442_46660# 0.15211f
C10652 a_20974_43370# a_21855_43396# 0.029556f
C10653 a_14401_32519# a_13678_32519# 0.050672f
C10654 a_n97_42460# a_16823_43084# 0.205258f
C10655 a_5907_45546# VDD 0.390381f
C10656 a_n2956_37592# a_n3565_39304# 0.0261f
C10657 a_10193_42453# a_14539_43914# 0.278963f
C10658 a_526_44458# a_3905_42865# 0.321601f
C10659 a_3232_43370# a_6709_45028# 0.086072f
C10660 a_6171_45002# a_7229_43940# 0.010208f
C10661 a_10249_46116# a_11186_47026# 0.172467f
C10662 a_n881_46662# a_3147_46376# 0.073958f
C10663 a_n1613_43370# a_3483_46348# 0.029573f
C10664 a_16327_47482# a_18985_46122# 0.051538f
C10665 a_12861_44030# a_10809_44734# 0.156561f
C10666 a_4883_46098# a_10903_43370# 0.025531f
C10667 a_n4209_39304# VCM 0.05604f
C10668 a_n4334_38528# VDD 0.385889f
C10669 a_3726_37500# a_5088_37509# 0.189392f
C10670 a_n3420_39072# VIN_P 0.030377f
C10671 a_n3420_37984# C2_P_btm 0.03058f
C10672 a_n3565_39304# VREF 0.098117f
C10673 a_4520_42826# a_5111_42852# 0.047152f
C10674 a_9482_43914# a_15433_44458# 0.20244f
C10675 a_13556_45296# a_14815_43914# 0.378519f
C10676 a_11823_42460# a_14021_43940# 0.034191f
C10677 a_n2293_42834# a_n356_44636# 0.027771f
C10678 a_20447_31679# a_17730_32519# 0.051365f
C10679 a_19963_31679# a_19237_31679# 0.05162f
C10680 a_n2293_46098# a_3483_46348# 0.044283f
C10681 a_472_46348# a_1176_45822# 0.146555f
C10682 a_10227_46804# a_8696_44636# 0.089585f
C10683 a_n2497_47436# a_n913_45002# 0.019337f
C10684 a_14180_46812# a_10809_44734# 0.012862f
C10685 a_19237_31679# VDD 0.749539f
C10686 a_n3674_39304# a_n3674_38680# 0.17962f
C10687 a_n1741_47186# DATA[3] 0.033504f
C10688 a_n815_47178# DATA[0] 0.068508f
C10689 a_n23_47502# VDD 0.152616f
C10690 a_11415_45002# a_10907_45822# 0.050963f
C10691 a_2107_46812# a_1423_45028# 0.022467f
C10692 a_9145_43396# VDD 2.43736f
C10693 a_13259_45724# a_13575_42558# 0.097619f
C10694 a_3600_43914# a_3737_43940# 0.126609f
C10695 a_10490_45724# a_11652_45724# 0.044431f
C10696 a_11415_45002# a_21359_45002# 0.015551f
C10697 a_20202_43084# a_11827_44484# 0.032881f
C10698 a_18479_47436# a_19862_44208# 0.138185f
C10699 a_11322_45546# a_11525_45546# 0.055031f
C10700 a_13507_46334# a_12465_44636# 0.029101f
C10701 a_9313_45822# a_9804_47204# 0.171044f
C10702 a_12861_44030# a_n881_46662# 0.135351f
C10703 a_n971_45724# a_n743_46660# 0.122713f
C10704 a_n237_47217# a_n1925_46634# 0.079348f
C10705 a_15803_42450# a_16522_42674# 0.089677f
C10706 a_15959_42545# a_16104_42674# 0.057222f
C10707 a_19862_44208# a_4190_30871# 0.023868f
C10708 a_458_43396# a_648_43396# 0.045837f
C10709 a_3080_42308# a_2982_43646# 0.095684f
C10710 a_14180_46482# VDD 0.077608f
C10711 a_n2293_42834# a_n3674_38680# 0.010983f
C10712 a_742_44458# a_1793_42852# 0.010622f
C10713 a_15861_45028# a_16019_45002# 0.04712f
C10714 a_8696_44636# a_1307_43914# 0.030679f
C10715 a_n2840_45002# a_n2661_45010# 0.189331f
C10716 a_13507_46334# a_13887_32519# 0.08088f
C10717 a_3090_45724# a_7499_43940# 0.025901f
C10718 a_4791_45118# a_3483_46348# 0.088998f
C10719 a_4646_46812# a_6540_46812# 0.029952f
C10720 a_4651_46660# a_5732_46660# 0.102355f
C10721 a_3877_44458# a_5072_46660# 0.021873f
C10722 a_n1925_46634# a_8270_45546# 0.109762f
C10723 a_n881_46662# a_14180_46812# 0.028137f
C10724 a_n1741_47186# a_12594_46348# 0.150956f
C10725 a_21811_47423# a_21363_46634# 0.010128f
C10726 a_4883_46098# a_21188_46660# 0.012559f
C10727 a_4817_46660# a_5167_46660# 0.218775f
C10728 a_n2661_46634# a_11735_46660# 0.044956f
C10729 a_13747_46662# a_14976_45028# 0.016638f
C10730 a_11453_44696# a_20107_46660# 0.050203f
C10731 a_n1151_42308# a_5164_46348# 0.110485f
C10732 a_n3565_38502# a_n4064_37440# 0.028296f
C10733 a_n4064_38528# a_n3565_37414# 0.029213f
C10734 a_n3420_38528# a_n3420_37440# 0.051118f
C10735 a_16522_42674# VDD 0.077608f
C10736 a_n1059_45260# VDD 4.75361f
C10737 a_14579_43548# a_5534_30871# 0.030066f
C10738 a_13467_32519# a_14209_32519# 0.048306f
C10739 a_20556_43646# a_20749_43396# 0.018955f
C10740 a_19479_31679# VIN_N 0.028718f
C10741 a_3422_30871# a_1606_42308# 0.022481f
C10742 a_1423_45028# a_n2661_44458# 0.164701f
C10743 a_526_44458# a_4093_43548# 0.107158f
C10744 a_10903_43370# a_8685_43396# 0.031035f
C10745 a_20841_46902# a_20731_47026# 0.097745f
C10746 a_21363_46634# a_22000_46634# 0.017308f
C10747 a_20623_46660# a_20528_46660# 0.049827f
C10748 a_n1613_43370# a_n357_42282# 0.030838f
C10749 a_6755_46942# a_15015_46420# 0.133517f
C10750 a_4915_47217# a_13904_45546# 0.013453f
C10751 C8_N_btm VREF 3.6701f
C10752 C9_N_btm VIN_N 1.82823f
C10753 VDD EN_OFFSET_CAL 0.489629f
C10754 C7_N_btm VREF_GND 1.61142f
C10755 C6_N_btm VCM 0.877241f
C10756 a_n97_42460# a_13070_42354# 0.02477f
C10757 a_20447_31679# a_17538_32519# 0.051306f
C10758 a_15004_44636# a_14673_44172# 0.039287f
C10759 a_n863_45724# a_1847_42826# 0.216819f
C10760 a_n2312_39304# a_n3565_39304# 0.104981f
C10761 a_768_44030# a_6171_45002# 0.027851f
C10762 a_n2442_46660# a_n2810_45028# 0.045466f
C10763 a_n2438_43548# a_n2472_45002# 0.023014f
C10764 a_n2293_46098# a_n357_42282# 0.014918f
C10765 a_n1853_46287# a_n1099_45572# 0.067343f
C10766 a_n2497_47436# a_n2661_44458# 0.138848f
C10767 a_n2840_43370# VDD 0.246858f
C10768 a_7281_43914# a_7542_44172# 0.060549f
C10769 a_n1059_45260# a_16414_43172# 0.094309f
C10770 a_948_46660# VDD 0.278482f
C10771 a_10193_42453# a_19987_42826# 0.164153f
C10772 a_2324_44458# a_2437_43646# 0.011046f
C10773 a_15227_44166# a_16922_45042# 0.533576f
C10774 a_7903_47542# a_6575_47204# 0.046223f
C10775 a_6151_47436# a_11459_47204# 0.034818f
C10776 a_14097_32519# a_13258_32519# 0.051815f
C10777 en_comp COMP_P 1.91962f
C10778 a_17730_32519# a_13467_32519# 0.054292f
C10779 a_n2293_43922# a_12545_42858# 0.022686f
C10780 a_13925_46122# VDD 0.251868f
C10781 a_20512_43084# a_13678_32519# 0.059475f
C10782 a_18341_45572# a_18799_45938# 0.027606f
C10783 a_11652_45724# a_6171_45002# 0.072138f
C10784 a_10227_46804# a_14205_43396# 0.422372f
C10785 a_9049_44484# a_8953_45002# 0.031391f
C10786 a_4883_46098# a_8685_43396# 0.011038f
C10787 a_11599_46634# a_14976_45028# 0.020184f
C10788 a_4915_47217# a_14035_46660# 0.075669f
C10789 a_12861_44030# a_17609_46634# 0.183853f
C10790 a_n743_46660# a_601_46902# 0.022066f
C10791 a_n2438_43548# a_33_46660# 0.588568f
C10792 a_n133_46660# a_171_46873# 0.163873f
C10793 a_n1925_46634# a_1123_46634# 0.018809f
C10794 a_10227_46804# a_11813_46116# 0.094518f
C10795 a_n4209_39304# a_n4064_38528# 0.029379f
C10796 a_n3690_39392# a_n3690_38528# 0.050585f
C10797 a_1169_39043# comp_n 0.3874f
C10798 a_n3420_39072# a_n3565_38502# 0.034254f
C10799 a_n4064_39072# a_n4209_38502# 0.030674f
C10800 a_n3565_39304# a_n3420_38528# 0.028052f
C10801 a_1606_42308# VDD 0.629724f
C10802 a_15781_43660# a_15743_43084# 0.050751f
C10803 a_16409_43396# a_16977_43638# 0.17072f
C10804 a_16243_43396# a_17499_43370# 0.043633f
C10805 a_n356_44636# a_5379_42460# 0.038779f
C10806 a_n2956_37592# a_n3690_37440# 0.015408f
C10807 a_11967_42832# a_14635_42282# 0.018349f
C10808 a_18494_42460# a_18214_42558# 0.012583f
C10809 a_15599_45572# VDD 0.390565f
C10810 a_20447_31679# a_19721_31679# 0.070259f
C10811 a_4646_46812# a_7871_42858# 0.26422f
C10812 a_1823_45246# a_3080_42308# 0.049986f
C10813 a_15227_44166# a_15743_43084# 0.513622f
C10814 a_n743_46660# a_12594_46348# 0.0427f
C10815 a_n2661_46634# a_2324_44458# 0.0278f
C10816 a_4791_45118# a_n357_42282# 0.020355f
C10817 a_n443_46116# a_310_45028# 0.06667f
C10818 a_3090_45724# a_15227_46910# 0.010657f
C10819 a_15009_46634# a_13059_46348# 0.054389f
C10820 a_2107_46812# a_9569_46155# 0.018199f
C10821 a_11599_46634# a_18051_46116# 0.03664f
C10822 a_8912_37509# VDD 18.3523f
C10823 a_10890_34112# a_18194_34908# 0.419705f
C10824 VDAC_N RST_Z 0.154233f
C10825 a_n4318_40392# VDD 0.573389f
C10826 a_17333_42852# a_18249_42858# 0.311255f
C10827 a_18083_42858# a_18817_42826# 0.0532f
C10828 a_n443_42852# a_14579_43548# 0.04846f
C10829 a_11827_44484# a_n2661_42834# 0.046936f
C10830 a_13259_45724# a_16823_43084# 0.017563f
C10831 a_10227_46804# a_4958_30871# 0.036177f
C10832 SMPL_ON_N a_19963_31679# 0.029334f
C10833 a_8199_44636# a_2324_44458# 0.412215f
C10834 a_3090_45724# a_2957_45546# 0.167712f
C10835 a_18326_43940# VDD 0.129408f
C10836 a_14539_43914# a_14021_43940# 0.043922f
C10837 a_12465_44636# SINGLE_ENDED 0.067716f
C10838 a_4185_45028# a_4921_42308# 0.059648f
C10839 SMPL_ON_N VDD 0.497737f
C10840 a_n2312_38680# a_n4318_40392# 0.023897f
C10841 a_10586_45546# a_2711_45572# 0.295169f
C10842 a_8016_46348# a_8696_44636# 0.031525f
C10843 a_12891_46348# a_13076_44458# 0.182315f
C10844 a_768_44030# a_12607_44458# 0.215512f
C10845 a_3090_45724# a_9482_43914# 0.029795f
C10846 a_526_44458# a_7499_43078# 0.2203f
C10847 a_n1741_47186# a_n452_47436# 0.013149f
C10848 a_n2109_47186# a_n746_45260# 0.295988f
C10849 a_14209_32519# RST_Z 0.049869f
C10850 a_n784_42308# a_1606_42308# 15.027599f
C10851 a_1067_42314# a_1576_42282# 0.017282f
C10852 a_22959_43396# VDD 0.303237f
C10853 a_9313_44734# a_4361_42308# 0.082952f
C10854 a_3905_42865# a_3626_43646# 0.036343f
C10855 a_7499_43078# a_9223_42460# 0.013802f
C10856 a_n357_42282# a_13258_32519# 0.022774f
C10857 a_18451_43940# a_18797_44260# 0.013377f
C10858 a_n755_45592# a_3065_45002# 0.027852f
C10859 a_n1925_42282# a_n2661_43370# 0.027962f
C10860 a_17715_44484# a_11827_44484# 0.037803f
C10861 a_12465_44636# a_n743_46660# 0.026136f
C10862 a_6545_47178# a_6540_46812# 0.013617f
C10863 a_n2312_40392# a_n2442_46660# 5.91846f
C10864 a_n2312_39304# a_n2472_46634# 0.016291f
C10865 COMP_P a_22537_40625# 0.120662f
C10866 a_20974_43370# a_4361_42308# 0.122936f
C10867 a_17538_32519# a_13467_32519# 0.051209f
C10868 a_5891_43370# a_7309_42852# 0.071511f
C10869 a_5263_45724# VDD 0.202719f
C10870 a_n2810_45028# a_n3565_39304# 0.021534f
C10871 a_n1925_42282# a_2998_44172# 0.02835f
C10872 a_n1613_43370# a_8952_43230# 0.213002f
C10873 a_3232_43370# a_7229_43940# 0.180766f
C10874 a_6431_45366# a_5205_44484# 0.018787f
C10875 a_10249_46116# a_10768_47026# 0.027091f
C10876 a_n881_46662# a_2804_46116# 0.050669f
C10877 a_n1151_42308# a_5066_45546# 0.5423f
C10878 a_16327_47482# a_18819_46122# 0.324239f
C10879 a_13487_47204# a_6945_45028# 0.015556f
C10880 a_4883_46098# a_11387_46155# 0.010865f
C10881 a_11599_46634# a_19900_46494# 0.055271f
C10882 a_n4209_39304# VREF_GND 0.02097f
C10883 a_n4209_38502# VDD 0.817081f
C10884 a_3726_37500# a_4338_37500# 0.212154f
C10885 a_9482_43914# a_14815_43914# 0.024524f
C10886 a_n743_46660# a_2711_45572# 0.525746f
C10887 a_16327_47482# a_16223_45938# 0.016725f
C10888 a_472_46348# a_1208_46090# 0.088629f
C10889 a_n2497_47436# a_n1059_45260# 0.073215f
C10890 a_22959_44484# VDD 0.303517f
C10891 a_n1991_42858# a_n1736_42282# 0.0101f
C10892 a_12545_42858# a_12800_43218# 0.05936f
C10893 a_17730_32519# RST_Z 0.049818f
C10894 a_n2312_38680# a_n4209_38502# 0.095213f
C10895 a_n1741_47186# DATA[2] 0.017604f
C10896 a_7499_43078# a_8605_42826# 0.026478f
C10897 a_n237_47217# VDD 4.05131f
C10898 a_18494_42460# a_15493_43940# 0.02195f
C10899 a_11189_46129# a_2711_45572# 0.011492f
C10900 a_4646_46812# a_6709_45028# 0.031325f
C10901 a_4419_46090# a_4880_45572# 0.032829f
C10902 a_n971_45724# a_5891_43370# 0.084717f
C10903 a_5534_30871# a_n3420_38528# 0.041746f
C10904 a_19721_31679# a_13467_32519# 0.051394f
C10905 a_8270_45546# VDD 1.26092f
C10906 a_768_44030# a_5663_43940# 0.011502f
C10907 a_10193_42453# a_11962_45724# 0.044438f
C10908 a_n1613_43370# a_n1441_43940# 0.012196f
C10909 a_16327_47482# a_11341_43940# 0.063063f
C10910 a_11415_45002# a_21101_45002# 0.018873f
C10911 a_10809_44734# a_10951_45334# 0.015679f
C10912 a_10490_45724# a_11525_45546# 0.06936f
C10913 a_12741_44636# a_18494_42460# 0.114105f
C10914 a_9313_45822# a_8128_46384# 0.013269f
C10915 a_13717_47436# a_n881_46662# 0.039579f
C10916 a_21496_47436# a_4883_46098# 0.257837f
C10917 a_n746_45260# a_n1925_46634# 0.036469f
C10918 a_15764_42576# a_16522_42674# 0.05936f
C10919 a_n4318_37592# a_n4064_38528# 0.020352f
C10920 a_4093_43548# a_3626_43646# 0.011002f
C10921 a_15861_45028# a_15595_45028# 0.072432f
C10922 a_n2293_46634# a_9803_43646# 0.01299f
C10923 a_n443_46116# a_2804_46116# 0.018109f
C10924 a_3877_44458# a_6540_46812# 0.244975f
C10925 a_4646_46812# a_5732_46660# 0.050752f
C10926 a_4651_46660# a_5907_46634# 0.043482f
C10927 a_5807_45002# a_15368_46634# 0.029781f
C10928 a_4883_46098# a_21363_46634# 0.066909f
C10929 a_4817_46660# a_5385_46902# 0.170485f
C10930 a_13747_46662# a_3090_45724# 0.139869f
C10931 a_13661_43548# a_14976_45028# 0.162789f
C10932 a_13507_46334# a_22000_46634# 0.183978f
C10933 a_11453_44696# a_19551_46910# 0.047386f
C10934 a_n1151_42308# a_5068_46348# 0.089946f
C10935 a_n1741_47186# a_12005_46116# 0.174477f
C10936 a_7754_40130# a_7754_39964# 0.301877f
C10937 a_16104_42674# VDD 0.134357f
C10938 a_743_42282# a_20749_43396# 0.09037f
C10939 a_14579_43548# a_14543_43071# 0.032593f
C10940 a_13678_32519# a_5649_42852# 0.506367f
C10941 a_3357_43084# CLK 2.63944f
C10942 a_n2017_45002# VDD 3.8321f
C10943 a_n2293_43922# a_12563_42308# 0.015547f
C10944 a_n971_45724# a_n3674_37592# 0.022388f
C10945 a_526_44458# a_1756_43548# 0.01292f
C10946 a_n881_46662# a_n1099_45572# 0.088565f
C10947 a_21363_46634# a_21188_46660# 0.233657f
C10948 a_20273_46660# a_20731_47026# 0.027606f
C10949 a_2063_45854# a_10907_45822# 0.22153f
C10950 C7_N_btm VREF 1.818f
C10951 C8_N_btm VIN_N 0.907642f
C10952 VDD DATA[5] 0.504354f
C10953 C6_N_btm VREF_GND 0.836236f
C10954 C5_N_btm VCM 0.719982f
C10955 a_3422_30871# VDAC_N 0.480156f
C10956 a_2711_45572# a_4361_42308# 0.031943f
C10957 a_n2293_42834# a_3499_42826# 0.029158f
C10958 a_n863_45724# a_791_42968# 0.338631f
C10959 a_14537_43396# a_11341_43940# 0.032289f
C10960 a_5891_43370# a_9313_44734# 0.028253f
C10961 a_n2293_46098# a_310_45028# 0.017313f
C10962 a_12549_44172# a_6171_45002# 0.029809f
C10963 a_768_44030# a_3232_43370# 0.224083f
C10964 a_6755_46942# a_15765_45572# 0.026052f
C10965 a_2107_46812# a_3357_43084# 0.033995f
C10966 a_n2293_46634# a_n913_45002# 0.024406f
C10967 a_15368_46634# a_15143_45578# 0.105334f
C10968 a_n2438_43548# a_n2661_45010# 0.220364f
C10969 a_n4318_38680# a_n4064_39616# 0.021342f
C10970 a_17538_32519# RST_Z 0.050782f
C10971 a_4190_30871# a_n3420_38528# 0.031855f
C10972 a_n913_45002# a_5342_30871# 0.122483f
C10973 a_n1059_45260# a_15567_42826# 0.048229f
C10974 a_1123_46634# VDD 0.469393f
C10975 a_13507_46334# a_20512_43084# 0.497215f
C10976 a_3090_45724# a_18911_45144# 0.190188f
C10977 a_13661_43548# a_15433_44458# 0.038412f
C10978 a_12549_44172# a_14673_44172# 0.024138f
C10979 a_11415_45002# a_14797_45144# 0.021281f
C10980 a_8049_45260# a_15765_45572# 0.012841f
C10981 a_5257_43370# a_5518_44484# 0.095452f
C10982 a_4915_47217# a_n1435_47204# 0.038318f
C10983 a_7227_47204# a_6575_47204# 0.028925f
C10984 a_6151_47436# a_9313_45822# 0.032544f
C10985 a_22400_42852# a_13258_32519# 0.039834f
C10986 a_5934_30871# a_8515_42308# 0.222946f
C10987 en_comp a_n4318_37592# 0.03345f
C10988 a_n2293_43922# a_12089_42308# 0.183316f
C10989 a_13759_46122# VDD 0.399995f
C10990 a_20512_43084# a_21855_43396# 0.013929f
C10991 a_3422_30871# a_14209_32519# 0.031148f
C10992 a_n2017_45002# a_n784_42308# 0.0226f
C10993 a_18341_45572# a_18596_45572# 0.056391f
C10994 a_18909_45814# a_19256_45572# 0.051162f
C10995 a_10227_46804# a_14358_43442# 0.019948f
C10996 a_20202_43084# a_19279_43940# 0.020761f
C10997 a_9290_44172# a_9313_44734# 0.140741f
C10998 a_16327_47482# a_10341_43396# 0.159266f
C10999 a_11599_46634# a_3090_45724# 0.133107f
C11000 a_4915_47217# a_13885_46660# 0.179458f
C11001 a_12861_44030# a_16292_46812# 0.059827f
C11002 a_n743_46660# a_33_46660# 0.025563f
C11003 a_n2438_43548# a_171_46873# 0.029723f
C11004 a_10227_46804# a_11735_46660# 0.54163f
C11005 a_n4209_39590# a_n4064_37984# 0.032388f
C11006 a_1169_39043# a_1666_39043# 0.08488f
C11007 a_n2302_39072# a_n2216_39072# 0.011479f
C11008 a_n4064_39616# a_n4209_38216# 0.027937f
C11009 a_n3420_39616# a_n3565_38216# 0.028042f
C11010 a_n3565_39590# a_n3420_37984# 0.031465f
C11011 a_5934_30871# EN_VIN_BSTR_N 0.073476f
C11012 a_16243_43396# a_16759_43396# 0.106647f
C11013 a_2479_44172# a_n2293_42282# 0.059476f
C11014 a_n2956_37592# a_n3565_37414# 0.304738f
C11015 a_11967_42832# a_13291_42460# 0.015813f
C11016 a_18494_42460# a_19332_42282# 0.040916f
C11017 a_18184_42460# a_18214_42558# 0.056496f
C11018 a_20447_31679# a_18114_32519# 0.051474f
C11019 a_3357_43084# a_n2661_44458# 0.027126f
C11020 a_4646_46812# a_7227_42852# 0.032378f
C11021 a_n443_46116# a_n1099_45572# 0.368941f
C11022 a_n743_46660# a_12005_46116# 0.024033f
C11023 a_n881_46662# a_n1925_42282# 0.041426f
C11024 a_15009_46634# a_15227_46910# 0.08213f
C11025 a_3877_44458# a_1823_45246# 0.231164f
C11026 a_2107_46812# a_9625_46129# 0.184645f
C11027 a_n4209_37414# VCM 0.03628f
C11028 a_n3565_37414# VREF 0.046045f
C11029 a_n3420_37440# VIN_P 0.137523f
C11030 VDAC_N VDD 4.61811f
C11031 a_6886_37412# RST_Z 0.031637f
C11032 a_10890_34112# EN_VIN_BSTR_N 1.06104f
C11033 a_19721_31679# RST_Z 0.050546f
C11034 a_18083_42858# a_18249_42858# 0.699797f
C11035 a_n2840_44458# VDD 0.247948f
C11036 a_n443_42852# a_13667_43396# 0.035517f
C11037 a_12883_44458# a_13076_44458# 0.142643f
C11038 a_12607_44458# a_13720_44458# 0.122704f
C11039 a_16388_46812# a_16375_45002# 0.039999f
C11040 a_18597_46090# a_n913_45002# 0.126328f
C11041 a_11453_44696# a_3357_43084# 0.020072f
C11042 a_18079_43940# VDD 0.162408f
C11043 a_12465_44636# START 0.065727f
C11044 a_n2661_42834# a_n2661_42282# 0.019795f
C11045 a_20447_31679# a_13887_32519# 0.051465f
C11046 a_n913_45002# a_743_42282# 0.25834f
C11047 a_9313_44734# a_10807_43548# 0.033005f
C11048 a_22731_47423# VDD 0.196667f
C11049 a_19963_31679# a_14209_32519# 0.051256f
C11050 a_14537_43396# a_10341_43396# 0.013753f
C11051 a_21811_47423# SINGLE_ENDED 0.215228f
C11052 a_n2840_45546# a_n2661_45546# 0.175179f
C11053 a_n2293_46634# a_n2661_44458# 0.029279f
C11054 a_12549_44172# a_12607_44458# 0.033279f
C11055 a_12891_46348# a_12883_44458# 0.018059f
C11056 a_8270_45546# a_1423_45028# 0.023554f
C11057 a_768_44030# a_8975_43940# 0.124155f
C11058 a_4190_30871# VIN_N 0.049977f
C11059 SMPL_ON_P a_n1605_47204# 0.194856f
C11060 a_n1741_47186# a_n815_47178# 0.031488f
C11061 a_n2109_47186# a_n971_45724# 1.21934f
C11062 a_14209_32519# VDD 0.284895f
C11063 a_9313_44734# a_13467_32519# 0.057668f
C11064 a_2107_46812# a_9672_43914# 0.079349f
C11065 a_13259_45724# a_14797_45144# 0.092924f
C11066 a_n357_42282# a_3065_45002# 0.023226f
C11067 a_3316_45546# a_413_45260# 0.110075f
C11068 a_3483_46348# a_6298_44484# 0.017162f
C11069 a_16327_47482# a_n97_42460# 0.113034f
C11070 a_19321_45002# a_15493_43940# 0.050579f
C11071 a_5907_45546# a_3357_43084# 0.023698f
C11072 a_526_44458# a_n2661_43370# 0.054473f
C11073 a_2063_45854# a_9863_46634# 0.10786f
C11074 a_6151_47436# a_6540_46812# 0.043688f
C11075 a_n2312_39304# a_n2661_46634# 0.105298f
C11076 a_n784_42308# VDAC_N 0.010218f
C11077 COMP_P a_22589_40599# 0.204694f
C11078 a_20974_43370# a_13467_32519# 0.017399f
C11079 a_5891_43370# a_5837_42852# 0.010625f
C11080 a_4099_45572# VDD 0.296272f
C11081 en_comp a_1273_38525# 0.03792f
C11082 a_n2956_37592# a_n4209_39304# 0.102982f
C11083 a_8696_44636# a_11827_44484# 0.039f
C11084 a_526_44458# a_2998_44172# 0.028337f
C11085 a_10903_43370# a_12429_44172# 0.116356f
C11086 a_n1613_43370# a_9127_43156# 0.267842f
C11087 a_3232_43370# a_7276_45260# 0.027376f
C11088 a_6171_45002# a_5205_44484# 0.0168f
C11089 a_10467_46802# a_11735_46660# 0.096658f
C11090 a_10554_47026# a_10768_47026# 0.097745f
C11091 a_10623_46897# a_11186_47026# 0.049827f
C11092 a_n881_46662# a_2698_46116# 0.058407f
C11093 a_13507_46334# a_10903_43370# 0.016027f
C11094 a_19321_45002# a_12741_44636# 0.113088f
C11095 a_12861_44030# a_6945_45028# 0.108969f
C11096 a_10227_46804# a_2324_44458# 0.051051f
C11097 a_11599_46634# a_20075_46420# 0.021805f
C11098 a_20916_46384# a_20202_43084# 0.181561f
C11099 a_2112_39137# VDD 0.28506f
C11100 a_n4209_39304# VREF 0.195875f
C11101 a_n3565_38216# C2_P_btm 0.040789f
C11102 a_n3565_39304# VIN_P 0.038656f
C11103 a_3935_42891# a_4520_42826# 0.017436f
C11104 a_13556_45296# a_13857_44734# 0.01375f
C11105 a_19963_31679# a_17730_32519# 0.054244f
C11106 a_n357_42282# a_458_43396# 0.016095f
C11107 a_n755_45592# a_n229_43646# 0.049717f
C11108 a_768_44030# a_10193_42453# 0.030504f
C11109 a_472_46348# a_805_46414# 0.360492f
C11110 a_1209_47178# a_2437_43646# 0.025116f
C11111 a_n2497_47436# a_n2017_45002# 0.125552f
C11112 a_13885_46660# a_10809_44734# 0.026009f
C11113 a_17730_32519# VDD 0.291149f
C11114 a_3626_43646# a_7174_31319# 0.022247f
C11115 a_10922_42852# a_11136_42852# 0.097745f
C11116 a_12089_42308# a_12800_43218# 0.15794f
C11117 a_743_42282# a_1755_42282# 0.058846f
C11118 a_n746_45260# VDD 1.41433f
C11119 a_7499_43078# a_8037_42858# 0.160087f
C11120 a_n1741_47186# DATA[1] 0.021536f
C11121 a_18184_42460# a_15493_43940# 0.022388f
C11122 a_9290_44172# a_2711_45572# 0.030631f
C11123 a_4646_46812# a_7229_43940# 0.104864f
C11124 a_4190_30871# CAL_N 0.045535f
C11125 a_18114_32519# a_13467_32519# 0.055508f
C11126 a_6755_46942# CLK 0.031541f
C11127 a_768_44030# a_5495_43940# 0.017815f
C11128 a_10809_44734# a_10775_45002# 0.022389f
C11129 a_2324_44458# a_1307_43914# 0.129761f
C11130 a_10193_42453# a_11652_45724# 0.197229f
C11131 a_11415_45002# a_21005_45260# 0.01592f
C11132 a_15227_44166# a_17767_44458# 0.023473f
C11133 a_10490_45724# a_11322_45546# 0.246478f
C11134 a_12741_44636# a_18184_42460# 0.041879f
C11135 a_n1925_42282# a_3537_45260# 0.055426f
C11136 a_18597_46090# a_11453_44696# 0.022871f
C11137 a_9863_47436# a_9804_47204# 0.109361f
C11138 a_n1435_47204# a_n881_46662# 0.068194f
C11139 a_13507_46334# a_4883_46098# 4.09671f
C11140 a_n971_45724# a_n1925_46634# 0.163523f
C11141 a_15764_42576# a_16104_42674# 0.029366f
C11142 a_14021_43940# a_17499_43370# 0.011011f
C11143 a_8049_45260# CLK 0.033207f
C11144 a_n2017_45002# a_15764_42576# 0.014981f
C11145 a_13507_46334# a_5649_42852# 0.136078f
C11146 a_n2293_46634# a_9145_43396# 0.238561f
C11147 a_n443_46116# a_2698_46116# 0.012019f
C11148 a_3877_44458# a_5732_46660# 0.040487f
C11149 a_4646_46812# a_5907_46634# 0.037052f
C11150 a_4651_46660# a_5167_46660# 0.102946f
C11151 a_16327_47482# a_11415_45002# 0.94171f
C11152 a_13661_43548# a_3090_45724# 0.177565f
C11153 a_5807_45002# a_14976_45028# 0.026261f
C11154 a_13507_46334# a_21188_46660# 0.03408f
C11155 a_11453_44696# a_19123_46287# 0.021733f
C11156 a_n1741_47186# a_10903_43370# 0.066687f
C11157 a_n3565_38502# a_n3420_37440# 0.034147f
C11158 a_n4209_38502# a_n4064_37440# 0.028279f
C11159 a_n4064_38528# a_n4209_37414# 0.027936f
C11160 a_n3420_38528# a_n3565_37414# 0.029229f
C11161 a_3754_39964# VDAC_Pi 0.296508f
C11162 a_21855_43396# a_5649_42852# 0.057783f
C11163 a_13467_32519# a_13887_32519# 0.058303f
C11164 a_n2109_45247# VDD 0.266396f
C11165 a_8953_45002# a_9838_44484# 0.013986f
C11166 a_n467_45028# a_n23_44458# 0.038286f
C11167 a_626_44172# a_n2661_44458# 0.031248f
C11168 a_526_44458# a_1568_43370# 0.220609f
C11169 a_8953_45546# a_9803_43646# 0.091141f
C11170 a_n971_45724# a_n327_42558# 0.01976f
C11171 a_n443_42852# a_15493_43396# 0.025952f
C11172 a_n1613_43370# a_n1099_45572# 0.025553f
C11173 a_18285_46348# a_18280_46660# 0.089884f
C11174 a_20273_46660# a_20528_46660# 0.056391f
C11175 a_9313_45822# a_9049_44484# 0.119007f
C11176 a_3090_45724# a_4185_45028# 0.770164f
C11177 a_2107_46812# a_8049_45260# 0.029889f
C11178 a_13059_46348# a_12741_44636# 0.02008f
C11179 C6_N_btm VREF 1.41944f
C11180 C7_N_btm VIN_N 1.52449f
C11181 VDD DATA[4] 0.326957f
C11182 C5_N_btm VREF_GND 0.676559f
C11183 C4_N_btm VCM 0.716447f
C11184 a_n97_42460# a_11633_42558# 0.011546f
C11185 a_n13_43084# a_133_42852# 0.171361f
C11186 a_3626_43646# a_5932_42308# 0.062334f
C11187 a_n356_44636# a_n2293_43922# 0.025509f
C11188 a_3537_45260# a_3737_43940# 0.012872f
C11189 a_18114_32519# a_22315_44484# 0.017551f
C11190 a_20447_31679# a_14401_32519# 0.054145f
C11191 a_19963_31679# a_17538_32519# 0.051095f
C11192 a_n863_45724# a_685_42968# 0.052365f
C11193 a_n2312_39304# a_n4209_39304# 0.19527f
C11194 a_n2956_39768# a_n2956_37592# 0.047483f
C11195 a_n2293_46098# a_n1099_45572# 0.069723f
C11196 a_n1853_46287# a_n452_45724# 0.080546f
C11197 a_12891_46348# a_6171_45002# 0.040434f
C11198 a_6755_46942# a_15903_45785# 0.192397f
C11199 a_n2293_46634# a_n1059_45260# 0.051525f
C11200 a_10903_43370# a_10586_45546# 0.238199f
C11201 a_17538_32519# VDD 0.352922f
C11202 a_n3674_39304# a_n4064_39616# 0.020873f
C11203 a_383_46660# VDD 0.198466f
C11204 a_n1059_45260# a_5342_30871# 0.030512f
C11205 a_n357_42282# a_14635_42282# 0.010701f
C11206 a_18579_44172# a_19862_44208# 0.091151f
C11207 a_n356_44636# a_n97_42460# 1.46232f
C11208 a_22612_30879# VCM 0.473529f
C11209 a_5257_43370# a_5343_44458# 0.063407f
C11210 a_8953_45546# a_n913_45002# 0.052161f
C11211 a_3090_45724# a_18587_45118# 0.039584f
C11212 a_13661_43548# a_14815_43914# 0.060575f
C11213 a_3218_45724# a_3260_45572# 0.010055f
C11214 a_11415_45002# a_14537_43396# 0.04406f
C11215 a_12741_44636# a_13556_45296# 0.046411f
C11216 a_4915_47217# a_13381_47204# 0.045103f
C11217 a_6851_47204# a_6575_47204# 0.027563f
C11218 a_6151_47436# a_11031_47542# 0.03901f
C11219 a_n1741_47186# a_4883_46098# 0.031761f
C11220 a_n2293_43922# a_12379_42858# 0.030458f
C11221 a_20512_43084# a_4361_42308# 0.02826f
C11222 a_n2956_37592# a_n4318_37592# 0.023082f
C11223 a_n2017_45002# a_196_42282# 0.010023f
C11224 a_13351_46090# VDD 0.238036f
C11225 a_18479_45785# a_18596_45572# 0.183223f
C11226 a_18341_45572# a_19256_45572# 0.116691f
C11227 a_10227_46804# a_14579_43548# 0.118896f
C11228 a_11322_45546# a_6171_45002# 0.069025f
C11229 w_10694_33990# a_17364_32525# 0.017447f
C11230 a_n2442_46660# a_n4318_39304# 0.023691f
C11231 a_11453_44696# a_6755_46942# 0.026496f
C11232 a_n2438_43548# a_n133_46660# 0.848709f
C11233 a_12861_44030# a_15559_46634# 0.066578f
C11234 a_n743_46660# a_171_46873# 0.075858f
C11235 a_768_44030# a_4646_46812# 0.047094f
C11236 a_10227_46804# a_11186_47026# 0.018916f
C11237 a_n4209_39304# a_n3420_38528# 0.029412f
C11238 a_n3565_39304# a_n3565_38502# 0.041674f
C11239 a_n3420_39072# a_n4209_38502# 0.032647f
C11240 a_n2661_42834# a_n4318_38216# 0.023647f
C11241 a_16243_43396# a_16977_43638# 0.053479f
C11242 a_16547_43609# a_16409_43396# 0.206231f
C11243 a_4905_42826# a_5111_42852# 0.105155f
C11244 a_18494_42460# a_18907_42674# 0.11494f
C11245 a_18184_42460# a_19332_42282# 0.042769f
C11246 a_n2810_45028# a_n3565_37414# 0.135518f
C11247 a_8953_45002# a_n2661_43370# 0.034058f
C11248 a_1823_45246# a_4235_43370# 0.029154f
C11249 a_n913_45002# a_20193_45348# 0.224918f
C11250 a_19963_31679# a_19721_31679# 9.01086f
C11251 a_n443_46116# a_380_45546# 0.073277f
C11252 a_n2109_47186# a_2711_45572# 0.032969f
C11253 a_11453_44696# a_8049_45260# 0.032046f
C11254 a_16327_47482# a_13259_45724# 0.584328f
C11255 a_19321_45002# a_18985_46122# 0.019556f
C11256 a_n743_46660# a_10903_43370# 0.080542f
C11257 a_n881_46662# a_526_44458# 0.060324f
C11258 a_5700_37509# RST_Z 0.051902f
C11259 a_6886_37412# VDD 0.235486f
C11260 a_18083_42858# a_17333_42852# 0.284837f
C11261 a_18114_32519# RST_Z 0.049686f
C11262 a_19721_31679# VDD 0.527265f
C11263 a_n443_42852# a_10695_43548# 0.042055f
C11264 a_742_44458# a_n356_44636# 0.207503f
C11265 a_12607_44458# a_13076_44458# 0.200168f
C11266 a_8016_46348# a_2324_44458# 0.048711f
C11267 a_11189_46129# a_10903_43370# 0.151119f
C11268 a_n2293_46098# a_n1925_42282# 0.020467f
C11269 a_17973_43940# VDD 0.265874f
C11270 a_5342_30871# a_1606_42308# 0.023615f
C11271 a_19479_31679# a_17364_32525# 0.05375f
C11272 a_4223_44672# a_7499_43940# 0.030206f
C11273 a_n1059_45260# a_743_42282# 0.198704f
C11274 a_4883_46098# SINGLE_ENDED 0.1664f
C11275 a_22223_47212# VDD 0.236555f
C11276 a_22315_44484# a_22485_44484# 0.109468f
C11277 a_n2840_45546# a_n2810_45572# 0.162234f
C11278 a_12891_46348# a_12607_44458# 0.067773f
C11279 a_768_44030# a_10057_43914# 0.041949f
C11280 a_4190_30871# VIN_P 0.049977f
C11281 a_13887_32519# RST_Z 0.048316f
C11282 a_n1741_47186# a_n1605_47204# 0.011722f
C11283 a_n2109_47186# a_n452_47436# 0.039314f
C11284 a_n2497_47436# a_n746_45260# 0.046973f
C11285 a_22591_43396# VDD 0.280354f
C11286 a_n357_42282# a_19511_42282# 0.056757f
C11287 a_2382_45260# a_n2293_42282# 0.080755f
C11288 a_20731_47026# VDD 0.132317f
C11289 a_8953_45546# a_n2661_44458# 0.019448f
C11290 a_2107_46812# a_9028_43914# 0.110155f
C11291 a_13259_45724# a_14537_43396# 0.083218f
C11292 a_3218_45724# a_413_45260# 0.016434f
C11293 a_13904_45546# a_14127_45572# 0.011458f
C11294 a_3483_46348# a_5518_44484# 0.081879f
C11295 a_n2661_45546# a_3232_43370# 0.038743f
C11296 a_3090_45724# a_11967_42832# 0.12811f
C11297 a_n1151_42308# a_7715_46873# 0.09029f
C11298 a_4883_46098# a_n743_46660# 5.6639f
C11299 a_n2312_39304# a_n2956_39768# 5.91067f
C11300 a_22775_42308# a_22485_38105# 0.330766f
C11301 a_7309_42852# VDD 0.177437f
C11302 a_n2810_45028# a_n4209_39304# 0.021684f
C11303 a_21381_43940# a_4361_42308# 0.195418f
C11304 a_14401_32519# a_13467_32519# 0.050489f
C11305 a_3175_45822# VDD 0.193907f
C11306 a_10903_43370# a_11750_44172# 0.135933f
C11307 a_n1613_43370# a_8387_43230# 0.163582f
C11308 a_6171_45002# a_6431_45366# 0.017465f
C11309 a_3232_43370# a_5205_44484# 0.217288f
C11310 a_n2956_38680# a_n3674_39768# 0.023133f
C11311 a_11599_46634# a_19335_46494# 0.030852f
C11312 a_10467_46802# a_11186_47026# 0.082642f
C11313 a_10623_46897# a_10768_47026# 0.057222f
C11314 a_n881_46662# a_2521_46116# 0.050613f
C11315 a_16327_47482# a_18189_46348# 0.029513f
C11316 a_5257_43370# a_3090_45724# 0.020885f
C11317 a_n443_46116# a_526_44458# 0.366438f
C11318 a_13717_47436# a_6945_45028# 0.038878f
C11319 a_10227_46804# a_14840_46494# 0.275527f
C11320 a_n2312_40392# COMP_P 0.035637f
C11321 a_n2312_39304# a_n4318_37592# 0.023445f
C11322 a_9482_43914# a_13857_44734# 0.011887f
C11323 a_19479_31679# a_19237_31679# 9.049419f
C11324 a_2711_45572# a_19319_43548# 0.225335f
C11325 a_12549_44172# a_10193_42453# 0.116594f
C11326 a_n237_47217# a_3357_43084# 0.022871f
C11327 a_16327_47482# a_17478_45572# 0.012405f
C11328 a_n1925_46634# a_2711_45572# 0.030736f
C11329 a_12379_42858# a_12800_43218# 0.089677f
C11330 a_10991_42826# a_11136_42852# 0.057222f
C11331 a_743_42282# a_1606_42308# 0.088097f
C11332 a_22591_44484# VDD 0.223346f
C11333 a_3537_45260# a_3539_42460# 0.264936f
C11334 a_9313_44734# a_3422_30871# 0.043499f
C11335 a_19778_44110# a_15493_43940# 0.033844f
C11336 a_18494_42460# a_11341_43940# 0.025825f
C11337 a_n971_45724# VDD 4.911799f
C11338 SMPL_ON_P CLK_DATA 0.200962f
C11339 a_n2109_47186# DATA[2] 0.05382f
C11340 a_n1741_47186# DATA[0] 0.051737f
C11341 a_4646_46812# a_7276_45260# 0.016809f
C11342 a_10249_46116# CLK 0.063525f
C11343 a_3422_30871# a_20974_43370# 0.020902f
C11344 a_n2956_38680# a_n4315_30879# 0.024632f
C11345 a_768_44030# a_5013_44260# 0.064017f
C11346 a_11415_45002# a_20567_45036# 0.011165f
C11347 a_10193_42453# a_11525_45546# 0.0979f
C11348 a_167_45260# a_n2661_43370# 0.055202f
C11349 a_15227_44166# a_16979_44734# 0.181002f
C11350 a_3090_45724# a_18989_43940# 0.095784f
C11351 a_12741_44636# a_19778_44110# 0.070586f
C11352 a_526_44458# a_3537_45260# 0.938783f
C11353 a_n1151_42308# a_13747_46662# 0.050569f
C11354 a_13381_47204# a_n881_46662# 0.025748f
C11355 a_13507_46334# a_21496_47436# 0.167302f
C11356 a_n3674_38216# a_n4064_38528# 0.020875f
C11357 a_n4318_37592# a_n3420_38528# 0.024768f
C11358 a_n913_45002# a_14113_42308# 0.029759f
C11359 a_13507_46334# a_13678_32519# 0.037522f
C11360 a_13259_45724# a_n356_44636# 0.026337f
C11361 a_1823_45246# a_3905_42865# 0.218008f
C11362 a_n755_45592# a_5343_44458# 0.349527f
C11363 a_3877_44458# a_5907_46634# 0.073504f
C11364 a_4646_46812# a_5167_46660# 0.033486f
C11365 a_4651_46660# a_5385_46902# 0.053479f
C11366 a_16327_47482# a_20202_43084# 0.475502f
C11367 a_4955_46873# a_4817_46660# 0.318259f
C11368 a_n2293_46634# a_8270_45546# 0.030248f
C11369 a_13507_46334# a_21363_46634# 0.029223f
C11370 a_11453_44696# a_18285_46348# 0.236771f
C11371 a_13747_46662# a_14084_46812# 0.038349f
C11372 a_5807_45002# a_3090_45724# 0.032418f
C11373 a_n2293_45010# VDD 1.885f
C11374 a_4190_30871# a_20749_43396# 0.018962f
C11375 a_n356_44636# a_18057_42282# 0.087032f
C11376 a_4361_42308# a_5649_42852# 0.064476f
C11377 a_21855_43396# a_13678_32519# 0.17881f
C11378 a_3357_43084# DATA[5] 0.032568f
C11379 a_n467_45028# a_n356_44636# 0.052527f
C11380 a_526_44458# a_1049_43396# 0.121121f
C11381 a_8953_45546# a_9145_43396# 0.019849f
C11382 a_18479_45785# a_17517_44484# 0.023114f
C11383 SMPL_ON_P a_n1794_35082# 6.16983f
C11384 a_20411_46873# a_20528_46660# 0.170785f
C11385 a_20841_46902# a_21188_46660# 0.051162f
C11386 a_13747_46662# a_19240_46482# 0.012097f
C11387 C5_N_btm VREF 0.987144f
C11388 C6_N_btm VIN_N 0.391905f
C11389 VDD DATA[3] 0.309692f
C11390 C4_N_btm VREF_GND 0.671882f
C11391 C3_N_btm VCM 0.716273f
C11392 a_9313_44734# VDD 0.389068f
C11393 a_n97_42460# a_11551_42558# 0.095523f
C11394 a_n356_44636# a_n2661_43922# 0.041936f
C11395 w_1575_34786# VDAC_P 0.107674f
C11396 a_3090_45724# a_15143_45578# 0.016572f
C11397 a_n1853_46287# a_n863_45724# 0.019522f
C11398 a_6755_46942# a_15599_45572# 0.024601f
C11399 a_n2293_46634# a_n2017_45002# 0.039556f
C11400 a_n2956_39768# a_n2810_45028# 0.04304f
C11401 a_1983_46706# a_2437_43646# 0.01301f
C11402 a_n4318_38680# a_n3420_39616# 0.02534f
C11403 a_20974_43370# VDD 0.550101f
C11404 a_14401_32519# RST_Z 0.048069f
C11405 a_601_46902# VDD 0.204253f
C11406 a_n2017_45002# a_5342_30871# 0.038471f
C11407 a_n913_45002# a_5534_30871# 0.274894f
C11408 a_n1059_45260# a_15279_43071# 0.021145f
C11409 a_18494_42460# a_10341_43396# 0.030934f
C11410 a_18579_44172# a_19478_44306# 0.040429f
C11411 a_22612_30879# VREF_GND 0.168163f
C11412 a_21588_30879# VCM 0.179761f
C11413 a_8953_45546# a_n1059_45260# 0.318691f
C11414 a_3090_45724# a_18315_45260# 0.061731f
C11415 a_12741_44636# a_9482_43914# 0.101234f
C11416 a_11415_45002# a_14180_45002# 0.025987f
C11417 a_6491_46660# a_6575_47204# 0.029984f
C11418 a_4915_47217# a_11459_47204# 0.03966f
C11419 a_6151_47436# a_9863_47436# 0.030884f
C11420 a_n1151_42308# a_11599_46634# 0.116147f
C11421 a_20512_43084# a_13467_32519# 0.021245f
C11422 a_3422_30871# a_13887_32519# 0.031713f
C11423 en_comp a_n3674_38216# 0.026738f
C11424 a_n2810_45028# a_n4318_37592# 0.023097f
C11425 a_n2017_45002# a_n473_42460# 0.017082f
C11426 a_12594_46348# VDD 1.03351f
C11427 a_18175_45572# a_18596_45572# 0.086708f
C11428 a_18341_45572# a_19431_45546# 0.041762f
C11429 a_18909_45814# a_18691_45572# 0.209641f
C11430 a_18479_45785# a_19256_45572# 0.044595f
C11431 a_n863_45724# a_n2661_43370# 0.076347f
C11432 a_n743_46660# a_n133_46660# 0.205551f
C11433 a_12861_44030# a_15368_46634# 0.066698f
C11434 a_768_44030# a_3877_44458# 0.012394f
C11435 a_10227_46804# a_10768_47026# 0.012196f
C11436 a_6123_31319# EN_VIN_BSTR_N 0.050716f
C11437 a_n4209_39590# a_n3420_37984# 0.032713f
C11438 a_n3420_39616# a_n4209_38216# 0.027924f
C11439 a_n3565_39590# a_n3565_38216# 0.031123f
C11440 a_961_42354# VDD 0.091526f
C11441 a_16243_43396# a_16409_43396# 0.575934f
C11442 a_n2956_37592# a_n4209_37414# 0.145558f
C11443 a_18184_42460# a_18907_42674# 0.071964f
C11444 a_18494_42460# a_18727_42674# 0.031761f
C11445 a_15037_45618# VDD 0.08759f
C11446 a_4905_42826# a_4520_42826# 0.147708f
C11447 a_8191_45002# a_n2661_43370# 0.013381f
C11448 a_10193_42453# a_17061_44734# 0.012286f
C11449 a_1823_45246# a_4093_43548# 0.17443f
C11450 a_19963_31679# a_18114_32519# 0.051445f
C11451 a_2905_45572# a_3218_45724# 0.021505f
C11452 a_n237_47217# a_2277_45546# 0.104529f
C11453 a_n443_46116# a_n452_45724# 0.188857f
C11454 a_19321_45002# a_18819_46122# 0.018323f
C11455 a_n881_46662# a_2981_46116# 0.026038f
C11456 a_n1613_43370# a_526_44458# 0.826565f
C11457 a_2107_46812# a_5937_45572# 0.027091f
C11458 a_11599_46634# a_19240_46482# 0.016662f
C11459 VDAC_N C10_N_btm 0.883474p
C11460 a_5088_37509# RST_Z 0.059771f
C11461 a_n4209_37414# VREF 0.056254f
C11462 a_n3565_37414# VIN_P 0.028947f
C11463 a_5700_37509# VDD 1.0734f
C11464 a_17701_42308# a_17333_42852# 0.061051f
C11465 a_18114_32519# VDD 0.552219f
C11466 a_n443_42852# a_9803_43646# 0.102893f
C11467 a_n452_44636# a_n356_44636# 0.318214f
C11468 a_12607_44458# a_12883_44458# 0.11453f
C11469 a_n971_45724# a_1423_45028# 0.021147f
C11470 a_3090_45724# a_n755_45592# 0.051041f
C11471 a_9290_44172# a_10903_43370# 0.340316f
C11472 a_11189_46129# a_11387_46155# 0.320331f
C11473 a_12549_44172# a_18479_45785# 0.105486f
C11474 a_n2293_46098# a_526_44458# 0.053029f
C11475 SMPL_ON_N a_19479_31679# 0.029207f
C11476 a_17737_43940# VDD 0.285511f
C11477 a_4223_44672# a_6671_43940# 0.03251f
C11478 a_n2017_45002# a_743_42282# 7.84646f
C11479 a_19963_31679# a_13887_32519# 0.051213f
C11480 a_n913_45002# a_4190_30871# 0.061913f
C11481 a_14537_43396# a_14955_43396# 0.027267f
C11482 a_21496_47436# SINGLE_ENDED 0.055146f
C11483 a_12465_44636# VDD 0.773277f
C11484 a_n2442_46660# a_n4318_40392# 0.023735f
C11485 a_n1920_47178# a_n1605_47204# 0.08571f
C11486 a_n2109_47186# a_n815_47178# 0.160027f
C11487 a_n2497_47436# a_n971_45724# 0.229429f
C11488 a_n1741_47186# SMPL_ON_P 0.178214f
C11489 a_13887_32519# VDD 0.424391f
C11490 a_n784_42308# a_961_42354# 0.038477f
C11491 a_5342_30871# VDAC_N 0.011631f
C11492 a_11967_42832# a_12281_43396# 0.027232f
C11493 a_3499_42826# a_n97_42460# 0.019497f
C11494 a_20528_46660# VDD 0.077608f
C11495 a_2324_44458# a_11827_44484# 0.03555f
C11496 a_5937_45572# a_n2661_44458# 0.061693f
C11497 a_19692_46634# a_17517_44484# 0.023737f
C11498 a_13259_45724# a_14180_45002# 0.04353f
C11499 a_2957_45546# a_413_45260# 0.012841f
C11500 a_n357_42282# a_2382_45260# 0.025504f
C11501 a_13904_45546# a_14033_45572# 0.010132f
C11502 a_4185_45028# a_n699_43396# 0.027874f
C11503 a_3483_46348# a_5343_44458# 0.046505f
C11504 a_n443_42852# a_n913_45002# 0.796158f
C11505 a_4646_46812# a_7542_44172# 0.012612f
C11506 a_13747_46662# a_15493_43940# 0.049242f
C11507 a_12549_44172# a_14021_43940# 0.150377f
C11508 a_n237_47217# a_6755_46942# 0.073038f
C11509 a_n2312_39304# a_n2840_46634# 0.018018f
C11510 a_n2312_40392# a_n2956_39768# 0.056063f
C11511 a_21613_42308# a_22485_38105# 0.026117f
C11512 a_5837_42852# VDD 0.1774f
C11513 a_20974_43370# a_21487_43396# 0.03755f
C11514 a_2711_45572# VDD 1.22011f
C11515 a_526_44458# a_2675_43914# 0.03283f
C11516 a_10903_43370# a_10807_43548# 0.193971f
C11517 a_n1613_43370# a_8605_42826# 0.159791f
C11518 a_n913_45002# a_375_42282# 0.01541f
C11519 a_4185_45028# a_22959_43948# 0.014665f
C11520 a_n2956_38680# a_n4318_39768# 0.023254f
C11521 a_n2956_39304# a_n3674_39768# 0.02324f
C11522 a_11599_46634# a_19553_46090# 0.021903f
C11523 a_6755_46942# a_8270_45546# 0.045608f
C11524 a_10428_46928# a_11186_47026# 0.055625f
C11525 a_n881_46662# a_167_45260# 0.108232f
C11526 a_16327_47482# a_17715_44484# 0.03083f
C11527 a_13747_46662# a_12741_44636# 0.099721f
C11528 a_4791_45118# a_526_44458# 0.042209f
C11529 a_n443_46116# a_2981_46116# 0.017561f
C11530 a_n1435_47204# a_6945_45028# 0.030745f
C11531 a_4883_46098# a_9290_44172# 0.055265f
C11532 a_10227_46804# a_15015_46420# 0.287571f
C11533 a_n237_47217# a_8049_45260# 0.109887f
C11534 a_n4209_39304# VIN_P 0.049227f
C11535 a_14209_32519# a_5342_30871# 0.028644f
C11536 a_n97_42460# a_133_42852# 0.012177f
C11537 a_n863_45724# a_1568_43370# 0.202455f
C11538 a_n2661_45546# a_3080_42308# 0.155045f
C11539 a_1138_42852# a_791_42968# 0.100783f
C11540 a_11691_44458# a_n2661_44458# 0.021716f
C11541 a_1423_45028# a_9313_44734# 0.241551f
C11542 a_n2312_40392# a_n4318_37592# 0.025292f
C11543 a_16327_47482# a_15861_45028# 0.030602f
C11544 a_8270_45546# a_8049_45260# 0.321896f
C11545 a_376_46348# a_472_46348# 0.318161f
C11546 a_n2497_47436# a_n2293_45010# 0.233882f
C11547 a_16388_46812# a_17957_46116# 0.140894f
C11548 a_10796_42968# a_11136_42852# 0.027606f
C11549 a_2982_43646# a_7174_31319# 0.081795f
C11550 a_n4318_39304# a_n4334_39392# 0.081919f
C11551 a_22485_44484# VDD 0.258874f
C11552 a_11827_44484# a_19862_44208# 0.015537f
C11553 a_7499_43078# a_7871_42858# 0.146369f
C11554 a_18184_42460# a_11341_43940# 0.029749f
C11555 a_n452_47436# VDD 0.092189f
C11556 a_n2109_47186# DATA[1] 0.049689f
C11557 a_n2956_38680# a_n2956_38216# 0.10753f
C11558 a_5937_45572# a_5907_45546# 0.104991f
C11559 a_4646_46812# a_5205_44484# 0.094488f
C11560 a_11453_44696# a_11691_44458# 0.035893f
C11561 a_4190_30871# VDAC_P 0.044618f
C11562 a_10554_47026# CLK 0.014924f
C11563 a_5891_43370# a_8685_43396# 0.145735f
C11564 a_3422_30871# a_14401_32519# 0.096501f
C11565 a_13249_42308# a_13291_42460# 0.068754f
C11566 a_n2956_39304# a_n4315_30879# 0.024812f
C11567 a_n443_42852# a_1755_42282# 0.055323f
C11568 a_2675_43914# a_3353_43940# 0.011812f
C11569 a_2324_44458# a_15595_45028# 0.04743f
C11570 a_8746_45002# a_10490_45724# 0.116339f
C11571 a_526_44458# a_3429_45260# 0.010386f
C11572 a_n1925_42282# a_3065_45002# 0.04956f
C11573 a_768_44030# a_5244_44056# 0.167173f
C11574 a_10193_42453# a_11322_45546# 0.024616f
C11575 a_3483_46348# a_8560_45348# 0.021507f
C11576 a_15227_44166# a_14539_43914# 0.520312f
C11577 a_12741_44636# a_18911_45144# 0.013476f
C11578 a_n746_45260# a_n2293_46634# 0.048005f
C11579 a_6151_47436# a_768_44030# 0.096889f
C11580 a_11459_47204# a_n881_46662# 0.0707f
C11581 a_18479_47436# a_11453_44696# 0.018416f
C11582 a_14113_42308# a_16522_42674# 0.183181f
C11583 a_1823_45246# a_3600_43914# 0.016141f
C11584 a_n443_42852# a_n2661_44458# 0.045408f
C11585 a_17339_46660# a_15493_43396# 0.075223f
C11586 a_n357_42282# a_5343_44458# 0.022768f
C11587 a_13059_46348# a_11341_43940# 0.025185f
C11588 a_12549_44172# a_19692_46634# 0.491923f
C11589 a_n443_46116# a_167_45260# 0.794635f
C11590 a_3877_44458# a_5167_46660# 0.032716f
C11591 a_4646_46812# a_5385_46902# 0.042888f
C11592 a_4651_46660# a_4817_46660# 0.57393f
C11593 a_11599_46634# a_12741_44636# 0.183316f
C11594 a_11453_44696# a_17829_46910# 0.013408f
C11595 a_n237_47217# a_8953_45546# 0.090521f
C11596 a_2063_45854# a_5204_45822# 0.174206f
C11597 a_13747_46662# a_13607_46688# 0.168294f
C11598 a_n3565_38502# a_n3565_37414# 0.030671f
C11599 a_n4209_38502# a_n3420_37440# 0.033073f
C11600 a_n3420_38528# a_n4209_37414# 0.027951f
C11601 a_n2293_43922# a_5742_30871# 0.098838f
C11602 a_n356_44636# a_17531_42308# 0.030778f
C11603 a_n2472_45002# VDD 0.217954f
C11604 a_2437_43646# CLK 0.101524f
C11605 a_4361_42308# a_13678_32519# 0.048617f
C11606 a_13467_32519# a_5649_42852# 0.042596f
C11607 a_3357_43084# DATA[4] 0.035981f
C11608 a_375_42282# a_n2661_44458# 0.025194f
C11609 a_526_44458# a_1209_43370# 0.057216f
C11610 a_9290_44172# a_8685_43396# 0.207262f
C11611 a_20273_46660# a_21188_46660# 0.118759f
C11612 a_20107_46660# a_20528_46660# 0.083408f
C11613 a_4915_47217# a_11823_42460# 0.016758f
C11614 a_13747_46662# a_16375_45002# 0.021583f
C11615 a_8270_45546# a_8953_45546# 1.06716f
C11616 a_n881_46662# a_n863_45724# 0.023273f
C11617 a_3090_45724# a_3483_46348# 0.060766f
C11618 C3_N_btm VREF_GND 0.67174f
C11619 C2_N_btm VCM 0.716172f
C11620 C4_N_btm VREF 0.98728f
C11621 C5_N_btm VIN_N 0.502041f
C11622 VDD DATA[2] 0.3216f
C11623 a_2982_43646# a_5932_42308# 0.073161f
C11624 a_n97_42460# a_5742_30871# 0.259664f
C11625 a_16137_43396# a_16877_42852# 0.010276f
C11626 a_19963_31679# a_14401_32519# 0.053905f
C11627 a_n356_44636# a_n2661_42834# 0.024765f
C11628 w_10694_33990# VDAC_N 0.143015f
C11629 a_n1853_46287# a_n1079_45724# 0.02186f
C11630 a_768_44030# a_5111_44636# 0.154519f
C11631 a_n2293_46634# a_n2109_45247# 0.016559f
C11632 a_2107_46812# a_2437_43646# 0.185914f
C11633 a_3080_42308# EN_VIN_BSTR_N 0.04304f
C11634 a_n3674_39304# a_n3420_39616# 0.152699f
C11635 a_14401_32519# VDD 0.562852f
C11636 a_3537_45260# a_8037_42858# 0.010068f
C11637 a_n913_45002# a_14543_43071# 0.036401f
C11638 a_n1059_45260# a_5534_30871# 0.025423f
C11639 a_18184_42460# a_10341_43396# 0.034231f
C11640 a_18579_44172# a_15493_43396# 0.070538f
C11641 a_5663_43940# a_6453_43914# 0.017005f
C11642 a_33_46660# VDD 0.272723f
C11643 a_21588_30879# VREF_GND 0.083908f
C11644 a_n2661_46634# CLK 0.032279f
C11645 a_22612_30879# VREF 1.73216f
C11646 a_8199_44636# a_n913_45002# 0.018004f
C11647 a_8953_45546# a_n2017_45002# 0.080521f
C11648 a_13661_43548# a_13857_44734# 0.012574f
C11649 a_11415_45002# a_13777_45326# 0.021087f
C11650 a_6851_47204# a_7227_47204# 0.241208f
C11651 a_6545_47178# a_6575_47204# 0.11927f
C11652 a_4915_47217# a_9313_45822# 0.366722f
C11653 a_n2109_47186# a_4883_46098# 0.029241f
C11654 a_18817_42826# VDD 0.204624f
C11655 a_6123_31319# a_5934_30871# 15.8951f
C11656 a_10807_43548# a_8685_43396# 0.029811f
C11657 a_12005_46116# VDD 0.518463f
C11658 a_9313_44734# a_15567_42826# 0.01457f
C11659 a_n2956_37592# a_n3674_38216# 0.023192f
C11660 a_8199_44636# CLK 0.231904f
C11661 a_n2017_45002# a_n961_42308# 0.012655f
C11662 a_18175_45572# a_19256_45572# 0.102355f
C11663 a_18341_45572# a_18691_45572# 0.206455f
C11664 a_3483_46348# a_14815_43914# 0.036548f
C11665 a_8746_45002# a_6171_45002# 0.069475f
C11666 a_20202_43084# a_20679_44626# 0.035147f
C11667 a_8270_45546# a_9028_43914# 0.233359f
C11668 a_n1613_43370# a_5275_47026# 0.039193f
C11669 a_n743_46660# a_n2438_43548# 0.426835f
C11670 a_n1925_46634# a_171_46873# 0.027689f
C11671 a_n4334_39392# a_n4334_38528# 0.050585f
C11672 a_n4209_39304# a_n3565_38502# 0.029672f
C11673 a_n3565_39304# a_n4209_38502# 5.79402f
C11674 a_n2946_39072# a_n2860_39072# 0.011479f
C11675 a_1184_42692# VDD 0.813074f
C11676 a_5934_30871# EN_VIN_BSTR_P 0.074693f
C11677 a_16243_43396# a_16547_43609# 0.165289f
C11678 a_16137_43396# a_16409_43396# 0.011989f
C11679 a_n2661_42834# a_n3674_38680# 0.03399f
C11680 a_18494_42460# a_18057_42282# 0.085802f
C11681 a_18184_42460# a_18727_42674# 0.044914f
C11682 a_n2810_45028# a_n4209_37414# 0.09606f
C11683 a_14033_45822# VDD 0.195067f
C11684 a_15227_44166# a_17324_43396# 0.010717f
C11685 a_n357_42282# a_453_43940# 0.027908f
C11686 a_13059_46348# a_10341_43396# 0.014853f
C11687 a_n755_45592# a_1414_42308# 0.013035f
C11688 a_2437_43646# a_n2661_44458# 0.036499f
C11689 a_n237_47217# a_1609_45822# 0.141985f
C11690 a_2905_45572# a_2957_45546# 0.137248f
C11691 a_n443_46116# a_n863_45724# 0.055503f
C11692 a_13747_46662# a_18985_46122# 0.035795f
C11693 a_2107_46812# a_8199_44636# 0.022874f
C11694 a_11599_46634# a_16375_45002# 0.407484f
C11695 VDAC_N C9_N_btm 0.44188p
C11696 a_4338_37500# RST_Z 0.01719f
C11697 a_5088_37509# VDD 1.15925f
C11698 a_17595_43084# a_17333_42852# 0.057438f
C11699 a_n443_42852# a_9145_43396# 2.32123f
C11700 a_5111_44636# a_7845_44172# 0.063408f
C11701 en_comp a_n2661_42282# 0.103098f
C11702 a_11453_44696# a_2437_43646# 0.189184f
C11703 a_n746_45260# a_626_44172# 0.011647f
C11704 a_11189_46129# a_11133_46155# 0.203074f
C11705 a_16388_46812# a_13259_45724# 0.030634f
C11706 a_5534_30871# a_1606_42308# 0.030581f
C11707 a_15682_43940# VDD 1.22657f
C11708 a_14537_43396# a_15095_43370# 0.019641f
C11709 a_20447_31679# a_13678_32519# 0.051589f
C11710 a_19479_31679# a_14209_32519# 0.051176f
C11711 a_4223_44672# a_5829_43940# 0.037008f
C11712 a_3422_30871# a_20512_43084# 0.125955f
C11713 a_n1059_45260# a_4190_30871# 0.133926f
C11714 a_13507_46334# SINGLE_ENDED 0.111959f
C11715 a_21811_47423# VDD 0.201359f
C11716 w_10694_33990# a_17730_32519# 0.03159f
C11717 a_10809_44734# a_11823_42460# 0.215753f
C11718 a_2324_44458# a_10907_45822# 0.025622f
C11719 a_n2109_47186# a_n1605_47204# 0.041602f
C11720 a_22223_43396# VDD 0.279195f
C11721 a_n784_42308# a_1184_42692# 0.026118f
C11722 a_564_42282# a_n1794_35082# 0.156633f
C11723 a_17364_32525# C7_N_btm 0.072179f
C11724 a_765_45546# CLK 0.0309f
C11725 a_22000_46634# VDD 0.257047f
C11726 a_8199_44636# a_n2661_44458# 0.069807f
C11727 a_n443_42852# a_n1059_45260# 0.130036f
C11728 a_4185_45028# a_4223_44672# 0.031094f
C11729 a_4646_46812# a_7281_43914# 0.021965f
C11730 a_13661_43548# a_15493_43940# 1.28948f
C11731 a_13259_45724# a_13777_45326# 0.043567f
C11732 a_4883_46098# a_n1925_46634# 0.030451f
C11733 a_13507_46334# a_n743_46660# 0.024694f
C11734 a_n971_45724# a_6969_46634# 0.235123f
C11735 a_11453_44696# a_n2661_46634# 0.032889f
C11736 a_n1151_42308# a_5257_43370# 0.058425f
C11737 a_5193_42852# VDD 0.187605f
C11738 a_20974_43370# a_20556_43646# 0.076332f
C11739 a_526_44458# a_895_43940# 0.018069f
C11740 a_10903_43370# a_10949_43914# 0.451961f
C11741 a_n1613_43370# a_8037_42858# 0.047354f
C11742 a_n1059_45260# a_375_42282# 0.0165f
C11743 a_4185_45028# a_15493_43940# 0.039364f
C11744 a_3232_43370# a_6171_45002# 0.314056f
C11745 a_n2956_39304# a_n4318_39768# 0.023377f
C11746 a_11599_46634# a_18985_46122# 0.570252f
C11747 a_10428_46928# a_10768_47026# 0.027606f
C11748 a_13661_43548# a_12741_44636# 0.13948f
C11749 a_n881_46662# a_2202_46116# 0.051959f
C11750 a_4883_46098# a_10355_46116# 0.23167f
C11751 a_10227_46804# a_14275_46494# 0.18614f
C11752 a_19321_45002# a_11415_45002# 0.065361f
C11753 a_n4209_38216# C3_P_btm 0.041776f
C11754 comp_n VDD 0.504807f
C11755 a_n2661_45546# a_4699_43561# 0.013733f
C11756 a_19479_31679# a_17730_32519# 0.052745f
C11757 a_n2312_39304# a_n3674_38216# 0.023615f
C11758 a_3877_44458# a_n2661_45546# 0.026409f
C11759 a_n881_46662# a_11823_42460# 0.036994f
C11760 a_n971_45724# a_3357_43084# 0.565799f
C11761 a_16327_47482# a_8696_44636# 0.087584f
C11762 a_n2293_46098# a_167_45260# 0.086636f
C11763 a_n2157_42858# a_n2104_42282# 0.011248f
C11764 a_17730_32519# C9_N_btm 0.215899f
C11765 a_4190_30871# a_1606_42308# 0.018892f
C11766 a_n4318_39304# a_n4209_39304# 0.135369f
C11767 a_20512_43084# VDD 0.317257f
C11768 a_n815_47178# VDD 0.380339f
C11769 a_3065_45002# a_3539_42460# 0.300764f
C11770 a_7499_43078# a_7227_42852# 0.126148f
C11771 a_n2109_47186# DATA[0] 0.08202f
C11772 a_21076_30879# a_14097_32519# 0.054945f
C11773 a_n2956_39304# a_n2956_38216# 0.05012f
C11774 a_584_46384# a_n356_44636# 0.268036f
C11775 a_19466_46812# a_19256_45572# 0.041135f
C11776 a_10623_46897# CLK 0.016177f
C11777 a_2324_44458# a_15415_45028# 0.03757f
C11778 a_10193_42453# a_10490_45724# 0.062365f
C11779 a_526_44458# a_3065_45002# 0.138202f
C11780 a_n443_46116# a_2455_43940# 0.010179f
C11781 a_20202_43084# a_18494_42460# 0.166633f
C11782 a_768_44030# a_3905_42865# 0.011432f
C11783 a_4185_45028# a_n2293_42834# 0.022725f
C11784 a_1823_45246# a_n2661_43370# 0.112095f
C11785 w_10694_33990# a_17538_32519# 0.039343f
C11786 a_15227_44166# a_16112_44458# 0.073746f
C11787 a_n971_45724# a_n2293_46634# 0.090091f
C11788 a_n1151_42308# a_5807_45002# 1.52318f
C11789 a_6151_47436# a_12549_44172# 0.214024f
C11790 a_6575_47204# a_8128_46384# 0.105633f
C11791 a_9313_45822# a_n881_46662# 1.00227f
C11792 a_n1741_47186# a_n743_46660# 0.017496f
C11793 a_21177_47436# a_13507_46334# 0.329096f
C11794 a_n3674_38216# a_n3420_38528# 0.152701f
C11795 a_n4318_38216# a_n4064_38528# 0.057645f
C11796 a_n97_42460# a_6293_42852# 0.018467f
C11797 a_14021_43940# a_16409_43396# 0.025204f
C11798 a_1823_45246# a_2998_44172# 0.062531f
C11799 a_8696_44636# a_14537_43396# 0.024289f
C11800 a_13507_46334# a_4361_42308# 0.040714f
C11801 a_n755_45592# a_n699_43396# 0.185444f
C11802 a_11453_44696# a_765_45546# 0.010973f
C11803 a_3877_44458# a_5385_46902# 0.021989f
C11804 a_4646_46812# a_4817_46660# 0.588038f
C11805 a_4651_46660# a_4955_46873# 0.140348f
C11806 a_4883_46098# a_20411_46873# 0.012008f
C11807 a_n237_47217# a_5937_45572# 0.08715f
C11808 a_2063_45854# a_5164_46348# 0.022664f
C11809 a_2113_38308# VDAC_Pi 0.170941f
C11810 a_4361_42308# a_21855_43396# 0.167446f
C11811 a_13467_32519# a_13678_32519# 10.9526f
C11812 a_n356_44636# a_17303_42282# 0.10316f
C11813 a_n2661_45010# VDD 0.842431f
C11814 a_3357_43084# DATA[3] 0.066637f
C11815 a_6171_45002# a_8975_43940# 0.175346f
C11816 a_526_44458# a_458_43396# 0.085782f
C11817 a_8199_44636# a_9145_43396# 0.020485f
C11818 SMPL_ON_P a_n3674_37592# 0.051734f
C11819 a_n971_45724# a_n473_42460# 0.094491f
C11820 a_13059_46348# a_11415_45002# 0.225168f
C11821 a_20841_46902# a_20623_46660# 0.209641f
C11822 a_20273_46660# a_21363_46634# 0.042415f
C11823 a_n743_46660# a_10586_45546# 0.018104f
C11824 a_8270_45546# a_5937_45572# 0.29626f
C11825 a_n1613_43370# a_n863_45724# 0.027265f
C11826 a_765_45546# a_17639_46660# 0.094916f
C11827 a_3090_45724# a_3147_46376# 0.010392f
C11828 C2_N_btm VREF_GND 0.671742f
C11829 C1_N_btm VCM 0.716121f
C11830 C3_N_btm VREF 0.984942f
C11831 C4_N_btm VIN_N 0.50261f
C11832 VDD DATA[1] 0.321585f
C11833 a_16137_43396# a_16245_42852# 0.016079f
C11834 a_3080_42308# a_5934_30871# 1.27306f
C11835 a_n2661_43370# a_n3674_39768# 0.144159f
C11836 a_9482_43914# a_11341_43940# 0.037822f
C11837 a_19479_31679# a_17538_32519# 0.051112f
C11838 a_768_44030# a_5147_45002# 0.191082f
C11839 a_11189_46129# a_10586_45546# 0.028266f
C11840 a_3090_45724# a_13249_42308# 0.032019f
C11841 a_n2293_46634# a_n2293_45010# 0.036081f
C11842 a_21381_43940# VDD 0.344882f
C11843 a_5111_44636# a_5111_42852# 0.148196f
C11844 a_n913_45002# a_13460_43230# 0.04239f
C11845 a_n2017_45002# a_5534_30871# 0.025363f
C11846 a_11967_42832# a_15493_43940# 0.299734f
C11847 a_19279_43940# a_19862_44208# 0.012567f
C11848 a_18579_44172# a_19328_44172# 0.053539f
C11849 a_1115_44172# a_1241_44260# 0.013015f
C11850 a_171_46873# VDD 0.539781f
C11851 a_22612_30879# VIN_N 0.18996f
C11852 a_21588_30879# VREF 0.860047f
C11853 a_5257_43370# a_4223_44672# 0.016657f
C11854 a_8199_44636# a_n1059_45260# 0.019728f
C11855 a_3503_45724# a_3775_45552# 0.13675f
C11856 a_4185_45028# a_413_45260# 0.191095f
C11857 a_n2293_46634# a_9313_44734# 0.022598f
C11858 a_11415_45002# a_13556_45296# 0.16025f
C11859 a_6151_47436# a_6575_47204# 0.047329f
C11860 a_4915_47217# a_11031_47542# 0.125943f
C11861 a_6123_31319# a_7963_42308# 0.192155f
C11862 a_18249_42858# VDD 0.250132f
C11863 a_10903_43370# VDD 2.60588f
C11864 a_9313_44734# a_5342_30871# 0.026413f
C11865 a_n2017_45002# a_n1329_42308# 0.018315f
C11866 a_3422_30871# a_5649_42852# 0.291966f
C11867 a_n2810_45028# a_n3674_38216# 0.023217f
C11868 en_comp a_n4318_38216# 0.064646f
C11869 a_19319_43548# a_19741_43940# 0.048788f
C11870 a_n2956_39768# a_n4318_39304# 0.02353f
C11871 a_18341_45572# a_18909_45814# 0.170692f
C11872 a_18479_45785# a_18691_45572# 0.036486f
C11873 a_18175_45572# a_19431_45546# 0.043567f
C11874 a_10193_42453# a_6171_45002# 0.411891f
C11875 a_8746_45002# a_3232_43370# 0.439467f
C11876 a_n2293_45546# a_n2661_43370# 0.131199f
C11877 a_20202_43084# a_20640_44752# 0.027593f
C11878 a_n1613_43370# a_5072_46660# 0.012366f
C11879 a_n1925_46634# a_n133_46660# 0.053144f
C11880 a_n1021_46688# a_n2438_43548# 0.053225f
C11881 a_12861_44030# a_3090_45724# 0.496275f
C11882 a_n4209_39590# a_n3565_38216# 0.03183f
C11883 a_n4064_40160# a_n4064_37984# 0.067467f
C11884 a_1576_42282# VDD 0.26017f
C11885 a_n3565_39590# a_n4209_38216# 0.0313f
C11886 a_16137_43396# a_16547_43609# 0.151161f
C11887 a_3080_42308# a_3935_42891# 0.017131f
C11888 a_18184_42460# a_18057_42282# 0.19301f
C11889 a_15227_44166# a_17499_43370# 0.021724f
C11890 a_6709_45028# a_n2661_43370# 0.041021f
C11891 a_19479_31679# a_19721_31679# 9.039419f
C11892 a_n357_42282# a_1414_42308# 0.027118f
C11893 a_n743_46660# a_11189_46129# 0.039903f
C11894 a_13747_46662# a_18819_46122# 0.039742f
C11895 a_n1151_42308# a_n755_45592# 0.03818f
C11896 a_4338_37500# VDD 0.525635f
C11897 EN_VIN_BSTR_P a_n217_35014# 0.651142f
C11898 VDAC_N C8_N_btm 0.220913p
C11899 a_3726_37500# RST_Z 1.60318f
C11900 a_n4209_37414# VIN_P 0.028788f
C11901 a_n4318_39304# a_n4318_37592# 0.023243f
C11902 a_18114_32519# C10_N_btm 0.460005f
C11903 a_16795_42852# a_17333_42852# 0.108694f
C11904 a_17595_43084# a_18083_42858# 0.046381f
C11905 a_3232_43370# a_5663_43940# 0.090892f
C11906 a_n357_42282# a_12281_43396# 0.022975f
C11907 a_5111_44636# a_7542_44172# 0.039468f
C11908 a_13059_46348# a_13259_45724# 0.812126f
C11909 a_12465_44636# a_3357_43084# 1.30897f
C11910 a_9290_44172# a_11133_46155# 0.051331f
C11911 a_n1641_46494# a_n1533_46116# 0.057222f
C11912 a_10227_46804# a_n913_45002# 0.344574f
C11913 a_8270_45546# a_n443_42852# 0.063811f
C11914 a_13747_46662# a_16223_45938# 0.02646f
C11915 a_6151_47436# a_5205_44484# 0.010575f
C11916 a_14955_43940# VDD 0.253201f
C11917 a_14537_43396# a_14205_43396# 0.080783f
C11918 a_21177_47436# SINGLE_ENDED 0.057266f
C11919 a_10227_46804# CLK 0.207445f
C11920 a_4883_46098# VDD 1.12729f
C11921 a_4223_44672# a_5745_43940# 0.040431f
C11922 a_4185_45028# a_5379_42460# 0.189676f
C11923 a_18989_43940# a_15493_43940# 0.025737f
C11924 a_n2017_45002# a_4190_30871# 0.025499f
C11925 a_12741_44636# a_20273_45572# 0.028616f
C11926 a_18597_46090# a_9313_44734# 0.029282f
C11927 a_11189_46129# a_11136_45572# 0.042798f
C11928 a_20202_43084# a_21188_45572# 0.013137f
C11929 a_11415_45002# a_21363_45546# 0.011178f
C11930 a_10809_44734# a_12427_45724# 0.01284f
C11931 a_5649_42852# VDD 0.438443f
C11932 a_13678_32519# RST_Z 0.048939f
C11933 a_n1920_47178# a_n1741_47186# 0.173125f
C11934 a_n2109_47186# SMPL_ON_P 0.049302f
C11935 COMP_P a_1606_42308# 2.67743f
C11936 a_n784_42308# a_1576_42282# 0.038241f
C11937 a_n3674_37592# a_n1794_35082# 0.096752f
C11938 a_9313_44734# a_743_42282# 0.024013f
C11939 a_21188_46660# VDD 0.284105f
C11940 a_18597_46090# a_20974_43370# 0.025672f
C11941 a_n443_42852# a_n2017_45002# 0.033337f
C11942 a_n443_46116# a_2982_43646# 0.140614f
C11943 a_13259_45724# a_13556_45296# 0.019616f
C11944 a_2711_45572# a_3357_43084# 0.037825f
C11945 a_12465_44636# a_n2293_46634# 0.012816f
C11946 a_n971_45724# a_6755_46942# 0.185154f
C11947 a_7227_47204# a_4646_46812# 0.01221f
C11948 a_4649_42852# VDD 0.194775f
C11949 a_526_44458# a_2479_44172# 0.08343f
C11950 a_10903_43370# a_10729_43914# 0.082892f
C11951 a_n1613_43370# a_7765_42852# 0.081834f
C11952 a_n2293_45010# a_626_44172# 0.024201f
C11953 a_n2017_45002# a_375_42282# 0.03181f
C11954 a_5111_44636# a_5205_44484# 0.200189f
C11955 a_5691_45260# a_6171_45002# 0.057463f
C11956 a_n913_45002# a_1307_43914# 0.298747f
C11957 a_9290_44172# a_12429_44172# 0.040422f
C11958 a_8746_45002# a_8975_43940# 0.016889f
C11959 a_11599_46634# a_18819_46122# 0.314824f
C11960 a_2063_45854# a_5066_45546# 0.055269f
C11961 a_16327_47482# a_15682_46116# 0.050548f
C11962 a_5807_45002# a_12741_44636# 0.041091f
C11963 a_n881_46662# a_1823_45246# 0.155149f
C11964 a_11459_47204# a_6945_45028# 0.010682f
C11965 a_4883_46098# a_9823_46155# 0.046689f
C11966 a_n971_45724# a_8049_45260# 0.078318f
C11967 a_10227_46804# a_14493_46090# 0.202633f
C11968 a_8530_39574# CAL_N 0.644218f
C11969 a_1666_39043# VDD 2.8964f
C11970 a_14209_32519# a_5534_30871# 0.057361f
C11971 a_13887_32519# a_5342_30871# 0.028465f
C11972 a_9482_43914# a_n2293_43922# 0.018115f
C11973 a_n2661_45546# a_4235_43370# 0.088313f
C11974 a_n2312_40392# a_n3674_38216# 0.025514f
C11975 SMPL_ON_N COMP_P 2.13156f
C11976 a_n2497_47436# a_n2661_45010# 0.281004f
C11977 a_16327_47482# a_16680_45572# 0.223571f
C11978 a_768_44030# a_7499_43078# 0.101779f
C11979 a_n237_47217# a_2437_43646# 0.076344f
C11980 a_16388_46812# a_17715_44484# 0.032772f
C11981 a_10341_42308# a_11554_42852# 0.170124f
C11982 a_743_42282# a_961_42354# 0.016854f
C11983 a_3626_43646# a_19647_42308# 0.170024f
C11984 a_5649_42852# a_n784_42308# 0.043382f
C11985 a_n1605_47204# VDD 0.20224f
C11986 a_3065_45002# a_3626_43646# 0.480498f
C11987 a_9625_46129# a_2711_45572# 0.019316f
C11988 a_10227_46804# a_n2661_44458# 0.034728f
C11989 a_19466_46812# a_19431_45546# 0.038922f
C11990 a_4646_46812# a_6171_45002# 0.032849f
C11991 a_2107_46812# a_1307_43914# 0.015866f
C11992 a_8685_43396# VDD 0.261626f
C11993 a_4190_30871# VDAC_N 0.048476f
C11994 a_10467_46802# CLK 0.028547f
C11995 a_12741_44636# a_18315_45260# 0.011294f
C11996 a_2324_44458# a_14797_45144# 0.048583f
C11997 a_10193_42453# a_8746_45002# 0.11003f
C11998 a_526_44458# a_2680_45002# 0.119733f
C11999 a_n443_46116# a_2253_43940# 0.011444f
C12000 a_1138_42852# a_n2661_43370# 0.023497f
C12001 a_11415_45002# a_19778_44110# 0.030651f
C12002 a_20202_43084# a_18184_42460# 0.299795f
C12003 a_768_44030# a_3600_43914# 0.182408f
C12004 a_3090_45724# a_18287_44626# 0.037072f
C12005 a_n237_47217# a_n2661_46634# 0.067716f
C12006 a_6151_47436# a_12891_46348# 0.169139f
C12007 a_7903_47542# a_8128_46384# 0.109077f
C12008 a_11031_47542# a_n881_46662# 0.183988f
C12009 a_20990_47178# a_13507_46334# 0.017412f
C12010 a_10227_46804# a_11453_44696# 0.08211f
C12011 a_3905_42865# a_5111_42852# 0.079376f
C12012 a_15599_45572# a_16751_45260# 0.012353f
C12013 a_13507_46334# a_13467_32519# 0.043891f
C12014 a_17339_46660# a_18451_43940# 0.012866f
C12015 a_n357_42282# a_n699_43396# 0.055761f
C12016 a_3160_47472# a_3699_46348# 0.109505f
C12017 a_11453_44696# a_17339_46660# 0.071641f
C12018 a_3877_44458# a_4817_46660# 0.017126f
C12019 a_4646_46812# a_4955_46873# 0.047208f
C12020 a_n443_46116# a_1823_45246# 0.217935f
C12021 a_13507_46334# a_20273_46660# 0.026778f
C12022 a_n237_47217# a_8199_44636# 0.089777f
C12023 a_n2661_46634# a_8270_45546# 0.037557f
C12024 a_n3565_38502# a_n4209_37414# 0.029366f
C12025 a_n4209_38502# a_n3565_37414# 0.030019f
C12026 a_4190_30871# a_14209_32519# 0.031783f
C12027 a_2437_43646# DATA[5] 0.059749f
C12028 a_n356_44636# a_4958_30871# 0.46356f
C12029 a_n2840_45002# VDD 0.289706f
C12030 a_3232_43370# a_8975_43940# 0.620589f
C12031 a_7499_43078# a_7845_44172# 0.112307f
C12032 a_20273_46660# a_20623_46660# 0.20669f
C12033 a_20107_46660# a_21188_46660# 0.102355f
C12034 a_n1613_43370# a_n1079_45724# 0.013012f
C12035 a_5807_45002# a_16375_45002# 0.042941f
C12036 a_8270_45546# a_8199_44636# 0.95539f
C12037 a_17339_46660# a_17639_46660# 0.081726f
C12038 C1_N_btm VREF_GND 0.673422f
C12039 C0_N_btm VCM 0.717064f
C12040 C2_N_btm VREF 0.987884f
C12041 C3_N_btm VIN_N 0.455045f
C12042 VDD DATA[0] 1.05526f
C12043 a_n2661_43370# a_n4318_39768# 0.068386f
C12044 a_2711_45572# a_743_42282# 0.039036f
C12045 a_2382_45260# a_3737_43940# 0.027805f
C12046 a_8270_45546# a_8192_45572# 0.048422f
C12047 a_11453_44696# a_1307_43914# 0.037741f
C12048 a_4883_46098# a_1423_45028# 0.022493f
C12049 a_9290_44172# a_10586_45546# 0.264957f
C12050 a_n881_46662# a_6709_45028# 0.011804f
C12051 a_12594_46348# a_8049_45260# 0.069217f
C12052 a_19741_43940# VDD 0.153579f
C12053 a_18599_43230# a_18695_43230# 0.013793f
C12054 a_17538_32519# C8_N_btm 0.090298f
C12055 a_5495_43940# a_5663_43940# 0.227135f
C12056 a_n913_45002# a_13635_43156# 0.036742f
C12057 a_18579_44172# a_18451_43940# 0.147572f
C12058 a_19279_43940# a_19478_44306# 0.03583f
C12059 a_21588_30879# VIN_N 0.106569f
C12060 a_n133_46660# VDD 0.483405f
C12061 a_8199_44636# a_n2017_45002# 0.020035f
C12062 a_584_46384# a_3499_42826# 0.036739f
C12063 a_2277_45546# a_2711_45572# 0.01233f
C12064 a_1823_45246# a_3537_45260# 0.482502f
C12065 a_11415_45002# a_9482_43914# 0.309633f
C12066 a_6491_46660# a_6851_47204# 0.132946f
C12067 a_4915_47217# a_9863_47436# 0.018512f
C12068 a_17333_42852# VDD 0.525529f
C12069 a_3422_30871# a_13678_32519# 0.452533f
C12070 a_11387_46155# VDD 0.099732f
C12071 en_comp a_n2472_42282# 0.018838f
C12072 a_n2293_42834# a_n2293_42282# 0.018879f
C12073 a_n2017_45002# COMP_P 0.012669f
C12074 a_n2956_37592# a_n4318_38216# 0.023067f
C12075 a_768_44030# a_1756_43548# 0.093469f
C12076 a_18175_45572# a_18691_45572# 0.105995f
C12077 a_18479_45785# a_18909_45814# 0.023226f
C12078 a_n755_45592# a_n2293_42834# 0.059468f
C12079 a_10193_42453# a_3232_43370# 0.016241f
C12080 a_10180_45724# a_6171_45002# 0.03378f
C12081 a_n2956_38216# a_n2661_43370# 0.028301f
C12082 a_10227_46804# a_9145_43396# 0.066362f
C12083 a_n1613_43370# a_6540_46812# 0.05541f
C12084 a_n2661_46634# a_1123_46634# 0.012266f
C12085 a_n1151_42308# a_14513_46634# 0.042579f
C12086 a_12465_44636# a_6755_46942# 0.021176f
C12087 a_n1021_46688# a_n743_46660# 0.11001f
C12088 a_n1925_46634# a_n2438_43548# 0.166008f
C12089 a_13487_47204# a_14084_46812# 0.012167f
C12090 a_12861_44030# a_15009_46634# 0.058082f
C12091 a_n237_47217# a_765_45546# 0.1364f
C12092 a_6123_31319# EN_VIN_BSTR_P 0.051746f
C12093 a_1067_42314# VDD 0.128996f
C12094 a_n4209_39304# a_n4209_38502# 0.042459f
C12095 a_14401_32519# a_5342_30871# 0.062032f
C12096 a_16137_43396# a_16243_43396# 0.182209f
C12097 a_7229_43940# a_n2661_43370# 0.040132f
C12098 a_19479_31679# a_18114_32519# 0.182316f
C12099 a_n863_45724# a_895_43940# 0.015488f
C12100 a_15009_46634# a_14180_46812# 0.123843f
C12101 a_n746_45260# a_n443_42852# 0.136813f
C12102 a_n743_46660# a_9290_44172# 0.048675f
C12103 a_5807_45002# a_18985_46122# 0.017912f
C12104 a_13661_43548# a_18819_46122# 0.02447f
C12105 a_2959_46660# a_3147_46376# 0.010696f
C12106 a_2107_46812# a_8016_46348# 0.022583f
C12107 a_10227_46804# a_14180_46482# 0.014179f
C12108 a_12465_44636# a_8049_45260# 0.027831f
C12109 a_3726_37500# VDD 0.341303f
C12110 a_n1057_35014# a_n217_35014# 0.481434f
C12111 VDAC_N C7_N_btm 0.11042p
C12112 a_17595_43084# a_17701_42308# 0.141211f
C12113 a_3232_43370# a_5495_43940# 0.060353f
C12114 a_20193_45348# a_9313_44734# 0.056112f
C12115 a_n746_45260# a_375_42282# 0.41439f
C12116 a_n1423_46090# a_n1533_46116# 0.097745f
C12117 a_9290_44172# a_11189_46129# 0.199578f
C12118 a_6755_46942# a_2711_45572# 0.612305f
C12119 a_10227_46804# a_n1059_45260# 0.036978f
C12120 a_13747_46662# a_16020_45572# 0.016423f
C12121 a_5755_42852# a_5932_42308# 0.012644f
C12122 a_13483_43940# VDD 0.219591f
C12123 a_14537_43396# a_14358_43442# 0.1418f
C12124 a_20990_47178# SINGLE_ENDED 0.067698f
C12125 a_19479_31679# a_13887_32519# 0.051118f
C12126 a_21496_47436# VDD 0.198362f
C12127 a_19963_31679# a_13678_32519# 0.051335f
C12128 a_20193_45348# a_20974_43370# 0.026944f
C12129 a_12741_44636# a_20107_45572# 0.029025f
C12130 a_20202_43084# a_21363_45546# 0.029873f
C12131 a_n2956_39768# a_n4318_40392# 0.023582f
C12132 a_8049_45260# a_2711_45572# 2.31131f
C12133 a_10809_44734# a_11962_45724# 0.033571f
C12134 a_13678_32519# VDD 0.455443f
C12135 a_n2497_47436# a_n1605_47204# 0.0417f
C12136 a_n2109_47186# a_n1741_47186# 0.18579f
C12137 a_n327_42558# a_n1794_35082# 0.053474f
C12138 a_n784_42308# a_1067_42314# 0.064066f
C12139 a_5891_43370# a_4361_42308# 0.028094f
C12140 a_765_45546# DATA[5] 0.027477f
C12141 a_21363_46634# VDD 0.357368f
C12142 a_8016_46348# a_n2661_44458# 0.030129f
C12143 a_n443_46116# a_2896_43646# 0.039985f
C12144 a_19321_45002# a_20623_43914# 0.294126f
C12145 a_15227_44166# a_17517_44484# 0.104904f
C12146 a_13661_43548# a_11341_43940# 0.15891f
C12147 a_13747_46662# a_21115_43940# 0.02491f
C12148 a_13259_45724# a_9482_43914# 0.321549f
C12149 a_n755_45592# a_413_45260# 0.032345f
C12150 a_n357_42282# a_327_44734# 0.078335f
C12151 a_2063_45854# a_7577_46660# 0.032724f
C12152 a_22959_47212# a_22612_30879# 0.156518f
C12153 a_9396_43370# a_9145_43396# 0.030617f
C12154 a_n4318_40392# a_n4318_37592# 0.023213f
C12155 a_n1059_45260# a_1307_43914# 0.016622f
C12156 a_10903_43370# a_10405_44172# 0.026421f
C12157 a_n1613_43370# a_7871_42858# 0.659491f
C12158 a_3483_46348# a_15493_43940# 0.026486f
C12159 a_5691_45260# a_3232_43370# 0.123939f
C12160 a_5147_45002# a_5205_44484# 0.018671f
C12161 a_10193_42453# a_8975_43940# 0.023559f
C12162 a_11599_46634# a_17957_46116# 0.031252f
C12163 a_9313_45822# a_6945_45028# 0.035455f
C12164 a_n881_46662# a_1138_42852# 0.148785f
C12165 a_13747_46662# a_11415_45002# 0.099293f
C12166 a_1123_46634# a_765_45546# 0.025395f
C12167 a_10227_46804# a_13925_46122# 0.635045f
C12168 a_8530_39574# a_11206_38545# 0.046219f
C12169 a_1169_39043# VDD 0.505762f
C12170 a_9482_43914# a_n2661_43922# 0.036658f
C12171 a_n863_45724# a_458_43396# 0.122956f
C12172 a_9290_44172# a_4361_42308# 0.1126f
C12173 a_n2661_45546# a_4093_43548# 0.343267f
C12174 a_n2312_39304# a_n4318_38216# 0.023429f
C12175 a_3090_45724# a_n1925_42282# 0.157861f
C12176 a_16327_47482# a_16855_45546# 0.305145f
C12177 a_12741_44636# a_3483_46348# 0.023452f
C12178 a_n2293_46098# a_1823_45246# 0.107882f
C12179 a_16721_46634# a_15682_46116# 0.010175f
C12180 a_16388_46812# a_17583_46090# 0.033313f
C12181 a_3626_43646# a_19511_42282# 0.182478f
C12182 a_2982_43646# a_13258_32519# 0.086314f
C12183 a_2382_45260# a_3539_42460# 0.110439f
C12184 SMPL_ON_P VDD 0.613427f
C12185 a_8953_45546# a_2711_45572# 0.032277f
C12186 a_768_44030# a_n2661_43370# 0.024666f
C12187 a_4646_46812# a_3232_43370# 0.305673f
C12188 a_n2956_38680# a_n2810_45572# 5.73878f
C12189 a_20193_45348# a_13887_32519# 0.277027f
C12190 a_10428_46928# CLK 0.032943f
C12191 a_10949_43914# a_12429_44172# 0.156922f
C12192 a_8035_47026# VDD 0.132317f
C12193 a_n755_45592# a_5379_42460# 0.038776f
C12194 a_895_43940# a_2455_43940# 0.01899f
C12195 a_12741_44636# a_17719_45144# 0.011019f
C12196 a_2324_44458# a_14537_43396# 0.341957f
C12197 a_10053_45546# a_10490_45724# 0.084842f
C12198 a_526_44458# a_2382_45260# 0.072916f
C12199 a_10180_45724# a_8746_45002# 0.304016f
C12200 w_10694_33990# a_14401_32519# 0.024342f
C12201 a_3483_46348# a_n2293_42834# 0.033766f
C12202 a_16327_47482# a_19862_44208# 0.209324f
C12203 a_768_44030# a_2998_44172# 0.571981f
C12204 a_3090_45724# a_18248_44752# 0.027743f
C12205 a_n746_45260# a_n2661_46634# 0.037885f
C12206 a_4915_47217# a_768_44030# 0.187438f
C12207 a_6151_47436# a_11309_47204# 0.065131f
C12208 a_9863_47436# a_n881_46662# 0.164043f
C12209 a_n2109_47186# a_n743_46660# 0.029623f
C12210 SMPL_ON_P a_n2312_38680# 0.041837f
C12211 a_n1741_47186# a_n1925_46634# 0.012189f
C12212 a_20990_47178# a_21177_47436# 0.159555f
C12213 a_n4318_38216# a_n3420_38528# 0.31769f
C12214 a_n3674_38680# a_n4064_38528# 0.557806f
C12215 a_14021_43940# a_16243_43396# 0.017079f
C12216 a_15493_43396# a_16823_43084# 0.029968f
C12217 a_3905_42865# a_4520_42826# 0.054799f
C12218 a_13661_43548# a_10341_43396# 0.053085f
C12219 a_15903_45785# a_16019_45002# 0.139976f
C12220 a_11652_45724# a_n2661_43370# 0.028174f
C12221 a_12549_44172# a_15781_43660# 0.062935f
C12222 a_13507_46334# a_20411_46873# 0.035522f
C12223 a_4646_46812# a_4651_46660# 0.844575f
C12224 a_3160_47472# a_3483_46348# 0.154179f
C12225 a_3877_44458# a_4955_46873# 0.029242f
C12226 a_12549_44172# a_15227_44166# 0.354423f
C12227 a_4791_45118# a_1823_45246# 0.015359f
C12228 a_n443_46116# a_1138_42852# 0.017807f
C12229 a_n971_45724# a_5937_45572# 0.027865f
C12230 a_n237_47217# a_8349_46414# 0.047427f
C12231 a_13467_32519# a_4361_42308# 0.121732f
C12232 a_2437_43646# DATA[4] 0.060047f
C12233 a_3422_30871# a_n1794_35082# 0.828871f
C12234 a_3232_43370# a_10057_43914# 0.025371f
C12235 a_4185_45028# a_10341_43396# 0.019539f
C12236 a_7229_43940# a_5883_43914# 0.026061f
C12237 a_7499_43078# a_7542_44172# 0.069089f
C12238 a_20107_46660# a_21363_46634# 0.043567f
C12239 a_20273_46660# a_20841_46902# 0.17072f
C12240 a_n1613_43370# a_n2293_45546# 0.020156f
C12241 a_13747_46662# a_13259_45724# 0.093177f
C12242 C0_N_btm VREF_GND 0.350401f
C12243 C0_dummy_N_btm VCM 0.311452f
C12244 RST_Z SINGLE_ENDED 0.0318f
C12245 C1_N_btm VREF 0.98698f
C12246 C2_N_btm VIN_N 0.502408f
C12247 VDD CLK_DATA 0.422202f
C12248 a_3626_43646# a_4921_42308# 0.431551f
C12249 a_3080_42308# a_6123_31319# 1.45722f
C12250 a_20193_45348# a_22485_44484# 0.027057f
C12251 a_22959_45036# a_22959_44484# 0.025171f
C12252 a_19479_31679# a_14401_32519# 0.053843f
C12253 a_10193_42453# a_16137_43396# 0.329316f
C12254 a_n755_45592# a_n13_43084# 0.113444f
C12255 a_10355_46116# a_10586_45546# 0.012906f
C12256 a_n2293_46098# a_n2293_45546# 0.04779f
C12257 a_n1613_43370# a_6709_45028# 0.037165f
C12258 a_3080_42308# EN_VIN_BSTR_P 0.043709f
C12259 a_18599_43230# a_18504_43218# 0.049827f
C12260 a_5013_44260# a_5663_43940# 0.083171f
C12261 a_n913_45002# a_12895_43230# 0.029875f
C12262 a_11967_42832# a_11341_43940# 0.046075f
C12263 a_18579_44172# a_18326_43940# 0.096332f
C12264 a_n2438_43548# VDD 3.40589f
C12265 a_1823_45246# a_3429_45260# 0.047931f
C12266 a_n971_45724# a_8333_44056# 0.017284f
C12267 a_3090_45724# a_16922_45042# 0.206138f
C12268 a_13507_46334# a_3422_30871# 0.074924f
C12269 a_18597_46090# a_20512_43084# 0.023158f
C12270 a_11415_45002# a_13348_45260# 0.036052f
C12271 a_6545_47178# a_6851_47204# 0.134581f
C12272 a_4915_47217# a_9067_47204# 0.061984f
C12273 a_n1151_42308# a_12861_44030# 0.029342f
C12274 a_18083_42858# VDD 0.408512f
C12275 a_7227_42308# a_6123_31319# 0.189956f
C12276 a_20512_43084# a_743_42282# 0.082751f
C12277 a_9313_44734# a_5534_30871# 0.039673f
C12278 en_comp a_n3674_38680# 0.014975f
C12279 a_n2810_45028# a_n4318_38216# 0.023084f
C12280 a_n2956_38216# a_n2302_37984# 0.041408f
C12281 a_n2017_45002# a_n4318_37592# 0.043579f
C12282 a_11133_46155# VDD 0.176249f
C12283 a_6755_46942# a_15682_43940# 0.028635f
C12284 a_768_44030# a_1568_43370# 0.077231f
C12285 a_18175_45572# a_18909_45814# 0.053479f
C12286 a_18479_45785# a_18341_45572# 0.21997f
C12287 a_n357_42282# a_n2293_42834# 4.06139f
C12288 a_9290_44172# a_5891_43370# 0.302383f
C12289 a_4185_45028# a_n2293_43922# 0.093999f
C12290 a_16375_45002# a_17719_45144# 0.201099f
C12291 a_526_44458# a_5343_44458# 0.015378f
C12292 a_13661_43548# a_n97_42460# 0.02781f
C12293 a_n1613_43370# a_5732_46660# 0.268372f
C12294 a_n1151_42308# a_14180_46812# 0.037471f
C12295 a_n2312_38680# a_n2438_43548# 0.046935f
C12296 a_n1925_46634# a_n743_46660# 0.193773f
C12297 a_n4315_30879# a_n4064_37984# 0.034375f
C12298 a_n1794_35082# VDD 3.49323f
C12299 a_n4209_39590# a_n4209_38216# 0.031951f
C12300 a_n4064_40160# a_n3420_37984# 0.053114f
C12301 a_4235_43370# a_3935_42891# 0.082011f
C12302 a_4093_43548# a_4520_42826# 0.077799f
C12303 a_18184_42460# a_17303_42282# 0.027385f
C12304 a_n863_45724# a_2479_44172# 0.047943f
C12305 a_n357_42282# a_1115_44172# 0.011627f
C12306 a_4185_45028# a_n97_42460# 0.022167f
C12307 a_1138_42852# a_1049_43396# 0.022078f
C12308 a_14084_46812# a_14180_46812# 0.318161f
C12309 a_n971_45724# a_n443_42852# 0.329303f
C12310 a_11599_46634# a_13259_45724# 0.249721f
C12311 a_n743_46660# a_10355_46116# 0.011802f
C12312 a_n2293_46634# a_10903_43370# 0.046902f
C12313 a_5807_45002# a_18819_46122# 0.012467f
C12314 a_13747_46662# a_18189_46348# 0.022348f
C12315 a_768_44030# a_10809_44734# 0.037504f
C12316 a_2609_46660# a_3483_46348# 0.010427f
C12317 a_2905_45572# a_n755_45592# 0.168143f
C12318 a_n1696_34930# a_n217_35014# 0.559484f
C12319 a_n1057_35014# EN_VIN_BSTR_P 1.06139f
C12320 VDAC_N C6_N_btm 55.2142f
C12321 a_n4318_39304# a_n3674_38216# 0.023484f
C12322 a_3232_43370# a_5013_44260# 0.081759f
C12323 a_10227_46804# a_16104_42674# 0.012196f
C12324 a_10057_43914# a_8975_43940# 0.069663f
C12325 a_2063_45854# a_9482_43914# 0.018952f
C12326 a_4883_46098# a_3357_43084# 0.060164f
C12327 a_10227_46804# a_n2017_45002# 0.030377f
C12328 a_n1991_46122# a_n1533_46116# 0.034619f
C12329 a_13747_46662# a_17478_45572# 0.073886f
C12330 a_4791_45118# a_6709_45028# 0.017539f
C12331 a_12429_44172# VDD 0.169047f
C12332 a_14537_43396# a_14579_43548# 0.046172f
C12333 a_20447_31679# a_13467_32519# 0.051601f
C12334 a_20193_45348# a_14401_32519# 0.175398f
C12335 a_20894_47436# SINGLE_ENDED 0.044283f
C12336 a_13507_46334# VDD 1.4135f
C12337 a_8270_45546# a_1307_43914# 0.050297f
C12338 a_10809_44734# a_11652_45724# 0.073342f
C12339 a_526_44458# a_4880_45572# 0.02064f
C12340 a_768_44030# a_5883_43914# 0.087568f
C12341 a_n2109_47186# a_n1920_47178# 0.070142f
C12342 a_n2497_47436# SMPL_ON_P 0.131317f
C12343 a_21855_43396# VDD 0.289066f
C12344 a_n784_42308# a_n1794_35082# 0.063076f
C12345 a_9313_44734# a_4190_30871# 0.02726f
C12346 a_11967_42832# a_10341_43396# 0.076124f
C12347 a_20623_46660# VDD 0.194217f
C12348 a_n357_42282# a_413_45260# 0.032207f
C12349 a_n755_45592# a_n37_45144# 0.050738f
C12350 a_n863_45724# a_2680_45002# 0.024737f
C12351 a_18597_46090# a_21381_43940# 0.080234f
C12352 a_15227_44166# a_17061_44734# 0.07208f
C12353 a_13259_45724# a_13348_45260# 0.016055f
C12354 a_n2661_45546# a_4558_45348# 0.050441f
C12355 a_n881_46662# a_768_44030# 0.057002f
C12356 a_4883_46098# a_n2293_46634# 0.046481f
C12357 a_2063_45854# a_7715_46873# 0.178294f
C12358 a_22959_47212# a_21588_30879# 0.018188f
C12359 a_6491_46660# a_4646_46812# 0.042695f
C12360 a_22400_42852# a_22537_39537# 0.019618f
C12361 a_20974_43370# a_4190_30871# 0.214288f
C12362 a_8791_43396# a_9145_43396# 0.092458f
C12363 a_22612_30879# a_17364_32525# 0.062457f
C12364 a_526_44458# a_453_43940# 0.028123f
C12365 a_n2661_45010# a_626_44172# 0.0195f
C12366 a_n2293_45010# a_375_42282# 0.021456f
C12367 a_n443_42852# a_9313_44734# 0.02484f
C12368 a_9290_44172# a_10807_43548# 0.364112f
C12369 a_8746_45002# a_10440_44484# 0.027688f
C12370 a_n237_47217# a_8034_45724# 0.0717f
C12371 a_4883_46098# a_9625_46129# 0.164961f
C12372 a_11599_46634# a_18189_46348# 0.101491f
C12373 a_13661_43548# a_11415_45002# 0.107787f
C12374 a_13747_46662# a_20202_43084# 0.308003f
C12375 a_n881_46662# a_1176_45822# 0.048496f
C12376 a_10227_46804# a_13759_46122# 0.920747f
C12377 a_8530_39574# VDAC_P 0.064895f
C12378 a_13887_32519# a_5534_30871# 0.047233f
C12379 a_5649_42852# a_5342_30871# 0.091782f
C12380 a_2075_43172# a_2905_42968# 0.023236f
C12381 a_9482_43914# a_n2661_42834# 0.076592f
C12382 a_n755_45592# a_104_43370# 0.029812f
C12383 a_10903_43370# a_743_42282# 0.029178f
C12384 a_20193_45348# a_20205_45028# 0.012189f
C12385 a_10193_42453# a_14021_43940# 0.033291f
C12386 a_n2312_40392# a_n4318_38216# 0.025276f
C12387 a_11599_46634# a_17478_45572# 0.025658f
C12388 a_3090_45724# a_526_44458# 0.058033f
C12389 a_n2293_46098# a_1138_42852# 0.029886f
C12390 a_16327_47482# a_16115_45572# 0.163022f
C12391 a_8270_45546# a_8034_45724# 0.031124f
C12392 a_n901_46420# a_n1076_46494# 0.234322f
C12393 a_16388_46812# a_15682_46116# 0.044769f
C12394 a_1799_45572# a_1848_45724# 0.080562f
C12395 a_n971_45724# a_2437_43646# 0.204278f
C12396 a_n2840_42826# a_n4318_38216# 0.012711f
C12397 a_10991_42826# a_11554_42852# 0.049827f
C12398 a_n2472_42826# a_n2472_42282# 0.025171f
C12399 a_n1059_45260# a_8791_43396# 0.196029f
C12400 a_18494_42460# a_20269_44172# 0.017863f
C12401 a_n2293_43922# a_11967_42832# 0.022597f
C12402 a_2382_45260# a_3626_43646# 0.041715f
C12403 a_3065_45002# a_2982_43646# 0.026494f
C12404 a_5883_43914# a_7845_44172# 0.02286f
C12405 a_n1741_47186# VDD 0.912651f
C12406 a_20820_30879# a_14097_32519# 0.052932f
C12407 a_n2497_47436# CLK_DATA 0.026654f
C12408 a_n2438_43548# a_1423_45028# 0.242599f
C12409 a_11453_44696# a_11827_44484# 0.170003f
C12410 a_12465_44636# a_11691_44458# 0.15589f
C12411 a_12741_44636# a_13249_42308# 0.028381f
C12412 a_3090_45724# a_17668_45572# 0.071363f
C12413 a_5937_45572# a_2711_45572# 0.063757f
C12414 a_13059_46348# a_8696_44636# 0.020156f
C12415 a_3877_44458# a_3232_43370# 0.016642f
C12416 a_n2956_39304# a_n2810_45572# 0.043323f
C12417 a_11823_42460# a_14635_42282# 0.087526f
C12418 a_20193_45348# a_22223_43396# 0.020364f
C12419 a_10949_43914# a_11750_44172# 0.05299f
C12420 a_7832_46660# VDD 0.077608f
C12421 a_11967_42832# a_n97_42460# 0.489711f
C12422 a_895_43940# a_2253_43940# 0.053882f
C12423 a_2479_44172# a_2455_43940# 0.025354f
C12424 a_2324_44458# a_14180_45002# 0.026932f
C12425 a_6945_45028# a_6709_45028# 0.060282f
C12426 a_10053_45546# a_8746_45002# 0.075884f
C12427 a_10180_45724# a_10193_42453# 0.145672f
C12428 a_526_44458# a_2274_45254# 0.019853f
C12429 a_22612_30879# a_19237_31679# 0.062542f
C12430 a_12861_44030# a_15493_43940# 0.370814f
C12431 a_768_44030# a_2889_44172# 0.011283f
C12432 a_n971_45724# a_n2661_46634# 0.190714f
C12433 a_n443_46116# a_768_44030# 0.177051f
C12434 a_4915_47217# a_12549_44172# 0.316329f
C12435 a_9067_47204# a_n881_46662# 0.073421f
C12436 a_n2497_47436# a_n2438_43548# 0.206216f
C12437 a_n1920_47178# a_n1925_46634# 0.013665f
C12438 a_18597_46090# a_4883_46098# 0.084375f
C12439 a_5742_30871# a_4958_30871# 0.032374f
C12440 a_15959_42545# a_15890_42674# 0.209641f
C12441 a_3905_42865# a_3935_42891# 0.240349f
C12442 a_10586_45546# VDD 0.582083f
C12443 a_2711_45572# a_11691_44458# 0.058464f
C12444 a_n2293_46634# a_8685_43396# 0.335608f
C12445 a_n755_45592# a_949_44458# 0.011024f
C12446 a_22959_45572# a_20447_31679# 0.154273f
C12447 a_5257_43370# a_n97_42460# 0.167676f
C12448 a_8696_44636# a_13556_45296# 0.022968f
C12449 a_16147_45260# a_6171_45002# 0.072853f
C12450 a_12549_44172# a_15681_43442# 0.080982f
C12451 a_13507_46334# a_20107_46660# 0.031344f
C12452 a_3877_44458# a_4651_46660# 0.032518f
C12453 a_2063_45854# a_4419_46090# 0.025095f
C12454 a_3160_47472# a_3147_46376# 0.208295f
C12455 a_2905_45572# a_3483_46348# 0.024106f
C12456 a_12549_44172# a_18834_46812# 0.01219f
C12457 a_12861_44030# a_12741_44636# 0.366155f
C12458 a_4883_46098# a_19123_46287# 0.022559f
C12459 a_n971_45724# a_8199_44636# 0.247183f
C12460 a_n237_47217# a_8016_46348# 0.017823f
C12461 a_n443_46116# a_1176_45822# 0.092452f
C12462 a_n4209_38502# a_n4209_37414# 0.028607f
C12463 a_5742_30871# VCM 0.211981f
C12464 a_7174_31319# EN_VIN_BSTR_N 0.051994f
C12465 a_20447_31679# RST_Z 0.050985f
C12466 a_743_42282# a_5649_42852# 0.030921f
C12467 a_2437_43646# DATA[3] 0.075788f
C12468 a_4190_30871# a_13887_32519# 0.032018f
C12469 a_3232_43370# a_10440_44484# 0.042872f
C12470 a_20107_46660# a_20623_46660# 0.105914f
C12471 a_8270_45546# a_8016_46348# 0.036831f
C12472 a_13661_43548# a_13259_45724# 0.250875f
C12473 RST_Z START 0.033428f
C12474 C0_dummy_P_btm VCM 0.311452f
C12475 C0_N_btm VREF 0.443884f
C12476 C1_N_btm VIN_N 0.39234f
C12477 VDD SINGLE_ENDED 0.210835f
C12478 a_3539_42460# a_3905_42558# 0.015463f
C12479 a_2711_45572# a_4190_30871# 0.051595f
C12480 a_20193_45348# a_20512_43084# 0.160912f
C12481 a_8375_44464# a_5891_43370# 0.094782f
C12482 a_n357_42282# a_n13_43084# 0.194173f
C12483 a_10903_43370# a_8049_45260# 0.114138f
C12484 a_19692_46634# a_10193_42453# 0.010323f
C12485 a_15368_46634# a_11823_42460# 0.014491f
C12486 a_768_44030# a_3537_45260# 0.341201f
C12487 a_n1613_43370# a_7229_43940# 0.059621f
C12488 a_4185_45028# a_13259_45724# 0.194989f
C12489 a_5013_44260# a_5495_43940# 0.251039f
C12490 a_20362_44736# a_20365_43914# 0.012553f
C12491 a_3537_45260# a_5755_42852# 0.088502f
C12492 a_n913_45002# a_13113_42826# 0.018663f
C12493 a_19279_43940# a_19328_44172# 0.120319f
C12494 a_n743_46660# VDD 1.75634f
C12495 a_22612_30879# EN_OFFSET_CAL 0.118817f
C12496 a_1823_45246# a_3065_45002# 0.607468f
C12497 a_3147_46376# a_413_45260# 0.015235f
C12498 a_11415_45002# a_13159_45002# 0.141106f
C12499 a_17701_42308# VDD 0.243354f
C12500 a_6545_47178# a_6491_46660# 0.181574f
C12501 a_4915_47217# a_6575_47204# 0.849579f
C12502 a_2063_45854# a_11599_46634# 0.19861f
C12503 a_6761_42308# a_6123_31319# 0.187371f
C12504 a_3422_30871# a_4361_42308# 0.096125f
C12505 a_n2956_37592# a_n3674_38680# 0.02294f
C12506 a_n2956_38216# a_n4064_37984# 0.054267f
C12507 a_n2017_45002# a_n1736_42282# 0.017988f
C12508 a_11189_46129# VDD 0.944289f
C12509 a_18175_45572# a_18341_45572# 0.577068f
C12510 a_n2661_45546# a_n2661_43370# 0.145941f
C12511 a_13259_45724# a_18587_45118# 0.099974f
C12512 a_8199_44636# a_9313_44734# 0.016063f
C12513 a_4185_45028# a_n2661_43922# 0.022579f
C12514 a_16375_45002# a_17613_45144# 0.040514f
C12515 a_9049_44484# a_6171_45002# 0.026882f
C12516 a_n1925_42282# a_n699_43396# 0.024581f
C12517 a_n1925_46634# a_n1021_46688# 0.011448f
C12518 a_n2104_46634# a_n2438_43548# 0.052991f
C12519 a_n1613_43370# a_5907_46634# 0.338694f
C12520 a_n1151_42308# a_14035_46660# 0.026112f
C12521 a_4883_46098# a_6755_46942# 0.060162f
C12522 a_12861_44030# a_13607_46688# 0.019182f
C12523 a_n971_45724# a_765_45546# 0.140618f
C12524 a_1273_38525# a_2112_39137# 0.225378f
C12525 a_5932_42308# EN_VIN_BSTR_N 0.066129f
C12526 a_564_42282# VDD 0.293756f
C12527 a_11967_42832# a_12800_43218# 0.025258f
C12528 a_10907_45822# CLK 0.035046f
C12529 a_14401_32519# a_5534_30871# 0.339008f
C12530 a_5205_44484# a_n2661_43370# 0.033807f
C12531 a_n2661_45546# a_2998_44172# 0.060624f
C12532 a_n755_45592# a_175_44278# 0.01086f
C12533 a_13059_46348# a_14205_43396# 0.049915f
C12534 a_1138_42852# a_1209_43370# 0.01435f
C12535 a_14084_46812# a_14035_46660# 0.086342f
C12536 a_2063_45854# a_1848_45724# 0.057473f
C12537 a_n1151_42308# a_n1099_45572# 0.046104f
C12538 a_4883_46098# a_8049_45260# 0.469963f
C12539 a_11599_46634# a_14383_46116# 0.026426f
C12540 a_n743_46660# a_9823_46155# 0.196587f
C12541 a_12861_44030# a_16375_45002# 0.033138f
C12542 a_13747_46662# a_17715_44484# 0.025502f
C12543 a_12549_44172# a_10809_44734# 2.27272f
C12544 a_n1550_35448# a_n217_35014# 0.08192f
C12545 a_n1696_34930# EN_VIN_BSTR_P 0.336365f
C12546 VDAC_N C5_N_btm 27.606901f
C12547 a_16795_42852# a_17595_43084# 0.010079f
C12548 a_18479_45785# a_14021_43940# 0.025329f
C12549 a_n913_45002# a_n2661_42282# 0.054259f
C12550 a_10440_44484# a_8975_43940# 0.045841f
C12551 a_3232_43370# a_5244_44056# 0.017099f
C12552 a_n1917_44484# a_n1821_44484# 0.013793f
C12553 a_10355_46116# a_9290_44172# 0.01806f
C12554 a_12465_44636# a_2437_43646# 0.18195f
C12555 a_13747_46662# a_15861_45028# 0.021551f
C12556 a_4791_45118# a_7229_43940# 0.026326f
C12557 a_11750_44172# VDD 0.131662f
C12558 a_4361_42308# a_15803_42450# 0.055869f
C12559 a_13556_45296# a_14205_43396# 0.012255f
C12560 a_20193_45348# a_21381_43940# 0.01388f
C12561 a_21177_47436# VDD 0.179587f
C12562 a_11415_45002# a_20273_45572# 0.01364f
C12563 a_n2497_47436# a_n1741_47186# 0.098118f
C12564 a_4361_42308# VDD 0.42717f
C12565 a_13467_32519# RST_Z 0.048721f
C12566 a_14209_32519# C5_N_btm 0.042017f
C12567 a_196_42282# a_n1794_35082# 0.032791f
C12568 a_2479_44172# a_2982_43646# 0.019219f
C12569 a_5343_44458# a_8037_42858# 0.019942f
C12570 a_14955_43940# a_15037_43940# 0.171361f
C12571 a_20841_46902# VDD 0.20446f
C12572 a_n755_45592# a_n143_45144# 0.07862f
C12573 a_n863_45724# a_2382_45260# 0.119625f
C12574 a_n2661_45546# a_4574_45260# 0.014727f
C12575 a_310_45028# a_413_45260# 0.025313f
C12576 a_15227_44166# a_16241_44734# 0.105126f
C12577 a_13259_45724# a_13159_45002# 0.047761f
C12578 a_2063_45854# a_7411_46660# 0.029159f
C12579 a_4791_45118# a_5907_46634# 0.016954f
C12580 a_n881_46662# a_12549_44172# 0.225257f
C12581 a_n1613_43370# a_768_44030# 0.028683f
C12582 SMPL_ON_N a_22612_30879# 5.22049f
C12583 a_11453_44696# a_21588_30879# 0.075738f
C12584 a_6491_46660# a_3877_44458# 0.02519f
C12585 a_6545_47178# a_4646_46812# 0.02302f
C12586 a_22400_42852# a_22889_38993# 0.13715f
C12587 a_21613_42308# a_22775_42308# 0.225363f
C12588 a_20974_43370# a_21259_43561# 0.049502f
C12589 a_14401_32519# a_4190_30871# 0.10855f
C12590 a_n4318_40392# a_n3674_38216# 0.023361f
C12591 a_n2293_43922# a_n2293_42282# 0.19201f
C12592 a_21588_30879# a_17364_32525# 0.05857f
C12593 a_4927_45028# a_5691_45260# 0.018415f
C12594 a_5111_44636# a_3232_43370# 0.134191f
C12595 a_526_44458# a_1414_42308# 0.097596f
C12596 a_3483_46348# a_11341_43940# 0.017129f
C12597 a_13259_45724# a_11967_42832# 0.141918f
C12598 a_9290_44172# a_10949_43914# 0.113864f
C12599 a_8746_45002# a_10334_44484# 0.019787f
C12600 a_n881_46662# a_1208_46090# 0.076994f
C12601 a_4883_46098# a_8953_45546# 0.078639f
C12602 a_11599_46634# a_17715_44484# 0.031427f
C12603 a_768_44030# a_n2293_46098# 0.039783f
C12604 a_5807_45002# a_11415_45002# 0.05094f
C12605 a_8530_39574# a_8912_37509# 0.426772f
C12606 a_7754_38470# VDAC_P 0.063714f
C12607 a_n4064_39616# VCM 0.068103f
C12608 a_13678_32519# a_5342_30871# 0.028488f
C12609 a_n2661_42282# a_1755_42282# 0.145244f
C12610 a_4190_30871# a_18817_42826# 0.011301f
C12611 a_1847_42826# a_2905_42968# 0.097535f
C12612 a_n755_45592# a_n97_42460# 1.02989f
C12613 a_n357_42282# a_104_43370# 0.026213f
C12614 a_22959_45036# a_19721_31679# 0.156264f
C12615 a_n2312_39304# a_n3674_38680# 0.023326f
C12616 a_n2293_46098# a_1176_45822# 0.027035f
C12617 a_16327_47482# a_16333_45814# 0.168559f
C12618 a_n2661_46634# a_2711_45572# 0.032616f
C12619 a_10796_42968# a_11554_42852# 0.056391f
C12620 a_10991_42826# a_11301_43218# 0.013793f
C12621 a_743_42282# a_1067_42314# 0.010185f
C12622 a_2982_43646# a_19511_42282# 0.014171f
C12623 a_n1920_47178# VDD 0.229556f
C12624 a_18494_42460# a_19862_44208# 0.019692f
C12625 a_n2833_47464# CLK_DATA 0.331592f
C12626 a_5111_44636# a_4905_42826# 0.128918f
C12627 a_5883_43914# a_7542_44172# 0.187537f
C12628 a_11691_44458# a_15682_43940# 0.013321f
C12629 a_8199_44636# a_2711_45572# 0.098064f
C12630 a_19466_46812# a_18341_45572# 0.02497f
C12631 a_20193_45348# a_5649_42852# 0.052027f
C12632 a_10729_43914# a_11750_44172# 0.144893f
C12633 a_10949_43914# a_10807_43548# 0.034945f
C12634 a_895_43940# a_1443_43940# 0.016028f
C12635 a_2127_44172# a_2455_43940# 0.096132f
C12636 a_2479_44172# a_2253_43940# 0.010537f
C12637 a_11823_42460# a_13291_42460# 0.257506f
C12638 a_5257_43370# a_n2661_43922# 0.030003f
C12639 a_10053_45546# a_10193_42453# 0.086012f
C12640 a_21588_30879# a_19237_31679# 0.055917f
C12641 a_9049_44484# a_8746_45002# 0.025877f
C12642 a_768_44030# a_2675_43914# 0.026212f
C12643 a_16327_47482# a_15493_43396# 0.025969f
C12644 a_4915_47217# a_12891_46348# 0.156543f
C12645 a_4791_45118# a_768_44030# 0.03019f
C12646 a_6575_47204# a_n881_46662# 0.708623f
C12647 a_n2109_47186# a_n1925_46634# 0.033276f
C12648 a_20894_47436# a_20990_47178# 0.313533f
C12649 a_5934_30871# a_7174_31319# 0.473128f
C12650 a_n3674_38680# a_n3420_38528# 0.07337f
C12651 a_15803_42450# a_15890_42674# 0.07009f
C12652 a_n3674_37592# a_n4064_39072# 0.019349f
C12653 a_4699_43561# a_3080_42308# 0.223965f
C12654 a_1568_43370# a_1427_43646# 0.046825f
C12655 a_3905_42865# a_3681_42891# 0.101054f
C12656 en_comp a_5742_30871# 0.092249f
C12657 a_11322_45546# a_n2661_43370# 0.01285f
C12658 a_n357_42282# a_949_44458# 0.016511f
C12659 a_19963_31679# a_20447_31679# 0.069779f
C12660 a_1138_42852# a_895_43940# 0.017458f
C12661 a_19692_46634# a_14021_43940# 0.775991f
C12662 a_8696_44636# a_9482_43914# 0.042504f
C12663 a_10227_46804# a_20731_47026# 0.016434f
C12664 a_3877_44458# a_4646_46812# 0.056449f
C12665 a_2063_45854# a_4185_45028# 0.023928f
C12666 a_2905_45572# a_3147_46376# 0.02017f
C12667 a_12549_44172# a_17609_46634# 0.487224f
C12668 a_12465_44636# a_765_45546# 0.019565f
C12669 a_4883_46098# a_18285_46348# 0.026239f
C12670 a_n971_45724# a_8349_46414# 0.01782f
C12671 a_n237_47217# a_7920_46348# 0.059304f
C12672 a_15890_42674# VDD 0.203548f
C12673 a_5742_30871# VREF_GND 0.191352f
C12674 a_8685_43396# a_15279_43071# 0.011343f
C12675 a_2437_43646# DATA[2] 0.046972f
C12676 a_21487_43396# a_4361_42308# 0.077645f
C12677 a_20447_31679# VDD 0.671143f
C12678 a_3232_43370# a_10334_44484# 0.040395f
C12679 a_8953_45546# a_8685_43396# 0.062741f
C12680 a_20411_46873# a_20273_46660# 0.219954f
C12681 a_20107_46660# a_20841_46902# 0.053479f
C12682 a_n881_46662# a_n2661_45546# 0.02866f
C12683 a_5807_45002# a_13259_45724# 0.096565f
C12684 C0_P_btm VCM 0.717283f
C12685 C0_N_btm VIN_N 0.529671f
C12686 VDD START 0.114358f
C12687 a_n97_42460# a_9885_42558# 0.011255f
C12688 a_5891_43370# VDD 2.12137f
C12689 a_7640_43914# a_5891_43370# 0.011186f
C12690 a_n2293_46098# a_n2472_45546# 0.015672f
C12691 a_n881_46662# a_5205_44484# 0.013688f
C12692 a_14976_45028# a_11823_42460# 0.010375f
C12693 a_18533_43940# VDD 0.182147f
C12694 a_5244_44056# a_5495_43940# 0.107037f
C12695 a_3537_45260# a_5111_42852# 0.123919f
C12696 a_n913_45002# a_12545_42858# 0.548984f
C12697 a_n1021_46688# VDD 0.226043f
C12698 a_21588_30879# EN_OFFSET_CAL 0.047538f
C12699 a_13259_45724# a_15143_45578# 0.060775f
C12700 a_1823_45246# a_2680_45002# 0.073588f
C12701 a_11415_45002# a_13017_45260# 0.100288f
C12702 a_6151_47436# a_6491_46660# 0.31912f
C12703 a_4915_47217# a_7903_47542# 0.042037f
C12704 a_17595_43084# VDD 0.168112f
C12705 a_6761_42308# a_7227_42308# 0.173849f
C12706 a_5932_42308# a_5934_30871# 1.37963f
C12707 a_3422_30871# a_13467_32519# 0.421402f
C12708 a_n2956_38216# a_n2946_37984# 0.150404f
C12709 a_n2810_45028# a_n3674_38680# 0.022953f
C12710 a_9290_44172# VDD 2.74561f
C12711 a_20202_43084# a_11967_42832# 0.02752f
C12712 a_18175_45572# a_18479_45785# 0.280208f
C12713 a_13259_45724# a_18315_45260# 0.144632f
C12714 a_4185_45028# a_n2661_42834# 0.023267f
C12715 a_16375_45002# a_17023_45118# 0.014031f
C12716 a_n1925_42282# a_4223_44672# 0.053508f
C12717 a_9049_44484# a_3232_43370# 0.17048f
C12718 a_7499_43078# a_6171_45002# 0.029896f
C12719 a_526_44458# a_n699_43396# 0.285f
C12720 a_n2293_46634# a_n2438_43548# 0.807205f
C12721 a_n1613_43370# a_5167_46660# 0.177362f
C12722 a_n2661_46634# a_33_46660# 0.050833f
C12723 a_n1151_42308# a_13885_46660# 0.333314f
C12724 a_4883_46098# a_10249_46116# 0.01923f
C12725 a_n4315_30879# a_n3420_37984# 0.034791f
C12726 a_n3674_37592# VDD 0.357168f
C12727 a_n4064_39072# a_n2302_39072# 0.250408f
C12728 a_n4064_40160# a_n3565_38216# 0.02828f
C12729 a_n4064_39616# a_n4064_38528# 0.05063f
C12730 a_n863_45724# a_453_43940# 0.02533f
C12731 a_8191_45002# a_8560_45348# 0.03364f
C12732 a_13059_46348# a_14358_43442# 0.041731f
C12733 a_14084_46812# a_13885_46660# 0.237373f
C12734 a_n2661_46634# a_12005_46116# 0.038027f
C12735 a_5807_45002# a_18189_46348# 0.033239f
C12736 a_12891_46348# a_10809_44734# 0.102888f
C12737 a_768_44030# a_6945_45028# 0.014703f
C12738 a_n743_46660# a_9569_46155# 0.104962f
C12739 a_n443_46116# a_n2661_45546# 0.136593f
C12740 a_n1696_34930# a_n1057_35014# 0.419419f
C12741 a_n1550_35448# EN_VIN_BSTR_P 0.573018f
C12742 VDAC_N C4_N_btm 13.8047f
C12743 a_n4318_39304# a_n4318_38216# 0.023477f
C12744 a_5111_44636# a_5495_43940# 0.037006f
C12745 a_5147_45002# a_5663_43940# 0.019985f
C12746 a_n1059_45260# a_n2661_42282# 0.028862f
C12747 a_10903_43370# a_5534_30871# 0.134296f
C12748 a_10440_44484# a_10057_43914# 0.026774f
C12749 a_10334_44484# a_8975_43940# 0.044798f
C12750 a_3232_43370# a_3905_42865# 0.027169f
C12751 a_n2312_38680# a_n3674_37592# 0.026177f
C12752 a_n1641_46494# a_n1545_46494# 0.013793f
C12753 a_13717_47436# a_413_45260# 4.36729f
C12754 a_13507_46334# a_3357_43084# 0.050295f
C12755 a_21811_47423# a_2437_43646# 0.025192f
C12756 a_n971_45724# a_1307_43914# 0.019541f
C12757 a_13661_43548# a_15861_45028# 0.047089f
C12758 a_13747_46662# a_8696_44636# 0.02273f
C12759 a_5342_30871# a_n1794_35082# 0.035143f
C12760 a_10807_43548# VDD 0.68049f
C12761 a_3422_30871# a_22315_44484# 0.19914f
C12762 a_19479_31679# a_13678_32519# 0.051236f
C12763 a_20990_47178# VDD 0.210484f
C12764 a_19787_47423# START 0.220891f
C12765 a_22612_30879# VDAC_N 0.011363f
C12766 a_n1059_45260# a_16823_43084# 0.318918f
C12767 a_19963_31679# a_13467_32519# 0.051345f
C12768 a_10809_44734# a_11322_45546# 0.22629f
C12769 a_20623_46660# a_3357_43084# 0.013905f
C12770 a_11415_45002# a_20107_45572# 0.019157f
C12771 a_22000_46634# a_2437_43646# 0.010034f
C12772 a_10227_46804# a_9313_44734# 0.875947f
C12773 a_15227_44166# a_6171_45002# 0.021072f
C12774 a_13467_32519# VDD 0.354212f
C12775 a_n2497_47436# a_n1920_47178# 0.049461f
C12776 a_n2288_47178# a_n2109_47186# 0.177673f
C12777 a_n784_42308# a_n3674_37592# 0.254719f
C12778 a_n473_42460# a_n1794_35082# 0.049561f
C12779 a_3905_42865# a_4905_42826# 0.404829f
C12780 a_2479_44172# a_2896_43646# 0.026857f
C12781 a_1414_42308# a_3626_43646# 0.015112f
C12782 a_5343_44458# a_7765_42852# 0.010279f
C12783 a_20273_46660# VDD 0.247553f
C12784 a_n755_45592# a_n467_45028# 0.26002f
C12785 a_n863_45724# a_2274_45254# 0.17549f
C12786 a_n2661_45546# a_3537_45260# 0.780422f
C12787 a_n1925_42282# a_n2293_42834# 0.024873f
C12788 a_18189_46348# a_18315_45260# 0.101775f
C12789 a_310_45028# a_n37_45144# 0.112458f
C12790 a_n443_46116# a_1427_43646# 0.05874f
C12791 a_10903_43370# a_11691_44458# 0.020718f
C12792 a_15227_44166# a_14673_44172# 0.357896f
C12793 a_13259_45724# a_13017_45260# 0.078313f
C12794 a_19321_45002# a_19862_44208# 0.090113f
C12795 a_10193_42453# a_16147_45260# 0.193225f
C12796 a_2063_45854# a_5257_43370# 0.426517f
C12797 a_n881_46662# a_12891_46348# 0.026595f
C12798 SMPL_ON_N a_21588_30879# 0.119776f
C12799 a_11453_44696# a_20916_46384# 0.021978f
C12800 a_6545_47178# a_3877_44458# 0.026367f
C12801 a_6151_47436# a_4646_46812# 0.153739f
C12802 a_13258_32519# a_22485_38105# 0.057047f
C12803 a_22400_42852# a_22613_38993# 0.038807f
C12804 a_8292_43218# VDD 0.08228f
C12805 a_21381_43940# a_4190_30871# 0.023285f
C12806 a_22612_30879# a_14209_32519# 0.059911f
C12807 a_5111_44636# a_5691_45260# 0.130044f
C12808 a_5147_45002# a_3232_43370# 0.253159f
C12809 a_n2661_45010# a_375_42282# 0.017053f
C12810 a_526_44458# a_1467_44172# 0.041836f
C12811 a_9290_44172# a_10729_43914# 0.042243f
C12812 a_n357_42282# a_n2293_43922# 0.02281f
C12813 a_n755_45592# a_n2661_43922# 0.037767f
C12814 a_n881_46662# a_805_46414# 0.011286f
C12815 a_n971_45724# a_8034_45724# 0.027525f
C12816 a_4883_46098# a_5937_45572# 0.015486f
C12817 a_11599_46634# a_17583_46090# 0.031836f
C12818 a_9067_47204# a_6945_45028# 0.014009f
C12819 a_3754_38470# a_11206_38545# 0.078412f
C12820 a_8530_39574# VDAC_N 0.06498f
C12821 a_7754_38470# a_8912_37509# 0.575911f
C12822 a_n2302_39072# VDD 0.355374f
C12823 a_n2302_37690# a_n2216_37690# 0.011479f
C12824 a_n4064_39616# VREF_GND 0.241027f
C12825 a_n2661_42282# a_1606_42308# 0.082268f
C12826 a_1847_42826# a_2075_43172# 0.103349f
C12827 a_5649_42852# a_5534_30871# 0.234793f
C12828 a_4190_30871# a_18249_42858# 0.029356f
C12829 a_1423_45028# a_5891_43370# 0.301629f
C12830 a_1307_43914# a_9313_44734# 0.021168f
C12831 a_13249_42308# a_11341_43940# 0.032308f
C12832 a_n755_45592# a_n447_43370# 0.017822f
C12833 a_n357_42282# a_n97_42460# 0.900712f
C12834 a_n2312_40392# a_n3674_38680# 0.025175f
C12835 a_10227_46804# a_15037_45618# 0.012118f
C12836 a_n1741_47186# a_3357_43084# 0.03857f
C12837 a_1799_45572# a_n755_45592# 0.024036f
C12838 a_n1423_46090# a_n1076_46494# 0.051162f
C12839 a_12359_47026# a_10809_44734# 0.010386f
C12840 a_13059_46348# a_2324_44458# 0.0606f
C12841 a_11415_45002# a_3483_46348# 0.057381f
C12842 a_16327_47482# a_15765_45572# 0.048221f
C12843 a_10835_43094# a_11554_42852# 0.086334f
C12844 a_n2840_42826# a_n3674_38680# 0.019613f
C12845 a_22315_44484# VDD 0.213791f
C12846 a_13467_32519# a_n784_42308# 0.014901f
C12847 a_3422_30871# RST_Z 0.0872f
C12848 a_2382_45260# a_2982_43646# 0.468592f
C12849 a_16922_45042# a_15493_43940# 0.019907f
C12850 a_n2109_47186# VDD 2.71791f
C12851 a_3232_43370# a_4093_43548# 0.091441f
C12852 a_18184_42460# a_19862_44208# 0.028217f
C12853 a_5883_43914# a_7281_43914# 0.029594f
C12854 a_n2438_43548# a_626_44172# 0.025123f
C12855 a_10903_43370# a_n443_42852# 0.176275f
C12856 a_4646_46812# a_5111_44636# 0.078281f
C12857 a_n2293_42282# a_3318_42354# 0.01699f
C12858 a_20193_45348# a_13678_32519# 0.055785f
C12859 a_10729_43914# a_10807_43548# 0.238591f
C12860 a_895_43940# a_1241_43940# 0.054548f
C12861 a_2127_44172# a_2253_43940# 0.143754f
C12862 a_n755_45592# a_3318_42354# 0.152654f
C12863 a_12741_44636# a_16922_45042# 0.139755f
C12864 a_5257_43370# a_n2661_42834# 0.01982f
C12865 a_10053_45546# a_10180_45724# 0.144403f
C12866 a_2324_44458# a_13556_45296# 0.026317f
C12867 a_7499_43078# a_8746_45002# 0.153858f
C12868 a_12861_44030# a_11341_43940# 0.064865f
C12869 a_526_44458# a_327_44734# 0.076983f
C12870 a_6667_45809# a_6977_45572# 0.013793f
C12871 a_768_44030# a_895_43940# 0.06559f
C12872 a_22612_30879# a_17730_32519# 0.060497f
C12873 a_10227_46804# a_12465_44636# 0.057431f
C12874 a_18597_46090# a_13507_46334# 0.093881f
C12875 a_18479_47436# a_4883_46098# 0.038695f
C12876 SMPL_ON_P a_n2442_46660# 0.092029f
C12877 a_2063_45854# a_5807_45002# 0.074286f
C12878 a_4915_47217# a_11309_47204# 0.045252f
C12879 a_6151_47436# a_9804_47204# 0.095181f
C12880 a_7903_47542# a_n881_46662# 0.178742f
C12881 a_n3674_38680# a_n3690_38528# 0.071909f
C12882 COMP_P comp_n 0.032515f
C12883 a_15764_42576# a_15890_42674# 0.181217f
C12884 a_15803_42450# a_15959_42545# 0.110532f
C12885 a_15493_43940# a_15743_43084# 0.206331f
C12886 a_1049_43396# a_1427_43646# 0.010711f
C12887 a_4235_43370# a_3080_42308# 0.098951f
C12888 a_2437_43646# a_n2661_45010# 0.15182f
C12889 a_n755_45592# a_n452_44636# 0.015469f
C12890 a_n357_42282# a_742_44458# 0.085409f
C12891 a_4791_45118# a_5111_42852# 0.012003f
C12892 a_19963_31679# a_22959_45572# 0.020087f
C12893 a_17715_44484# a_11967_42832# 0.081495f
C12894 a_13507_46334# a_743_42282# 0.026943f
C12895 a_13507_46334# a_19123_46287# 0.034113f
C12896 a_12549_44172# a_16292_46812# 0.013094f
C12897 a_n237_47217# a_6419_46155# 0.029086f
C12898 a_n971_45724# a_8016_46348# 0.029312f
C12899 a_15959_42545# VDD 0.19373f
C12900 a_4190_30871# a_5649_42852# 0.434284f
C12901 a_21487_43396# a_13467_32519# 0.152042f
C12902 a_22959_45572# VDD 0.304443f
C12903 a_3357_43084# SINGLE_ENDED 0.131897f
C12904 a_19963_31679# RST_Z 0.050135f
C12905 a_2437_43646# DATA[1] 0.014934f
C12906 w_10694_33990# a_n1794_35082# 1.3413f
C12907 a_3232_43370# a_10157_44484# 0.049345f
C12908 a_7229_43940# a_6298_44484# 0.028942f
C12909 a_10227_46804# a_2711_45572# 0.130695f
C12910 a_20107_46660# a_20273_46660# 0.608339f
C12911 a_4883_46098# a_n443_42852# 0.074259f
C12912 a_n1613_43370# a_n2661_45546# 0.029057f
C12913 C0_P_btm VREF_GND 0.350485f
C12914 C1_P_btm VCM 0.716121f
C12915 C0_dummy_N_btm VIN_N 0.544204f
C12916 VDD RST_Z 4.72787f
C12917 a_8375_44464# VDD 0.086619f
C12918 a_13249_42308# a_10341_43396# 0.040208f
C12919 a_n2472_46090# a_n2472_45546# 0.025171f
C12920 a_n2293_46098# a_n2661_45546# 3.03243f
C12921 a_n743_46660# a_3357_43084# 0.034228f
C12922 a_17339_46660# a_2711_45572# 0.02331f
C12923 a_n881_46662# a_6431_45366# 0.177591f
C12924 a_12465_44636# a_1307_43914# 0.022149f
C12925 a_n1613_43370# a_5205_44484# 0.551795f
C12926 a_768_44030# a_3065_45002# 0.288972f
C12927 a_3090_45724# a_11823_42460# 0.089008f
C12928 a_3483_46348# a_13259_45724# 0.230226f
C12929 a_14401_32519# C6_N_btm 0.054459f
C12930 a_19319_43548# VDD 0.561461f
C12931 a_5244_44056# a_5013_44260# 0.094334f
C12932 a_3537_45260# a_4520_42826# 0.066648f
C12933 a_n913_45002# a_12089_42308# 0.038293f
C12934 a_n1059_45260# a_12545_42858# 0.011705f
C12935 a_n1925_46634# VDD 0.783093f
C12936 a_4185_45028# a_17303_42282# 0.235259f
C12937 a_n2442_46660# CLK_DATA 0.063913f
C12938 a_1823_45246# a_2382_45260# 0.801932f
C12939 a_13259_45724# a_14495_45572# 0.020864f
C12940 a_167_45260# a_1667_45002# 0.05322f
C12941 a_11415_45002# a_11963_45334# 0.031636f
C12942 a_6151_47436# a_6545_47178# 0.39775f
C12943 a_4915_47217# a_7227_47204# 0.059062f
C12944 a_16795_42852# VDD 0.179044f
C12945 a_n2810_45572# a_n2302_37984# 0.130495f
C12946 a_n2017_45002# a_n2104_42282# 0.010745f
C12947 a_n2956_38216# a_n3420_37984# 0.208204f
C12948 a_10355_46116# VDD 0.222751f
C12949 a_9313_44734# a_13635_43156# 0.013436f
C12950 a_12861_44030# a_10341_43396# 0.018259f
C12951 a_13259_45724# a_17719_45144# 0.039832f
C12952 a_8016_46348# a_9313_44734# 0.020204f
C12953 a_3483_46348# a_n2661_43922# 0.038814f
C12954 a_2711_45572# a_1307_43914# 0.187968f
C12955 a_22612_30879# a_17538_32519# 0.060018f
C12956 a_16375_45002# a_16922_45042# 0.170835f
C12957 a_7499_43078# a_3232_43370# 0.318423f
C12958 a_n1613_43370# a_5385_46902# 0.182522f
C12959 a_13507_46334# a_6755_46942# 0.075659f
C12960 a_11599_46634# a_11813_46116# 0.106062f
C12961 a_n327_42558# VDD 0.198414f
C12962 a_n784_42308# RST_Z 0.033698f
C12963 a_1606_42308# C2_N_btm 0.021793f
C12964 a_n4064_40160# a_n4334_38304# 0.013157f
C12965 a_10341_43396# a_19700_43370# 0.013451f
C12966 a_5343_44458# a_8325_42308# 0.014133f
C12967 a_n863_45724# a_1414_42308# 0.711805f
C12968 a_6171_45002# a_n2661_43370# 2.37006f
C12969 a_13059_46348# a_14579_43548# 0.171744f
C12970 a_2711_45572# a_18579_44172# 0.170319f
C12971 a_n755_45592# a_n809_44244# 0.404418f
C12972 a_13607_46688# a_13885_46660# 0.11044f
C12973 a_n2661_46634# a_10903_43370# 0.663878f
C12974 a_13507_46334# a_8049_45260# 0.086137f
C12975 a_4791_45118# a_n2661_45546# 0.012117f
C12976 a_2063_45854# a_n755_45592# 0.074611f
C12977 a_n1613_43370# a_n1533_46116# 0.012221f
C12978 a_n743_46660# a_9625_46129# 0.206271f
C12979 a_12549_44172# a_6945_45028# 0.028827f
C12980 a_5807_45002# a_17715_44484# 0.045558f
C12981 a_n1550_35448# a_n1057_35014# 0.201872f
C12982 VDAC_N C3_N_btm 6.907279f
C12983 a_5111_44636# a_5013_44260# 0.029412f
C12984 a_5147_45002# a_5495_43940# 0.086203f
C12985 a_3232_43370# a_3600_43914# 0.087298f
C12986 a_n443_42852# a_8685_43396# 0.281116f
C12987 a_13249_42308# a_n97_42460# 0.067568f
C12988 a_n2017_45002# a_n2661_42282# 0.035164f
C12989 a_10157_44484# a_8975_43940# 0.045547f
C12990 a_n1917_44484# a_n1809_44850# 0.057222f
C12991 a_n2442_46660# a_n1794_35082# 0.02547f
C12992 a_n1641_46494# a_n1736_46482# 0.049827f
C12993 a_13059_46348# a_12839_46116# 0.098052f
C12994 a_16327_47482# a_n913_45002# 0.137194f
C12995 a_4915_47217# a_6171_45002# 0.022258f
C12996 a_n1435_47204# a_413_45260# 0.025027f
C12997 a_4883_46098# a_2437_43646# 0.458866f
C12998 a_13507_46334# a_19479_31679# 0.061466f
C12999 a_4791_45118# a_5205_44484# 0.053467f
C13000 a_13661_43548# a_8696_44636# 0.049791f
C13001 a_13747_46662# a_16680_45572# 0.047612f
C13002 a_10949_43914# VDD 0.797824f
C13003 a_19386_47436# START 0.042951f
C13004 a_n2293_42834# a_3539_42460# 0.019435f
C13005 a_20894_47436# VDD 0.188358f
C13006 a_5891_43370# a_10405_44172# 0.15894f
C13007 a_n743_46660# a_16237_45028# 0.038671f
C13008 a_22612_30879# a_19721_31679# 0.068873f
C13009 a_13259_45724# a_n357_42282# 0.056511f
C13010 a_768_44030# a_6298_44484# 0.015186f
C13011 a_4915_47217# a_14673_44172# 0.020025f
C13012 a_8034_45724# a_2711_45572# 0.035334f
C13013 a_10809_44734# a_10490_45724# 0.030973f
C13014 a_20205_31679# a_20692_30879# 0.055565f
C13015 a_n2497_47436# a_n2109_47186# 0.197671f
C13016 a_196_42282# a_n3674_37592# 0.1528f
C13017 a_n961_42308# a_n1794_35082# 0.028868f
C13018 a_3905_42865# a_3080_42308# 0.029566f
C13019 a_1414_42308# a_3540_43646# 0.022584f
C13020 a_5343_44458# a_7871_42858# 0.020081f
C13021 a_11967_42832# a_15095_43370# 0.098499f
C13022 a_13483_43940# a_13565_43940# 0.171361f
C13023 a_20411_46873# VDD 0.348821f
C13024 a_526_44458# a_n2293_42834# 1.7774f
C13025 a_13661_43548# a_20365_43914# 0.020045f
C13026 a_584_46384# a_648_43396# 0.050476f
C13027 a_n2293_45546# a_2382_45260# 0.078874f
C13028 a_n863_45724# a_1667_45002# 0.20954f
C13029 a_n443_46116# a_4817_46660# 0.020386f
C13030 a_n881_46662# a_11309_47204# 0.028783f
C13031 a_4883_46098# a_n2661_46634# 0.030655f
C13032 a_22731_47423# a_21588_30879# 0.014331f
C13033 a_6151_47436# a_3877_44458# 0.034088f
C13034 a_n1741_47186# a_6755_46942# 0.017537f
C13035 a_n3674_37592# a_n4064_37440# 0.651412f
C13036 a_22400_42852# a_22581_37893# 0.031385f
C13037 a_21887_42336# a_21613_42308# 0.071168f
C13038 a_n97_42460# a_19700_43370# 0.154491f
C13039 a_21381_43940# a_21259_43561# 0.013931f
C13040 a_n2956_37592# a_n4064_39616# 0.015429f
C13041 a_n4318_40392# a_n4318_38216# 0.023287f
C13042 a_5111_44636# a_4927_45028# 0.134309f
C13043 a_7499_43078# a_8975_43940# 0.519621f
C13044 a_21588_30879# a_14209_32519# 0.056208f
C13045 a_5147_45002# a_5691_45260# 0.035185f
C13046 a_n755_45592# a_n2661_42834# 0.059506f
C13047 a_n357_42282# a_n2661_43922# 0.088336f
C13048 a_n881_46662# a_472_46348# 0.022658f
C13049 a_4883_46098# a_8199_44636# 0.242f
C13050 a_11599_46634# a_15682_46116# 1.8289f
C13051 a_6755_46942# a_7832_46660# 0.025487f
C13052 a_584_46384# a_1337_46116# 0.044678f
C13053 a_6575_47204# a_6945_45028# 0.06375f
C13054 a_12861_44030# a_17957_46116# 0.01013f
C13055 a_3160_47472# a_526_44458# 0.026069f
C13056 a_3754_38470# VDAC_P 0.323951f
C13057 a_7754_38470# VDAC_N 0.110605f
C13058 a_8530_39574# a_6886_37412# 0.616015f
C13059 a_n4064_39072# VDD 1.74929f
C13060 a_n3420_39616# VCM 0.0424f
C13061 a_4361_42308# a_5342_30871# 0.047616f
C13062 a_743_42282# a_17701_42308# 0.014357f
C13063 a_13678_32519# a_5534_30871# 0.043974f
C13064 a_11967_42832# a_17303_42282# 0.058225f
C13065 a_1423_45028# a_8375_44464# 0.032906f
C13066 a_22223_45036# a_18114_32519# 0.15655f
C13067 a_n1991_46122# a_n1076_46494# 0.124988f
C13068 a_13059_46348# a_14840_46494# 0.031849f
C13069 a_n2840_42826# a_n2840_42282# 0.025171f
C13070 a_3422_30871# VDD 1.12305f
C13071 a_743_42282# a_564_42282# 0.169821f
C13072 a_19778_44110# a_19862_44208# 0.213467f
C13073 a_5883_43914# a_6453_43914# 0.051468f
C13074 a_n2288_47178# VDD 0.29372f
C13075 a_13507_46334# a_20193_45348# 0.253904f
C13076 a_15227_44166# a_18341_45572# 0.017357f
C13077 a_8016_46348# a_2711_45572# 0.028247f
C13078 a_4646_46812# a_5147_45002# 0.010619f
C13079 a_11415_45002# a_13249_42308# 0.071546f
C13080 a_8049_45260# a_10586_45546# 0.038262f
C13081 a_10729_43914# a_10949_43914# 0.418928f
C13082 a_n755_45592# a_2903_42308# 0.070479f
C13083 a_n443_42852# a_1067_42314# 0.011239f
C13084 a_3090_45724# a_14539_43914# 0.040638f
C13085 a_6945_45028# a_5205_44484# 0.058545f
C13086 a_n1613_43370# a_7281_43914# 0.030229f
C13087 a_7499_43078# a_10193_42453# 0.298293f
C13088 a_12861_44030# a_21115_43940# 0.035299f
C13089 a_10809_44734# a_6171_45002# 0.244599f
C13090 a_526_44458# a_413_45260# 0.103799f
C13091 a_768_44030# a_2479_44172# 0.056833f
C13092 a_21588_30879# a_17730_32519# 0.05582f
C13093 a_n1741_47186# a_n2442_46660# 0.014004f
C13094 a_6151_47436# a_8128_46384# 0.052868f
C13095 a_16327_47482# a_11453_44696# 0.038815f
C13096 a_n2497_47436# a_n1925_46634# 0.052533f
C13097 a_n3674_38680# a_n3565_38502# 0.128677f
C13098 a_15486_42560# a_15890_42674# 0.051162f
C13099 a_13575_42558# a_13921_42308# 0.013377f
C13100 a_15764_42576# a_15959_42545# 0.21686f
C13101 a_6123_31319# a_7174_31319# 13.9919f
C13102 a_n3674_37592# a_n3420_39072# 0.019892f
C13103 a_1049_43396# a_n1557_42282# 0.211757f
C13104 a_1209_43370# a_1427_43646# 0.08213f
C13105 a_4093_43548# a_3080_42308# 0.08049f
C13106 a_n863_45724# a_n699_43396# 0.23135f
C13107 a_18597_46090# a_4361_42308# 0.024928f
C13108 a_8270_45546# a_9801_43940# 0.014887f
C13109 a_8746_45002# a_n2661_43370# 0.052623f
C13110 a_n237_47217# a_6165_46155# 0.021223f
C13111 a_n443_46116# a_472_46348# 0.025699f
C13112 a_12861_44030# a_11415_45002# 0.081894f
C13113 a_13507_46334# a_18285_46348# 0.041986f
C13114 a_4883_46098# a_765_45546# 0.055532f
C13115 a_2063_45854# a_3483_46348# 0.164542f
C13116 a_n743_46660# a_6755_46942# 0.044888f
C13117 a_12549_44172# a_15559_46634# 0.012304f
C13118 a_13258_32519# EN_VIN_BSTR_N 0.040234f
C13119 a_15803_42450# VDD 0.448709f
C13120 a_5742_30871# VIN_N 0.042613f
C13121 a_7174_31319# EN_VIN_BSTR_P 0.052876f
C13122 a_743_42282# a_4361_42308# 7.66647f
C13123 a_4190_30871# a_13678_32519# 0.032285f
C13124 a_3357_43084# START 0.045418f
C13125 a_19963_31679# VDD 0.607916f
C13126 a_n356_44636# a_17124_42282# 0.025455f
C13127 a_3422_30871# a_n784_42308# 0.022792f
C13128 w_1575_34786# a_n1794_35082# 1.3413f
C13129 a_3232_43370# a_9838_44484# 0.053106f
C13130 a_3357_43084# a_5891_43370# 0.013053f
C13131 a_n913_45002# a_n356_44636# 0.640597f
C13132 a_8199_44636# a_8685_43396# 0.03394f
C13133 a_3090_45724# a_1823_45246# 0.038665f
C13134 a_20107_46660# a_20411_46873# 0.316529f
C13135 a_n743_46660# a_8049_45260# 2.07544f
C13136 C1_P_btm VREF_GND 0.673422f
C13137 C2_P_btm VCM 0.716172f
C13138 C0_P_btm VREF 0.443926f
C13139 a_7640_43914# VDD 0.196713f
C13140 a_4905_42826# a_5932_42308# 0.058059f
C13141 a_1307_43914# a_15682_43940# 0.028719f
C13142 a_11823_42460# a_12281_43396# 0.049968f
C13143 a_14539_43914# a_14815_43914# 0.099149f
C13144 a_n2293_46098# a_n2810_45572# 0.013787f
C13145 a_11453_44696# a_14537_43396# 0.029591f
C13146 a_20202_43084# a_n357_42282# 0.062522f
C13147 a_15227_44166# a_10193_42453# 0.205591f
C13148 a_n881_46662# a_6171_45002# 0.090566f
C13149 a_768_44030# a_2680_45002# 0.028861f
C13150 a_11189_46129# a_8049_45260# 0.03932f
C13151 a_n4318_38680# a_n4064_40160# 0.079598f
C13152 a_n2661_46634# DATA[0] 0.012107f
C13153 a_n2312_38680# VDD 0.540248f
C13154 a_4185_45028# a_4958_30871# 0.121495f
C13155 a_3905_42865# a_5013_44260# 0.182997f
C13156 a_13259_45724# a_22400_42852# 0.34531f
C13157 a_n913_45002# a_12379_42858# 0.066604f
C13158 a_n1059_45260# a_12089_42308# 0.022942f
C13159 a_n2293_46634# a_5891_43370# 0.105307f
C13160 a_n755_45592# a_3775_45552# 0.100709f
C13161 a_1823_45246# a_2274_45254# 0.255985f
C13162 a_13259_45724# a_13249_42308# 0.358931f
C13163 a_167_45260# a_327_44734# 0.199136f
C13164 a_11415_45002# a_11787_45002# 0.072246f
C13165 a_16414_43172# VDD 0.201389f
C13166 a_4915_47217# a_6851_47204# 0.172567f
C13167 a_6773_42558# a_6761_42308# 0.01129f
C13168 a_5932_42308# a_6123_31319# 1.49414f
C13169 a_10193_42453# a_7174_31319# 0.020527f
C13170 a_n2810_45572# a_n4064_37984# 0.094405f
C13171 a_n2956_38216# a_n3690_38304# 0.016795f
C13172 a_9823_46155# VDD 0.102474f
C13173 a_16147_45260# a_18175_45572# 0.108647f
C13174 a_526_44458# a_2779_44458# 0.090804f
C13175 a_3483_46348# a_n2661_42834# 0.0234f
C13176 a_2711_45572# a_16019_45002# 0.024255f
C13177 a_21588_30879# a_17538_32519# 0.055813f
C13178 a_n2661_46634# a_n133_46660# 0.022138f
C13179 a_n881_46662# a_4955_46873# 0.066882f
C13180 a_n1613_43370# a_4817_46660# 0.330391f
C13181 a_11599_46634# a_11735_46660# 0.268769f
C13182 a_n2104_46634# a_n1925_46634# 0.167849f
C13183 a_n784_42308# VDD 0.59759f
C13184 a_n4315_30879# a_n3565_38216# 0.043307f
C13185 a_1666_39587# a_2112_39137# 0.269764f
C13186 a_1606_42308# C1_N_btm 0.096405f
C13187 a_5932_42308# EN_VIN_BSTR_P 0.066893f
C13188 a_n4064_40160# a_n4209_38216# 0.047163f
C13189 a_n3420_39616# a_n4064_38528# 0.048102f
C13190 a_n4064_39616# a_n3420_38528# 0.052176f
C13191 a_n2946_39072# a_n4064_39072# 0.053263f
C13192 a_15781_43660# a_16137_43396# 0.089942f
C13193 a_10341_43396# a_19268_43646# 0.010402f
C13194 a_3232_43370# a_n2661_43370# 0.077167f
C13195 a_n863_45724# a_1467_44172# 0.021736f
C13196 a_n2293_46634# a_9290_44172# 0.102393f
C13197 a_n1151_42308# a_n863_45724# 0.081395f
C13198 a_12861_44030# a_13259_45724# 0.435853f
C13199 a_584_46384# a_n755_45592# 0.020619f
C13200 a_n743_46660# a_8953_45546# 0.062066f
C13201 a_12891_46348# a_6945_45028# 0.013255f
C13202 a_13747_46662# a_2324_44458# 0.025909f
C13203 a_n2302_37690# VDD 0.350119f
C13204 a_n1550_35448# a_n1696_34930# 0.04535f
C13205 VDAC_N C2_N_btm 3.46253f
C13206 a_n4318_39304# a_n3674_38680# 0.031218f
C13207 a_5147_45002# a_5013_44260# 0.189328f
C13208 a_3232_43370# a_2998_44172# 0.056614f
C13209 a_5111_44636# a_5244_44056# 0.01138f
C13210 a_n2661_44458# a_n356_44636# 0.055568f
C13211 a_10334_44484# a_10440_44484# 0.313533f
C13212 a_9838_44484# a_8975_43940# 0.055678f
C13213 a_n1917_44484# a_n2012_44484# 0.049827f
C13214 a_n1699_44726# a_n1809_44850# 0.097745f
C13215 a_4646_46812# a_7499_43078# 0.158236f
C13216 a_21496_47436# a_2437_43646# 0.01965f
C13217 a_13507_46334# a_22223_45572# 0.015966f
C13218 a_16327_47482# a_n1059_45260# 0.235708f
C13219 a_13747_46662# a_16855_45546# 0.02676f
C13220 a_5807_45002# a_8696_44636# 0.024228f
C13221 a_3483_46348# a_17715_44484# 0.059106f
C13222 a_743_42282# a_15890_42674# 0.010042f
C13223 a_10729_43914# VDD 0.681371f
C13224 a_5534_30871# a_n1794_35082# 0.033914f
C13225 a_4361_42308# a_15051_42282# 0.016131f
C13226 a_14537_43396# a_9145_43396# 0.129182f
C13227 a_n2293_42834# a_3626_43646# 0.019674f
C13228 a_18597_46090# START 0.020125f
C13229 a_1823_45246# a_3905_42558# 0.010516f
C13230 a_19787_47423# VDD 0.256911f
C13231 a_20273_46660# a_3357_43084# 0.02704f
C13232 a_21588_30879# a_19721_31679# 0.055771f
C13233 a_22612_30879# a_18114_32519# 0.061298f
C13234 a_10809_44734# a_8746_45002# 0.049227f
C13235 a_21487_43396# VDD 0.222231f
C13236 a_n2497_47436# a_n2288_47178# 0.067981f
C13237 a_n473_42460# a_n3674_37592# 0.054584f
C13238 a_n1329_42308# a_n1794_35082# 0.043579f
C13239 a_5891_43370# a_743_42282# 0.065685f
C13240 a_1414_42308# a_2982_43646# 0.071994f
C13241 a_20107_46660# VDD 0.442554f
C13242 a_13747_46662# a_19862_44208# 0.15289f
C13243 a_n2293_46634# a_10807_43548# 0.05087f
C13244 a_n971_45724# a_8147_43396# 0.116186f
C13245 a_n2293_45546# a_2274_45254# 0.07158f
C13246 a_n863_45724# a_327_44734# 0.353745f
C13247 a_n443_46116# a_4955_46873# 0.126551f
C13248 a_4791_45118# a_4817_46660# 0.020367f
C13249 a_22223_47212# a_21588_30879# 0.164932f
C13250 a_21335_42336# a_21613_42308# 0.110671f
C13251 a_9290_44172# a_9672_43914# 0.071844f
C13252 a_n2661_45010# a_1307_43914# 0.016415f
C13253 a_5147_45002# a_4927_45028# 0.168157f
C13254 a_7499_43078# a_10057_43914# 0.262644f
C13255 a_22612_30879# a_13887_32519# 0.060052f
C13256 a_n357_42282# a_n2661_42834# 0.239713f
C13257 a_n881_46662# a_376_46348# 0.016146f
C13258 a_11599_46634# a_2324_44458# 0.428445f
C13259 a_10227_46804# a_10903_43370# 0.041882f
C13260 a_2905_45572# a_526_44458# 0.142766f
C13261 a_7754_38470# a_6886_37412# 0.181496f
C13262 a_3754_38470# a_8912_37509# 1.88278f
C13263 a_n2946_39072# VDD 0.383374f
C13264 a_n3420_39616# VREF_GND 0.117023f
C13265 a_8530_39574# a_5700_37509# 0.947638f
C13266 a_13467_32519# a_5342_30871# 0.028573f
C13267 a_4190_30871# a_18083_42858# 0.023338f
C13268 a_11967_42832# a_4958_30871# 0.239255f
C13269 a_1423_45028# VDD 4.06861f
C13270 a_9290_44172# a_743_42282# 0.117511f
C13271 a_1423_45028# a_7640_43914# 0.105665f
C13272 a_8953_45546# a_4361_42308# 0.012234f
C13273 a_11827_44484# a_18114_32519# 0.09907f
C13274 a_n1853_46287# a_n1076_46494# 0.056078f
C13275 a_n1991_46122# a_n901_46420# 0.041816f
C13276 a_n2109_47186# a_3357_43084# 0.170493f
C13277 a_n1423_46090# a_n1641_46494# 0.209641f
C13278 a_16327_47482# a_15599_45572# 0.331892f
C13279 a_21398_44850# VDD 0.077608f
C13280 a_3626_43646# a_19332_42282# 0.013212f
C13281 a_19237_31679# C0_N_btm 0.040442f
C13282 a_4190_30871# a_n1794_35082# 0.039258f
C13283 a_3080_42308# a_7174_31319# 0.22305f
C13284 a_16922_45042# a_11341_43940# 0.028038f
C13285 a_6298_44484# a_7542_44172# 0.014735f
C13286 a_19778_44110# a_19478_44306# 0.099524f
C13287 a_5883_43914# a_5663_43940# 0.153361f
C13288 a_n2497_47436# VDD 1.33346f
C13289 a_15227_44166# a_18479_45785# 0.035756f
C13290 a_12465_44636# a_11827_44484# 0.785011f
C13291 a_n755_45592# a_2713_42308# 0.243663f
C13292 a_10405_44172# a_10949_43914# 0.05348f
C13293 a_10903_43370# a_1307_43914# 0.065094f
C13294 a_10809_44734# a_3232_43370# 0.158726f
C13295 a_3483_46348# a_5093_45028# 0.05597f
C13296 a_12861_44030# a_20935_43940# 0.02414f
C13297 SMPL_ON_P a_n2661_46634# 0.0112f
C13298 a_10227_46804# a_4883_46098# 0.200137f
C13299 a_18479_47436# a_13507_46334# 0.033523f
C13300 a_n3674_38680# a_n4334_38528# 0.05024f
C13301 a_15764_42576# a_15803_42450# 0.901878f
C13302 a_1209_43370# a_n1557_42282# 0.113851f
C13303 a_10807_43548# a_743_42282# 0.011093f
C13304 a_375_42282# a_n1794_35082# 0.036312f
C13305 a_19479_31679# a_20447_31679# 0.05179f
C13306 a_13507_46334# a_4190_30871# 0.186424f
C13307 a_22591_45572# a_19963_31679# 0.161955f
C13308 a_2711_45572# a_11827_44484# 0.033351f
C13309 a_1138_42852# a_453_43940# 0.018298f
C13310 a_15227_44166# a_14021_43940# 0.052407f
C13311 a_n1925_42282# a_n2293_43922# 2.06056f
C13312 a_n237_47217# a_5497_46414# 0.021428f
C13313 a_n443_46116# a_376_46348# 0.025241f
C13314 a_12861_44030# a_20202_43084# 0.020377f
C13315 a_4883_46098# a_17339_46660# 0.071433f
C13316 a_10227_46804# a_21188_46660# 0.22222f
C13317 a_12549_44172# a_15368_46634# 0.012256f
C13318 a_5807_45002# a_11813_46116# 0.037525f
C13319 a_5742_30871# VIN_P 0.042613f
C13320 a_15764_42576# VDD 0.258303f
C13321 a_n4064_39072# a_n4064_37440# 0.046264f
C13322 a_22485_38105# a_22629_38406# 0.206945f
C13323 a_3357_43084# RST_Z 0.031959f
C13324 a_22591_45572# VDD 0.314172f
C13325 a_3232_43370# a_5883_43914# 0.337937f
C13326 a_n1925_42282# a_n97_42460# 0.021883f
C13327 a_n1059_45260# a_n356_44636# 0.07487f
C13328 a_5205_44484# a_6298_44484# 0.085118f
C13329 a_7229_43940# a_5343_44458# 0.196399f
C13330 SMPL_ON_P COMP_P 0.03194f
C13331 C2_P_btm VREF_GND 0.671742f
C13332 C3_P_btm VCM 0.716273f
C13333 C1_P_btm VREF 0.98698f
C13334 C0_dummy_P_btm VIN_P 0.544204f
C13335 a_3422_30871# a_n4064_37440# 0.032121f
C13336 a_6109_44484# VDD 0.243629f
C13337 a_3626_43646# a_5379_42460# 0.057009f
C13338 a_n97_42460# a_9803_42558# 0.099148f
C13339 a_3080_42308# a_5932_42308# 14.0282f
C13340 a_11827_44484# a_22485_44484# 0.015798f
C13341 a_4883_46098# a_1307_43914# 0.026965f
C13342 a_n2438_43548# a_2437_43646# 0.045715f
C13343 a_n1925_46634# a_3357_43084# 0.034378f
C13344 a_n1613_43370# a_6171_45002# 0.026867f
C13345 a_768_44030# a_2382_45260# 0.094536f
C13346 a_9290_44172# a_8049_45260# 0.041148f
C13347 a_n3674_39304# a_n4064_40160# 0.024923f
C13348 a_n2104_46634# VDD 0.286113f
C13349 a_n913_45002# a_10341_42308# 0.070067f
C13350 a_n2017_45002# a_12089_42308# 0.043278f
C13351 a_n1925_42282# a_3823_42558# 0.010285f
C13352 a_16922_45042# a_10341_43396# 0.048996f
C13353 a_167_45260# a_413_45260# 0.120357f
C13354 a_1823_45246# a_1667_45002# 0.24808f
C13355 a_5815_47464# a_6151_47436# 0.235454f
C13356 a_4915_47217# a_6491_46660# 0.19739f
C13357 a_n1151_42308# a_9313_45822# 0.024431f
C13358 a_15567_42826# VDD 0.163583f
C13359 a_5342_30871# RST_Z 0.048618f
C13360 a_9569_46155# VDD 0.19288f
C13361 a_10193_42453# a_20712_42282# 0.157661f
C13362 a_n2810_45572# a_n2946_37984# 0.020842f
C13363 a_n2956_38216# a_n3565_38216# 0.307285f
C13364 a_16375_45002# a_16405_45348# 0.012425f
C13365 a_4883_46098# a_9396_43370# 0.172323f
C13366 a_526_44458# a_949_44458# 0.03455f
C13367 a_10809_44734# a_8975_43940# 0.169586f
C13368 a_10227_46804# a_8685_43396# 0.227547f
C13369 a_12861_44030# a_14955_43396# 0.024664f
C13370 a_n863_45724# a_n2293_42834# 0.107229f
C13371 a_22612_30879# a_14401_32519# 0.062739f
C13372 a_8953_45546# a_5891_43370# 0.321625f
C13373 a_n2661_46634# a_n2438_43548# 0.493975f
C13374 a_n1613_43370# a_4955_46873# 0.051259f
C13375 a_n2104_46634# a_n2312_38680# 0.154937f
C13376 a_n2293_46634# a_n1925_46634# 0.051324f
C13377 a_196_42282# VDD 0.291844f
C13378 a_1273_38525# a_1666_39043# 0.297741f
C13379 a_1606_42308# C0_N_btm 0.029189f
C13380 a_n3420_39072# a_n4064_39072# 4.91095f
C13381 a_n356_44636# a_1606_42308# 0.282657f
C13382 a_10341_43396# a_15743_43084# 0.464206f
C13383 a_5691_45260# a_n2661_43370# 0.015295f
C13384 a_8191_45002# a_n2293_42834# 0.084957f
C13385 a_n1151_42308# a_n1079_45724# 0.012662f
C13386 a_11599_46634# a_12839_46116# 0.042002f
C13387 a_15227_44166# a_19692_46634# 0.116169f
C13388 a_19333_46634# a_19466_46812# 0.167526f
C13389 a_584_46384# a_n357_42282# 0.107436f
C13390 a_11309_47204# a_6945_45028# 0.010402f
C13391 a_n743_46660# a_5937_45572# 0.02494f
C13392 a_5807_45002# a_15682_46116# 0.062679f
C13393 a_13661_43548# a_2324_44458# 0.307974f
C13394 a_n4064_37440# VDD 1.66017f
C13395 VDAC_N C1_N_btm 1.7375f
C13396 a_3422_30871# a_n3420_39072# 0.096346f
C13397 a_19721_31679# C2_N_btm 0.040789f
C13398 a_n357_42282# a_15095_43370# 0.034944f
C13399 a_5147_45002# a_5244_44056# 0.122327f
C13400 a_5883_43914# a_8975_43940# 0.50976f
C13401 a_n2267_44484# a_n1809_44850# 0.027606f
C13402 a_n2442_46660# a_n3674_37592# 0.032368f
C13403 a_n2497_47436# a_1423_45028# 1.36987f
C13404 a_13507_46334# a_2437_43646# 0.117533f
C13405 a_16327_47482# a_n2017_45002# 0.209709f
C13406 a_n1991_46122# a_n1736_46482# 0.06121f
C13407 a_n443_46116# a_3232_43370# 0.059286f
C13408 a_4791_45118# a_6171_45002# 0.031317f
C13409 a_n1151_42308# a_7705_45326# 0.042252f
C13410 a_13747_46662# a_16115_45572# 0.029803f
C13411 a_8953_45546# a_9290_44172# 0.373944f
C13412 a_4185_45028# a_2324_44458# 0.015434f
C13413 a_10405_44172# VDD 0.408512f
C13414 a_4361_42308# a_14113_42308# 0.075467f
C13415 a_19479_31679# a_13467_32519# 0.051245f
C13416 a_19386_47436# VDD 0.121241f
C13417 a_18780_47178# START 0.01578f
C13418 a_18479_47436# SINGLE_ENDED 0.040779f
C13419 a_20411_46873# a_3357_43084# 0.157199f
C13420 a_4646_46812# a_n2661_43370# 0.028718f
C13421 a_21588_30879# a_18114_32519# 0.055884f
C13422 a_768_44030# a_5343_44458# 0.066821f
C13423 a_3090_45724# a_7229_43940# 0.054969f
C13424 a_3483_46348# a_8696_44636# 0.06521f
C13425 a_10903_43370# a_11682_45822# 0.071222f
C13426 a_10809_44734# a_10193_42453# 0.02204f
C13427 a_20556_43646# VDD 0.34939f
C13428 COMP_P a_n1794_35082# 2.45644f
C13429 a_n473_42460# a_n327_42558# 0.171361f
C13430 a_13887_32519# C3_N_btm 0.030933f
C13431 a_9313_44734# a_16823_43084# 0.031008f
C13432 a_3905_42865# a_4235_43370# 0.041971f
C13433 a_19551_46910# VDD 0.226848f
C13434 a_n913_45002# a_133_42852# 0.046777f
C13435 a_17715_44484# a_17613_45144# 0.012898f
C13436 a_n2293_45546# a_1667_45002# 0.07132f
C13437 a_1823_45246# a_n699_43396# 0.08003f
C13438 a_n863_45724# a_413_45260# 0.140312f
C13439 a_12465_44636# a_21588_30879# 0.053175f
C13440 a_11453_44696# a_19594_46812# 0.041136f
C13441 a_n443_46116# a_4651_46660# 0.060179f
C13442 a_n237_47217# a_8667_46634# 0.171086f
C13443 a_n3674_37592# a_n3420_37440# 0.073321f
C13444 a_22400_42852# a_22527_39145# 0.228292f
C13445 a_n784_42308# a_n4064_37440# 0.014901f
C13446 a_n97_42460# a_15743_43084# 0.205305f
C13447 a_n4318_40392# a_n3674_38680# 0.023225f
C13448 a_9290_44172# a_9028_43914# 0.169653f
C13449 a_5147_45002# a_5111_44636# 0.562127f
C13450 a_4558_45348# a_4927_45028# 0.123258f
C13451 a_15861_45028# a_17613_45144# 0.016666f
C13452 a_21588_30879# a_13887_32519# 0.056445f
C13453 a_3537_45260# a_3232_43370# 0.530258f
C13454 a_n881_46662# a_n1076_46494# 0.018649f
C13455 a_4883_46098# a_8016_46348# 0.289691f
C13456 a_11599_46634# a_14840_46494# 0.051732f
C13457 a_8667_46634# a_8270_45546# 0.046604f
C13458 a_n2438_43548# a_765_45546# 0.081258f
C13459 a_7227_47204# a_6945_45028# 0.01947f
C13460 a_n3565_39590# VCM 0.097317f
C13461 a_n4064_39616# VIN_P 0.047639f
C13462 a_3754_38470# VDAC_N 0.169096f
C13463 a_n3420_39072# VDD 1.01449f
C13464 a_n2946_37690# a_n2860_37690# 0.011479f
C13465 a_7754_38470# a_5700_37509# 0.971846f
C13466 a_n4064_37440# a_n2302_37690# 0.239588f
C13467 a_8530_39574# a_5088_37509# 0.166912f
C13468 a_4361_42308# a_5534_30871# 0.049795f
C13469 a_1423_45028# a_6109_44484# 0.018788f
C13470 a_3232_43370# a_11541_44484# 0.050289f
C13471 a_13059_46348# a_14275_46494# 0.036863f
C13472 a_n1853_46287# a_n901_46420# 0.049679f
C13473 a_n1991_46122# a_n1641_46494# 0.219633f
C13474 a_n2157_46122# a_n1076_46494# 0.102355f
C13475 a_n743_46660# a_n443_42852# 0.378464f
C13476 a_n1741_47186# a_2437_43646# 4.86702f
C13477 a_12861_44030# a_15861_45028# 0.015193f
C13478 a_20980_44850# VDD 0.132317f
C13479 a_3537_45260# a_4905_42826# 0.339989f
C13480 a_6298_44484# a_7281_43914# 0.010383f
C13481 a_5343_44458# a_7845_44172# 0.103601f
C13482 a_19778_44110# a_15493_43396# 0.015561f
C13483 a_5883_43914# a_5495_43940# 0.09813f
C13484 a_n2833_47464# VDD 0.461379f
C13485 a_22959_46124# a_20692_30879# 0.155635f
C13486 a_15227_44166# a_18175_45572# 0.018929f
C13487 a_5204_45822# a_5263_45724# 0.109078f
C13488 a_n746_45260# a_n23_44458# 0.046452f
C13489 a_3877_44458# a_4558_45348# 0.028316f
C13490 a_12741_44636# a_11823_42460# 0.031865f
C13491 a_6969_46634# VDD 0.154507f
C13492 a_1414_42308# a_1443_43940# 0.018064f
C13493 a_20193_45348# a_13467_32519# 0.016015f
C13494 a_10405_44172# a_10729_43914# 0.083277f
C13495 a_n2293_42834# a_7765_42852# 0.010796f
C13496 a_6945_45028# a_6171_45002# 0.032875f
C13497 a_8049_45260# a_22959_45572# 0.176374f
C13498 a_3090_45724# a_15004_44636# 0.010872f
C13499 a_2711_45572# a_10907_45822# 0.016608f
C13500 a_11415_45002# a_16922_45042# 0.012903f
C13501 a_768_44030# a_453_43940# 0.110708f
C13502 a_3483_46348# a_5009_45028# 0.029292f
C13503 a_12861_44030# a_20623_43914# 0.033132f
C13504 a_n2288_47178# a_n2293_46634# 0.011283f
C13505 a_n1741_47186# a_n2661_46634# 0.22396f
C13506 SMPL_ON_P a_n2956_39768# 0.039986f
C13507 a_4915_47217# a_9804_47204# 0.072476f
C13508 a_n3674_38680# a_n4209_38502# 0.04481f
C13509 a_14113_42308# a_15890_42674# 0.022182f
C13510 a_15486_42560# a_15803_42450# 0.102355f
C13511 a_n3674_39768# a_n4318_38680# 0.024755f
C13512 a_4093_43548# a_4235_43370# 0.515101f
C13513 a_3422_30871# a_5342_30871# 0.026613f
C13514 a_458_43396# a_n1557_42282# 0.027865f
C13515 a_n97_42460# a_3539_42460# 0.021726f
C13516 a_n913_45002# a_5742_30871# 0.028271f
C13517 a_375_42282# a_564_42282# 0.022891f
C13518 a_n2293_46098# a_5663_43940# 0.142661f
C13519 a_8270_45546# a_9165_43940# 0.063297f
C13520 a_n1925_42282# a_n2661_43922# 0.028186f
C13521 a_10180_45724# a_n2661_43370# 0.038795f
C13522 a_n237_47217# a_5204_45822# 0.019965f
C13523 a_11453_44696# a_16388_46812# 0.019353f
C13524 a_10227_46804# a_21363_46634# 0.273017f
C13525 a_13507_46334# a_765_45546# 0.045587f
C13526 a_18597_46090# a_20411_46873# 0.070431f
C13527 a_768_44030# a_3090_45724# 0.115303f
C13528 a_n1925_46634# a_6755_46942# 0.12389f
C13529 a_15486_42560# VDD 0.275297f
C13530 a_22485_38105# CAL_P 0.026856f
C13531 a_19479_31679# RST_Z 0.049574f
C13532 a_2437_43646# SINGLE_ENDED 0.117817f
C13533 a_4190_30871# a_4361_42308# 0.06171f
C13534 a_3357_43084# VDD 1.66202f
C13535 a_5205_44484# a_5518_44484# 0.135771f
C13536 a_3232_43370# a_8701_44490# 0.062297f
C13537 a_526_44458# a_n97_42460# 0.277959f
C13538 a_n2017_45002# a_n356_44636# 0.036195f
C13539 SMPL_ON_P a_n4318_37592# 0.040097f
C13540 a_n1925_46634# a_8049_45260# 0.088663f
C13541 a_5257_43370# a_2324_44458# 0.067403f
C13542 C10_N_btm VDD 2.40001f
C13543 C3_P_btm VREF_GND 0.67174f
C13544 C4_P_btm VCM 0.716447f
C13545 C2_P_btm VREF 0.987884f
C13546 C0_P_btm VIN_P 0.529671f
C13547 a_3539_42460# a_3823_42558# 0.07742f
C13548 a_8975_43940# a_11541_44484# 0.028558f
C13549 a_n443_42852# a_4361_42308# 0.016253f
C13550 a_n863_45724# a_n13_43084# 0.041588f
C13551 a_15004_44636# a_14815_43914# 0.078606f
C13552 a_11827_44484# a_20512_43084# 0.030456f
C13553 a_n2956_39304# a_n2956_38680# 0.163045f
C13554 a_n743_46660# a_2437_43646# 0.031693f
C13555 a_n1613_43370# a_3232_43370# 0.091534f
C13556 a_8199_44636# a_10586_45546# 0.057648f
C13557 a_3065_45002# a_3935_42891# 0.01149f
C13558 a_n1549_44318# a_n1441_43940# 0.057222f
C13559 a_n913_45002# a_10922_42852# 0.01889f
C13560 a_n1059_45260# a_10341_42308# 0.032786f
C13561 a_n2293_46634# VDD 1.52629f
C13562 a_n2956_39768# CLK_DATA 0.015401f
C13563 a_526_44458# a_3823_42558# 0.183187f
C13564 a_18597_46090# a_3422_30871# 0.030159f
C13565 a_4646_46812# a_5883_43914# 0.019308f
C13566 a_167_45260# a_n37_45144# 0.277898f
C13567 a_n2293_46098# a_3232_43370# 0.054403f
C13568 a_4915_47217# a_6545_47178# 0.033555f
C13569 a_14097_32519# a_4958_30871# 0.030871f
C13570 a_5342_30871# VDD 0.496295f
C13571 a_9625_46129# VDD 0.996485f
C13572 a_526_44458# a_742_44458# 0.54618f
C13573 a_13259_45724# a_16922_45042# 0.401687f
C13574 a_10809_44734# a_10057_43914# 0.060542f
C13575 a_7499_43078# a_5111_44636# 0.753731f
C13576 a_21588_30879# a_14401_32519# 0.058775f
C13577 a_n2661_46634# a_n743_46660# 0.037388f
C13578 a_n2293_46634# a_n2312_38680# 0.131017f
C13579 a_n1741_47186# a_765_45546# 0.536367f
C13580 a_n1613_43370# a_4651_46660# 0.686447f
C13581 a_n881_46662# a_4646_46812# 0.024758f
C13582 a_n473_42460# VDD 0.27195f
C13583 a_n3565_39590# a_n4064_38528# 0.031177f
C13584 a_n4315_30879# a_n4209_38216# 0.053149f
C13585 a_1273_38525# a_1169_39043# 0.010455f
C13586 a_5742_30871# VDAC_P 0.030334f
C13587 a_n3420_39616# a_n3420_38528# 0.049464f
C13588 a_n4064_39616# a_n3565_38502# 0.02802f
C13589 a_n3565_39304# a_n2302_39072# 0.066757f
C13590 a_n3690_39392# a_n4064_39072# 0.085872f
C13591 a_n3420_39072# a_n2946_39072# 0.238708f
C13592 a_10341_43396# a_18783_43370# 0.010939f
C13593 a_n1059_45260# a_18494_42460# 0.187733f
C13594 a_7705_45326# a_n2293_42834# 0.071732f
C13595 a_n746_45260# a_n356_45724# 0.030083f
C13596 a_584_46384# a_310_45028# 0.024195f
C13597 a_n1151_42308# a_n2293_45546# 0.01733f
C13598 a_15227_44166# a_19466_46812# 0.310201f
C13599 a_2443_46660# a_167_45260# 0.012819f
C13600 a_n743_46660# a_8199_44636# 0.046048f
C13601 a_5807_45002# a_2324_44458# 0.232399f
C13602 a_n2946_37690# VDD 0.38221f
C13603 a_n2002_35448# a_n1550_35448# 0.150805f
C13604 VDAC_N C0_N_btm 0.901121f
C13605 VDAC_P C0_dummy_P_btm 0.88451f
C13606 a_16237_45028# VDD 0.248452f
C13607 a_9290_44172# a_5534_30871# 0.472376f
C13608 a_5147_45002# a_3905_42865# 0.048808f
C13609 a_10903_43370# a_12895_43230# 0.011631f
C13610 a_13259_45724# a_15743_43084# 0.021493f
C13611 a_10157_44484# a_10334_44484# 0.159555f
C13612 a_n2267_44484# a_n2012_44484# 0.05936f
C13613 a_n2129_44697# a_n1809_44850# 0.026556f
C13614 a_2063_45854# a_10951_45334# 0.016425f
C13615 a_21177_47436# a_2437_43646# 0.014824f
C13616 a_n1853_46287# a_n1736_46482# 0.170096f
C13617 a_4791_45118# a_3232_43370# 0.268929f
C13618 a_n1151_42308# a_6709_45028# 0.286957f
C13619 a_13747_46662# a_16333_45814# 0.018523f
C13620 a_9625_46129# a_9823_46155# 0.321686f
C13621 a_5342_30871# a_n784_42308# 0.049079f
C13622 a_743_42282# a_15803_42450# 0.037845f
C13623 a_9672_43914# VDD 0.150499f
C13624 a_5891_43370# a_8333_44056# 0.070354f
C13625 a_14539_43914# a_15493_43940# 0.625897f
C13626 a_n2293_42834# a_2982_43646# 0.019738f
C13627 a_18597_46090# VDD 0.930122f
C13628 a_18479_47436# START 0.313639f
C13629 w_10694_33990# a_3422_30871# 3.14233f
C13630 a_20107_46660# a_3357_43084# 0.025828f
C13631 a_3877_44458# a_n2661_43370# 0.038641f
C13632 a_n2833_47464# a_n2497_47436# 0.217831f
C13633 a_743_42282# VDD 0.597869f
C13634 a_n473_42460# a_n784_42308# 0.020033f
C13635 a_n4318_37592# a_n1794_35082# 0.847279f
C13636 a_3905_42865# a_4093_43548# 0.032751f
C13637 a_19123_46287# VDD 0.336379f
C13638 a_n1059_45260# a_133_42852# 0.045134f
C13639 en_comp a_n2293_42282# 0.026f
C13640 a_11967_42832# a_14579_43548# 0.060711f
C13641 a_12741_44636# a_14539_43914# 0.09527f
C13642 a_3090_45724# a_17517_44484# 0.020082f
C13643 a_1138_42852# a_n699_43396# 0.024181f
C13644 a_18189_46348# a_16922_45042# 0.015824f
C13645 a_13249_42308# a_8696_44636# 0.021669f
C13646 a_n2293_45546# a_327_44734# 0.027309f
C13647 a_10903_43370# a_11827_44484# 0.021644f
C13648 a_4791_45118# a_4905_42826# 0.516502f
C13649 a_167_45260# a_949_44458# 0.021626f
C13650 a_n863_45724# a_n37_45144# 0.056531f
C13651 a_n881_46662# a_9804_47204# 0.061323f
C13652 a_11453_44696# a_19321_45002# 0.023175f
C13653 a_4791_45118# a_4651_46660# 0.020454f
C13654 a_n443_46116# a_4646_46812# 0.077958f
C13655 a_n971_45724# a_8492_46660# 0.016456f
C13656 a_n3674_37592# a_n3690_37440# 0.071822f
C13657 a_22400_42852# a_22589_40055# 0.663766f
C13658 a_8791_43396# a_8685_43396# 0.086218f
C13659 a_2277_45546# VDD 0.209584f
C13660 a_n443_42852# a_5891_43370# 0.175668f
C13661 a_15861_45028# a_17023_45118# 0.076138f
C13662 a_8696_44636# a_17613_45144# 0.09062f
C13663 a_4574_45260# a_4927_45028# 0.047624f
C13664 a_3357_43084# a_1423_45028# 0.02044f
C13665 a_n881_46662# a_n901_46420# 0.053662f
C13666 a_n1613_43370# a_n1076_46494# 0.232314f
C13667 a_11599_46634# a_15015_46420# 0.040858f
C13668 a_10227_46804# a_11133_46155# 0.019137f
C13669 a_6851_47204# a_6945_45028# 0.013916f
C13670 a_2063_45854# a_n1925_42282# 0.025501f
C13671 a_n743_46660# a_765_45546# 0.148721f
C13672 a_n3565_39590# VREF_GND 0.041931f
C13673 a_n4064_37984# EN_VIN_BSTR_P 0.031797f
C13674 a_n3690_39392# VDD 0.363068f
C13675 a_8530_39574# a_4338_37500# 0.093669f
C13676 a_7754_38470# a_5088_37509# 0.394117f
C13677 a_685_42968# a_791_42968# 0.13675f
C13678 a_13467_32519# a_5534_30871# 0.041703f
C13679 a_626_44172# VDD 0.621601f
C13680 a_8199_44636# a_4361_42308# 0.024061f
C13681 a_n863_45724# a_104_43370# 0.046664f
C13682 a_n743_46660# a_509_45822# 0.039863f
C13683 a_13059_46348# a_14493_46090# 0.029059f
C13684 a_n1853_46287# a_n1641_46494# 0.033696f
C13685 a_n1991_46122# a_n1423_46090# 0.175891f
C13686 a_n2157_46122# a_n901_46420# 0.043559f
C13687 a_19692_46634# a_10809_44734# 0.014397f
C13688 a_12861_44030# a_8696_44636# 0.046746f
C13689 a_n4318_39304# a_n4064_39616# 0.059009f
C13690 a_743_42282# a_n784_42308# 0.087438f
C13691 a_3537_45260# a_3080_42308# 0.02683f
C13692 w_10694_33990# VDD 1.82872f
C13693 a_5343_44458# a_7542_44172# 0.014194f
C13694 a_19778_44110# a_19328_44172# 0.064774f
C13695 a_9290_44172# a_n443_42852# 0.483812f
C13696 a_22959_46124# a_20205_31679# 0.012679f
C13697 a_4646_46812# a_3537_45260# 0.361823f
C13698 a_3877_44458# a_4574_45260# 0.010367f
C13699 a_15227_44166# a_16147_45260# 0.282941f
C13700 a_n743_46660# a_16751_45260# 0.028358f
C13701 a_n746_45260# a_n356_44636# 0.418585f
C13702 a_n2293_46634# a_1423_45028# 0.025918f
C13703 a_1467_44172# a_1443_43940# 0.011516f
C13704 a_n2293_43922# a_3626_43646# 0.03147f
C13705 a_n2293_42834# a_7871_42858# 0.027f
C13706 a_6755_46942# VDD 1.05713f
C13707 a_8049_45260# a_19963_31679# 0.2062f
C13708 a_1823_45246# a_n2293_42834# 0.031316f
C13709 a_5257_43370# a_5708_44484# 0.056224f
C13710 a_768_44030# a_1414_42308# 0.072003f
C13711 a_13259_45724# a_17668_45572# 0.050071f
C13712 a_2324_44458# a_13017_45260# 0.021259f
C13713 a_12861_44030# a_20365_43914# 0.044371f
C13714 a_10227_46804# a_13507_46334# 0.120657f
C13715 a_n2497_47436# a_n2293_46634# 0.174929f
C13716 a_4915_47217# a_8128_46384# 0.070866f
C13717 a_6545_47178# a_n881_46662# 0.020203f
C13718 a_6491_46660# a_n1613_43370# 0.071408f
C13719 a_15051_42282# a_15803_42450# 0.043619f
C13720 a_15486_42560# a_15764_42576# 0.118759f
C13721 a_14113_42308# a_15959_42545# 0.036113f
C13722 a_n4318_39768# a_n4318_38680# 0.02372f
C13723 a_n3674_39768# a_n3674_39304# 0.037712f
C13724 a_5111_44636# a_5932_42308# 0.021257f
C13725 a_458_43396# a_766_43646# 0.017351f
C13726 a_8049_45260# VDD 1.89366f
C13727 a_n97_42460# a_3626_43646# 0.394673f
C13728 a_n863_45724# a_949_44458# 0.034335f
C13729 a_3357_43084# a_22591_45572# 0.181818f
C13730 a_19479_31679# a_19963_31679# 0.104687f
C13731 a_n2293_46098# a_5495_43940# 0.096987f
C13732 a_13661_43548# a_13667_43396# 0.168674f
C13733 a_1138_42852# a_1467_44172# 0.034446f
C13734 a_n1925_42282# a_n2661_42834# 0.029302f
C13735 a_13259_45724# a_17970_44736# 0.011308f
C13736 a_526_44458# a_n2661_43922# 0.154533f
C13737 a_n237_47217# a_5164_46348# 0.081549f
C13738 a_n443_46116# a_n901_46420# 0.367344f
C13739 a_11453_44696# a_13059_46348# 0.039573f
C13740 a_10227_46804# a_20623_46660# 0.156341f
C13741 a_13507_46334# a_17339_46660# 0.05814f
C13742 a_12549_44172# a_3090_45724# 0.082348f
C13743 a_18479_47436# a_20273_46660# 0.018124f
C13744 a_15051_42282# VDD 0.461307f
C13745 a_n4064_39072# a_n3420_37440# 0.051893f
C13746 a_n3420_39072# a_n4064_37440# 0.047151f
C13747 a_n2302_37984# a_n2216_37984# 0.011479f
C13748 a_4190_30871# a_13467_32519# 0.032722f
C13749 a_2437_43646# START 0.12936f
C13750 a_19479_31679# VDD 0.583964f
C13751 a_5205_44484# a_5343_44458# 0.129692f
C13752 a_n443_42852# a_10807_43548# 0.173997f
C13753 a_3357_43084# a_6109_44484# 0.016236f
C13754 a_3232_43370# a_8103_44636# 0.013825f
C13755 a_20202_43084# a_15743_43084# 0.021267f
C13756 a_10249_46116# a_10355_46116# 0.182836f
C13757 C9_N_btm VDD 0.345685f
C13758 C4_P_btm VREF_GND 0.671882f
C13759 C5_P_btm VCM 0.719982f
C13760 C3_P_btm VREF 0.984942f
C13761 C1_P_btm VIN_P 0.39234f
C13762 a_3422_30871# a_n3420_37440# 0.0344f
C13763 a_3539_42460# a_3318_42354# 0.161793f
C13764 a_3626_43646# a_3823_42558# 0.017529f
C13765 a_2982_43646# a_5379_42460# 0.068435f
C13766 a_n357_42282# a_n1853_43023# 0.04297f
C13767 a_n2956_38216# a_n4318_38680# 0.023204f
C13768 a_20193_45348# a_3422_30871# 0.042753f
C13769 a_n2840_46090# a_n2840_45546# 0.025171f
C13770 a_11453_44696# a_13556_45296# 0.027553f
C13771 a_15037_43940# VDD 0.190221f
C13772 a_n1331_43914# a_n1441_43940# 0.097745f
C13773 a_n2017_45002# a_10341_42308# 0.049998f
C13774 a_n913_45002# a_10991_42826# 0.029878f
C13775 a_n2442_46660# VDD 0.693209f
C13776 a_12549_44172# a_14815_43914# 0.026324f
C13777 a_13259_45724# a_13163_45724# 0.166368f
C13778 a_167_45260# a_n143_45144# 0.03701f
C13779 a_1823_45246# a_413_45260# 0.043122f
C13780 a_4915_47217# a_6151_47436# 0.783303f
C13781 a_n1741_47186# a_10227_46804# 0.020904f
C13782 a_1606_42308# a_5742_30871# 3.46204f
C13783 a_5534_30871# RST_Z 0.031803f
C13784 a_15279_43071# VDD 0.189193f
C13785 a_8953_45546# VDD 1.32809f
C13786 a_10193_42453# a_13258_32519# 0.061618f
C13787 a_n2956_38216# a_n4209_38216# 0.232905f
C13788 a_9313_44734# a_12089_42308# 0.011899f
C13789 a_17478_45572# a_17668_45572# 0.045837f
C13790 a_3090_45724# a_7542_44172# 0.137368f
C13791 a_8199_44636# a_5891_43370# 0.399007f
C13792 a_n2442_46660# a_n2312_38680# 0.068683f
C13793 a_n1613_43370# a_4646_46812# 1.38979f
C13794 a_n881_46662# a_3877_44458# 0.142507f
C13795 a_n2293_46634# a_n2104_46634# 0.042499f
C13796 a_n961_42308# VDD 0.24416f
C13797 a_14097_32519# VREF_GND 0.047244f
C13798 a_n3565_39304# a_n4064_39072# 0.344587f
C13799 a_10341_43396# a_18525_43370# 0.015853f
C13800 a_1568_43370# a_1847_42826# 0.153113f
C13801 a_n1059_45260# a_18184_42460# 0.52106f
C13802 a_13059_46348# a_9145_43396# 0.028786f
C13803 a_n863_45724# a_175_44278# 0.113317f
C13804 a_n755_45592# a_n1761_44111# 0.015303f
C13805 a_626_44172# a_1423_45028# 0.014461f
C13806 a_5111_44636# a_n2661_43370# 0.075649f
C13807 a_n971_45724# a_n356_45724# 0.030873f
C13808 a_584_46384# a_n1099_45572# 0.021537f
C13809 a_10227_46804# a_10586_45546# 0.306536f
C13810 a_15227_44166# a_19333_46634# 0.065741f
C13811 a_n3420_37440# VDD 2.26579f
C13812 VDAC_N C0_dummy_N_btm 0.885361f
C13813 VDAC_P C0_P_btm 0.901219f
C13814 CAL_P EN_VIN_BSTR_N 0.040136f
C13815 a_5342_30871# a_15567_42826# 0.024331f
C13816 a_20193_45348# VDD 0.793111f
C13817 a_10903_43370# a_13113_42826# 0.011891f
C13818 a_n2129_44697# a_n2012_44484# 0.172424f
C13819 w_1575_34786# a_n4064_39072# 0.017447f
C13820 a_13747_46662# a_15765_45572# 0.5661f
C13821 a_9625_46129# a_9569_46155# 0.204034f
C13822 a_13059_46348# a_14180_46482# 0.025233f
C13823 a_n2497_47436# a_626_44172# 0.249352f
C13824 a_3090_45724# a_n2661_45546# 0.561435f
C13825 a_2063_45854# a_10775_45002# 0.012226f
C13826 a_n1151_42308# a_7229_43940# 0.036511f
C13827 a_n2157_46122# a_n1736_46482# 0.086708f
C13828 a_3483_46348# a_2324_44458# 0.668551f
C13829 a_8199_44636# a_9290_44172# 0.516297f
C13830 a_743_42282# a_15764_42576# 0.054445f
C13831 a_9028_43914# VDD 0.17194f
C13832 a_18780_47178# VDD 0.245515f
C13833 w_1575_34786# a_3422_30871# 2.62797f
C13834 a_768_44030# a_n699_43396# 1.37533f
C13835 a_16327_47482# a_9313_44734# 0.169217f
C13836 a_10903_43370# a_10907_45822# 0.199567f
C13837 a_5066_45546# a_5263_45724# 0.022243f
C13838 a_20301_43646# VDD 0.296691f
C13839 a_5342_30871# a_n4064_37440# 0.028573f
C13840 a_4190_30871# RST_Z 0.087843f
C13841 a_22165_42308# a_17303_42282# 0.095988f
C13842 a_n1736_42282# a_n1794_35082# 0.071684f
C13843 COMP_P a_n3674_37592# 0.054748f
C13844 a_n961_42308# a_n784_42308# 0.154417f
C13845 a_10807_43548# a_11257_43940# 0.013221f
C13846 a_18285_46348# VDD 0.259614f
C13847 a_12741_44636# a_16112_44458# 0.019518f
C13848 a_13661_43548# a_15493_43396# 0.491785f
C13849 a_17715_44484# a_16922_45042# 0.039816f
C13850 a_n2293_45546# a_413_45260# 0.066602f
C13851 a_n863_45724# a_n143_45144# 0.033306f
C13852 a_10227_46804# a_n743_46660# 0.134234f
C13853 a_n881_46662# a_8128_46384# 0.206292f
C13854 a_21811_47423# a_20916_46384# 0.109084f
C13855 a_4791_45118# a_4646_46812# 0.485113f
C13856 a_n443_46116# a_3877_44458# 0.06318f
C13857 a_n3674_37592# a_n3565_37414# 0.129086f
C13858 a_19511_42282# a_21125_42558# 0.01129f
C13859 a_n784_42308# a_n3420_37440# 0.140549f
C13860 a_19319_43548# a_4190_30871# 0.188868f
C13861 a_1609_45822# VDD 0.270106f
C13862 a_n2956_37592# a_n3565_39590# 0.023811f
C13863 a_8147_43396# a_8685_43396# 0.077232f
C13864 a_4558_45348# a_5147_45002# 0.09356f
C13865 a_3065_45002# a_3232_43370# 0.049451f
C13866 a_8696_44636# a_17023_45118# 0.064781f
C13867 a_15861_45028# a_16922_45042# 0.259169f
C13868 a_22612_30879# a_13678_32519# 0.060546f
C13869 a_3537_45260# a_4927_45028# 0.216859f
C13870 a_n1613_43370# a_n901_46420# 0.406381f
C13871 a_11599_46634# a_14275_46494# 0.029786f
C13872 a_n237_47217# a_5066_45546# 1.48406f
C13873 a_12861_44030# a_15682_46116# 0.030474f
C13874 a_584_46384# a_n1925_42282# 0.194054f
C13875 a_2063_45854# a_526_44458# 0.039908f
C13876 a_n4064_38528# C5_P_btm 0.042017f
C13877 a_n3420_39616# VIN_P 0.04023f
C13878 a_n3565_39590# VREF 0.417978f
C13879 a_n4209_39590# VCM 0.179761f
C13880 a_n3565_39304# VDD 0.898174f
C13881 a_8530_39574# a_3726_37500# 1.35509f
C13882 a_7754_38470# a_4338_37500# 0.208561f
C13883 a_3754_38470# a_5700_37509# 0.124176f
C13884 a_n2946_37690# a_n4064_37440# 0.053228f
C13885 a_n863_45724# a_n97_42460# 0.581863f
C13886 a_13259_45724# a_3626_43646# 0.037016f
C13887 a_11823_42460# a_11341_43940# 0.087329f
C13888 a_8270_45546# a_5066_45546# 0.189476f
C13889 a_13059_46348# a_13925_46122# 0.056739f
C13890 a_n1853_46287# a_n1423_46090# 0.043126f
C13891 a_n2157_46122# a_n1641_46494# 0.105995f
C13892 a_5807_45002# a_6511_45714# 0.012932f
C13893 a_n2109_47186# a_2437_43646# 0.027184f
C13894 a_3626_43646# a_18057_42282# 0.01061f
C13895 a_3537_45260# a_4699_43561# 0.024682f
C13896 w_1575_34786# VDD 1.60056f
C13897 a_n2312_38680# a_n3565_39304# 0.418567f
C13898 a_10809_44734# a_20205_31679# 0.039075f
C13899 a_3877_44458# a_3537_45260# 0.12249f
C13900 a_2107_46812# a_9482_43914# 0.109711f
C13901 a_5342_30871# a_n3420_39072# 0.062032f
C13902 a_1467_44172# a_1241_43940# 0.011879f
C13903 a_1115_44172# a_1443_43940# 0.096132f
C13904 a_10249_46116# VDD 1.03004f
C13905 a_12861_44030# a_20269_44172# 0.047709f
C13906 a_768_44030# a_1467_44172# 0.022755f
C13907 a_8953_45546# a_1423_45028# 0.021907f
C13908 a_1138_42852# a_n2293_42834# 0.015752f
C13909 a_8049_45260# a_22591_45572# 0.036446f
C13910 a_n2497_47436# a_n2442_46660# 0.045496f
C13911 a_n2109_47186# a_n2661_46634# 0.038259f
C13912 a_n1151_42308# a_768_44030# 0.019901f
C13913 a_6151_47436# a_n881_46662# 1.58776f
C13914 a_18479_47436# a_20894_47436# 0.032517f
C13915 a_15051_42282# a_15764_42576# 0.042737f
C13916 a_14113_42308# a_15803_42450# 0.289859f
C13917 a_n4318_39768# a_n3674_39304# 0.024426f
C13918 a_n97_42460# a_3540_43646# 0.027089f
C13919 a_3537_45260# a_6761_42308# 0.057884f
C13920 a_n2661_42282# a_5649_42852# 0.052118f
C13921 a_3422_30871# a_5534_30871# 0.023427f
C13922 a_n863_45724# a_742_44458# 0.629795f
C13923 a_19479_31679# a_22591_45572# 0.011797f
C13924 a_9049_44484# a_n2661_43370# 0.030026f
C13925 a_10227_46804# a_4361_42308# 0.073929f
C13926 a_n2293_46098# a_5013_44260# 0.040459f
C13927 a_526_44458# a_n2661_42834# 0.06021f
C13928 a_13259_45724# a_17767_44458# 0.026768f
C13929 a_1138_42852# a_1115_44172# 0.012127f
C13930 a_768_44030# a_14084_46812# 0.013767f
C13931 a_n237_47217# a_5068_46348# 0.033474f
C13932 a_10227_46804# a_20841_46902# 0.164019f
C13933 a_2063_45854# a_2521_46116# 0.011365f
C13934 a_2107_46812# a_7715_46873# 0.032178f
C13935 a_18479_47436# a_20411_46873# 0.192791f
C13936 a_14113_42308# VDD 0.365578f
C13937 a_2112_39137# VDAC_Ni 0.018095f
C13938 a_743_42282# a_20556_43646# 0.028541f
C13939 a_4190_30871# a_19095_43396# 0.046015f
C13940 a_22223_45572# VDD 0.287831f
C13941 a_2437_43646# RST_Z 0.082469f
C13942 a_7229_43940# a_4223_44672# 0.014299f
C13943 a_9482_43914# a_n2661_44458# 0.017706f
C13944 a_n357_42282# a_19862_44208# 0.138067f
C13945 a_n2293_45010# a_n356_44636# 0.031375f
C13946 a_3232_43370# a_6298_44484# 0.256727f
C13947 a_5111_44636# a_5883_43914# 0.281106f
C13948 SMPL_ON_P a_n3674_38216# 0.044338f
C13949 a_4646_46812# a_6945_45028# 0.090679f
C13950 a_10249_46116# a_9823_46155# 0.082191f
C13951 a_n743_46660# a_8034_45724# 0.021079f
C13952 a_16327_47482# a_2711_45572# 0.101699f
C13953 C8_N_btm VDD 0.19922f
C13954 C5_P_btm VREF_GND 0.676559f
C13955 C6_P_btm VCM 0.877162f
C13956 C4_P_btm VREF 0.98728f
C13957 C2_P_btm VIN_P 0.502408f
C13958 a_11823_42460# a_10341_43396# 0.088285f
C13959 a_n2956_38216# a_n3674_39304# 0.023342f
C13960 a_13720_44458# a_14112_44734# 0.016359f
C13961 a_n2312_39304# a_n3565_39590# 0.491833f
C13962 a_20202_43084# a_21195_42852# 0.018373f
C13963 a_n1925_46634# a_2437_43646# 0.02753f
C13964 a_n2293_46634# a_3357_43084# 0.963711f
C13965 a_11453_44696# a_9482_43914# 0.042575f
C13966 a_12465_44636# a_14537_43396# 0.031033f
C13967 a_13565_43940# VDD 0.175245f
C13968 a_10903_43370# a_13070_42354# 0.04369f
C13969 a_2382_45260# a_3935_42891# 0.061675f
C13970 a_n1899_43946# a_n1441_43940# 0.03441f
C13971 a_11967_42832# a_15493_43396# 0.02628f
C13972 a_n913_45002# a_10796_42968# 0.545674f
C13973 a_n2472_46634# VDD 0.287589f
C13974 a_1138_42852# a_413_45260# 0.026098f
C13975 a_4791_45118# a_5013_44260# 0.02062f
C13976 a_768_44030# a_13857_44734# 0.011246f
C13977 a_10586_45546# a_11682_45822# 0.014019f
C13978 a_n2293_46098# a_4927_45028# 0.015237f
C13979 a_4915_47217# a_5815_47464# 0.064955f
C13980 a_4791_45118# a_6545_47178# 0.112353f
C13981 a_5534_30871# VDD 0.513761f
C13982 a_9313_44734# a_12379_42858# 0.05039f
C13983 a_3422_30871# a_4190_30871# 12.909901f
C13984 en_comp a_22400_42852# 0.721871f
C13985 a_5937_45572# VDD 2.20055f
C13986 a_n2810_45572# a_n3565_38216# 0.104999f
C13987 a_15861_45028# a_17668_45572# 0.065471f
C13988 a_2711_45572# a_14537_43396# 0.249285f
C13989 a_3090_45724# a_7281_43914# 0.170855f
C13990 a_8199_44636# a_8375_44464# 0.043989f
C13991 a_n2109_47186# a_765_45546# 0.126431f
C13992 a_n2472_46634# a_n2312_38680# 0.039578f
C13993 a_n2661_46634# a_n1925_46634# 4.75867f
C13994 a_n1613_43370# a_3877_44458# 1.43013f
C13995 a_n3565_39590# a_n3420_38528# 0.031237f
C13996 COMP_P RST_Z 0.03403f
C13997 a_1666_39587# a_1666_39043# 1.95282f
C13998 a_n4334_39392# a_n4064_39072# 0.410653f
C13999 a_n4209_39304# a_n2302_39072# 0.407162f
C14000 a_n4209_39590# a_n4064_38528# 0.032071f
C14001 a_1606_42308# C0_P_btm 0.029189f
C14002 a_n3420_39616# a_n3565_38502# 0.028014f
C14003 a_n4064_39616# a_n4209_38502# 0.02801f
C14004 a_n3565_39304# a_n2946_39072# 0.410957f
C14005 a_n3690_39392# a_n3420_39072# 0.414961f
C14006 a_n1329_42308# VDD 0.237697f
C14007 a_10341_43396# a_18429_43548# 0.012565f
C14008 a_15095_43370# a_15743_43084# 0.022008f
C14009 a_n2017_45002# a_18184_42460# 0.205351f
C14010 a_15227_44166# a_15781_43660# 0.016739f
C14011 a_7229_43940# a_n2293_42834# 0.148023f
C14012 a_11823_42460# a_n2293_43922# 0.494696f
C14013 a_5147_45002# a_n2661_43370# 0.034793f
C14014 a_1799_45572# a_167_45260# 0.061186f
C14015 a_3877_44458# a_n2293_46098# 0.030683f
C14016 a_n971_45724# a_3503_45724# 0.011412f
C14017 a_9804_47204# a_6945_45028# 0.028722f
C14018 a_n743_46660# a_8016_46348# 0.155955f
C14019 a_n3690_37440# VDD 0.363068f
C14020 VDAC_P C1_P_btm 1.74268f
C14021 CAL_P a_10890_34112# 0.041859f
C14022 a_11691_44458# VDD 3.25709f
C14023 a_n357_42282# a_14579_43548# 0.049501f
C14024 a_10903_43370# a_12545_42858# 0.026404f
C14025 a_n2433_44484# a_n2012_44484# 0.093133f
C14026 a_11823_42460# a_n97_42460# 0.324041f
C14027 a_10227_46804# a_15890_42674# 0.159412f
C14028 a_n2956_39768# a_n3674_37592# 0.031375f
C14029 a_13747_46662# a_15903_45785# 0.022255f
C14030 a_8953_45546# a_9569_46155# 0.014447f
C14031 a_13059_46348# a_12638_46436# 0.053952f
C14032 a_4791_45118# a_4927_45028# 0.03353f
C14033 a_18597_46090# a_3357_43084# 0.160577f
C14034 a_5257_43370# a_6472_45840# 0.012073f
C14035 a_n1151_42308# a_7276_45260# 0.062423f
C14036 a_8199_44636# a_10355_46116# 0.176325f
C14037 a_n1925_46634# a_8192_45572# 0.03394f
C14038 a_5534_30871# a_n784_42308# 9.92256f
C14039 a_743_42282# a_15486_42560# 0.010882f
C14040 a_8333_44056# VDD 0.124235f
C14041 a_14539_43914# a_11341_43940# 0.077754f
C14042 a_10227_46804# START 0.088203f
C14043 a_18479_47436# VDD 1.47669f
C14044 a_526_44458# a_3775_45552# 0.015665f
C14045 a_15015_46420# a_15143_45578# 0.011172f
C14046 a_14976_45028# a_6171_45002# 0.024858f
C14047 a_10227_46804# a_5891_43370# 0.2393f
C14048 a_2324_44458# a_13249_42308# 0.072143f
C14049 a_768_44030# a_4223_44672# 0.136643f
C14050 a_4190_30871# VDD 1.36846f
C14051 a_n4318_37592# a_n3674_37592# 3.06402f
C14052 a_n3674_38216# a_n1794_35082# 0.333493f
C14053 a_10807_43548# a_11173_43940# 0.013678f
C14054 a_17829_46910# VDD 0.37446f
C14055 a_20692_30879# a_13258_32519# 0.055049f
C14056 a_n2293_45546# a_n37_45144# 0.042299f
C14057 a_n863_45724# a_n467_45028# 0.037721f
C14058 a_n1151_42308# a_5167_46660# 0.011285f
C14059 a_4883_46098# a_20916_46384# 0.471396f
C14060 a_11453_44696# a_13747_46662# 0.046437f
C14061 a_4791_45118# a_3877_44458# 0.024145f
C14062 a_4700_47436# a_4646_46812# 0.010115f
C14063 a_n237_47217# a_7577_46660# 0.032223f
C14064 a_n971_45724# a_7927_46660# 0.035261f
C14065 a_13258_32519# a_21613_42308# 0.060546f
C14066 a_n3674_37592# a_n4334_37440# 0.050036f
C14067 a_22400_42852# a_22537_40625# 0.93502f
C14068 a_n2810_45028# a_n3565_39590# 0.021277f
C14069 a_2982_43646# a_10341_43396# 0.029008f
C14070 a_n443_42852# VDD 3.69394f
C14071 a_2813_43396# a_3457_43396# 0.026697f
C14072 a_16327_47482# a_18817_42826# 0.215236f
C14073 a_8696_44636# a_16922_45042# 0.10244f
C14074 a_9049_44484# a_5883_43914# 0.025986f
C14075 a_21588_30879# a_13678_32519# 0.056847f
C14076 a_3537_45260# a_5111_44636# 1.36722f
C14077 a_n863_45724# a_n2661_43922# 0.115404f
C14078 a_n1925_46634# a_765_45546# 0.029508f
C14079 a_n1613_43370# a_n1641_46494# 0.152421f
C14080 a_11599_46634# a_14493_46090# 0.018622f
C14081 a_10227_46804# a_9290_44172# 0.918064f
C14082 a_7927_46660# a_8023_46660# 0.013793f
C14083 a_12861_44030# a_2324_44458# 0.95556f
C14084 a_6545_47178# a_6945_45028# 0.09952f
C14085 a_584_46384# a_526_44458# 0.458472f
C14086 a_768_44030# a_12741_44636# 0.03898f
C14087 a_6755_46942# a_6969_46634# 0.085936f
C14088 a_n3420_38528# C4_P_btm 0.030945f
C14089 a_7754_40130# CAL_P 0.04831f
C14090 a_n3420_37984# EN_VIN_BSTR_P 0.031831f
C14091 a_n4334_39392# VDD 0.385989f
C14092 VDAC_Ni a_6886_37412# 0.178275f
C14093 a_n4209_39590# VREF_GND 0.083908f
C14094 a_7754_38470# a_3726_37500# 0.124796f
C14095 a_3754_38470# a_5088_37509# 0.632585f
C14096 a_n3420_37440# a_n4064_37440# 8.19012f
C14097 a_743_42282# a_5342_30871# 0.035916f
C14098 a_375_42282# VDD 0.591443f
C14099 a_1307_43914# a_5891_43370# 0.084799f
C14100 a_13059_46348# a_13759_46122# 0.249771f
C14101 a_19333_46634# a_10809_44734# 0.011589f
C14102 a_n2157_46122# a_n1423_46090# 0.053479f
C14103 a_n1853_46287# a_n1991_46122# 0.737461f
C14104 a_19692_46634# a_6945_45028# 0.669658f
C14105 a_5807_45002# a_6472_45840# 0.016039f
C14106 a_n4318_39304# a_n3420_39616# 0.256393f
C14107 a_4190_30871# a_n784_42308# 0.019472f
C14108 a_16922_45042# a_20365_43914# 0.021687f
C14109 a_3065_45002# a_3080_42308# 0.171466f
C14110 a_3537_45260# a_4235_43370# 0.010714f
C14111 a_15433_44458# a_14673_44172# 0.027789f
C14112 a_22223_46124# a_20205_31679# 0.160234f
C14113 a_11415_45002# a_11823_42460# 0.349238f
C14114 a_3877_44458# a_3429_45260# 0.02987f
C14115 a_13507_46334# a_11827_44484# 0.384415f
C14116 a_768_44030# a_n2293_42834# 0.036156f
C14117 a_5204_45822# a_2711_45572# 0.021829f
C14118 a_6655_43762# VDD 0.132357f
C14119 a_n755_45592# a_2351_42308# 0.057532f
C14120 a_10554_47026# VDD 0.205847f
C14121 a_1115_44172# a_1241_43940# 0.143754f
C14122 a_14539_43914# a_10341_43396# 0.041922f
C14123 a_n2293_43922# a_2982_43646# 0.094429f
C14124 a_18579_44172# a_18533_43940# 0.011624f
C14125 a_8568_45546# a_7499_43078# 0.070368f
C14126 a_12861_44030# a_19862_44208# 0.721035f
C14127 a_5937_45572# a_1423_45028# 0.083936f
C14128 a_9290_44172# a_1307_43914# 0.122831f
C14129 a_10227_46804# a_10807_43548# 0.025916f
C14130 a_8049_45260# a_3357_43084# 0.08902f
C14131 a_11599_46634# a_11453_44696# 0.075707f
C14132 a_n2833_47464# a_n2442_46660# 0.055535f
C14133 a_n1151_42308# a_12549_44172# 0.466584f
C14134 a_6151_47436# a_n1613_43370# 0.548675f
C14135 a_18479_47436# a_19787_47423# 0.029306f
C14136 a_5932_42308# a_7174_31319# 13.0265f
C14137 a_15051_42282# a_15486_42560# 0.234322f
C14138 a_14113_42308# a_15764_42576# 0.229529f
C14139 a_2479_44172# a_2905_42968# 0.163227f
C14140 a_n97_42460# a_2982_43646# 0.180648f
C14141 a_15493_43396# a_16867_43762# 0.02646f
C14142 a_n913_45002# a_10533_42308# 0.246621f
C14143 a_n2661_45546# a_n699_43396# 0.022358f
C14144 a_n863_45724# a_n452_44636# 0.01836f
C14145 a_19479_31679# a_3357_43084# 0.058337f
C14146 a_7499_43078# a_n2661_43370# 0.027764f
C14147 a_10227_46804# a_20273_46660# 0.037464f
C14148 a_n237_47217# a_4704_46090# 0.042359f
C14149 a_2063_45854# a_167_45260# 0.359284f
C14150 a_18597_46090# a_19123_46287# 0.188676f
C14151 a_18479_47436# a_20107_46660# 0.019527f
C14152 a_13657_42558# VDD 0.195727f
C14153 a_n3565_39304# a_n4064_37440# 0.028266f
C14154 a_n4064_39072# a_n3565_37414# 0.03075f
C14155 a_n3420_39072# a_n3420_37440# 0.052876f
C14156 a_22485_38105# a_22537_39537# 0.559814f
C14157 a_20301_43646# a_20556_43646# 0.114664f
C14158 a_2437_43646# VDD 1.17411f
C14159 a_20447_31679# C5_N_btm 0.040445f
C14160 a_3422_30871# COMP_P 0.208163f
C14161 a_n2661_45010# a_n23_44458# 0.049334f
C14162 a_3232_43370# a_5518_44484# 0.01014f
C14163 C7_N_btm VDD 0.121904f
C14164 C7_P_btm VCM 1.58335f
C14165 C6_P_btm VREF_GND 0.836236f
C14166 C5_P_btm VREF 0.987144f
C14167 C9_N_btm C10_N_btm 53.3168f
C14168 C3_P_btm VIN_P 0.455045f
C14169 a_4905_42826# a_4921_42308# 0.046918f
C14170 a_14537_43396# a_15682_43940# 0.01288f
C14171 a_1307_43914# a_10807_43548# 0.016974f
C14172 a_13720_44458# a_13857_44734# 0.126609f
C14173 a_20202_43084# a_21356_42826# 0.011854f
C14174 a_9625_46129# a_8049_45260# 0.04571f
C14175 a_n1613_43370# a_5111_44636# 0.601769f
C14176 a_768_44030# a_413_45260# 0.182253f
C14177 a_12465_44636# a_14180_45002# 0.015526f
C14178 a_5342_30871# a_15051_42282# 0.029795f
C14179 a_2382_45260# a_3681_42891# 0.067836f
C14180 a_14539_43914# a_n97_42460# 0.05616f
C14181 a_2998_44172# a_3600_43914# 0.012242f
C14182 a_n913_45002# a_10835_43094# 0.053818f
C14183 a_n1059_45260# a_10796_42968# 0.01348f
C14184 a_n2661_46634# VDD 2.23057f
C14185 a_16327_47482# a_20512_43084# 0.118893f
C14186 a_n2293_46098# a_5111_44636# 0.086926f
C14187 a_4185_45028# a_n913_45002# 0.855072f
C14188 a_3316_45546# a_3175_45822# 0.05019f
C14189 a_3503_45724# a_2711_45572# 0.058013f
C14190 a_13259_45724# a_11823_42460# 0.626941f
C14191 a_4646_46812# a_6298_44484# 1.65052f
C14192 a_4915_47217# a_5129_47502# 0.070911f
C14193 a_4791_45118# a_6151_47436# 0.019937f
C14194 a_14543_43071# VDD 0.18866f
C14195 a_9313_44734# a_10341_42308# 0.019286f
C14196 a_8199_44636# VDD 1.43837f
C14197 a_10193_42453# a_19511_42282# 0.133376f
C14198 a_5937_45572# a_6109_44484# 0.163331f
C14199 a_2711_45572# a_14180_45002# 0.147337f
C14200 a_12741_44636# a_17517_44484# 0.01998f
C14201 a_8016_46348# a_5891_43370# 0.183035f
C14202 a_17715_44484# a_17767_44458# 0.07408f
C14203 a_n2661_46634# a_n2312_38680# 0.106815f
C14204 a_1666_39587# a_1169_39043# 0.036194f
C14205 a_n4209_39304# a_n4064_39072# 0.19711f
C14206 a_1606_42308# C1_P_btm 0.096405f
C14207 a_14097_32519# VIN_N 0.052362f
C14208 a_n3565_39304# a_n3420_39072# 0.241179f
C14209 COMP_P VDD 3.52636f
C14210 a_10341_43396# a_17324_43396# 0.010417f
C14211 a_5343_44458# a_7963_42308# 0.108654f
C14212 a_n356_44636# a_1184_42692# 0.03675f
C14213 a_15681_43442# a_15781_43660# 0.167615f
C14214 a_15227_44166# a_15681_43442# 0.015868f
C14215 a_22959_45572# a_22959_45036# 0.026152f
C14216 a_n863_45724# a_n809_44244# 0.016179f
C14217 a_4558_45348# a_n2661_43370# 0.018142f
C14218 a_n1151_42308# a_n2661_45546# 0.044338f
C14219 a_18597_46090# a_8049_45260# 0.047215f
C14220 a_n971_45724# a_3316_45546# 0.086835f
C14221 a_11599_46634# a_14180_46482# 0.016275f
C14222 a_n2293_46634# a_8953_45546# 0.04453f
C14223 a_18834_46812# a_15227_44166# 0.231715f
C14224 a_8128_46384# a_6945_45028# 0.010979f
C14225 a_5807_45002# a_14275_46494# 0.013842f
C14226 a_13747_46662# a_13925_46122# 0.020304f
C14227 a_n3565_37414# VDD 0.785032f
C14228 VDAC_P C2_P_btm 3.46245f
C14229 a_15279_43071# a_5342_30871# 0.214197f
C14230 a_9290_44172# a_13635_43156# 0.394766f
C14231 a_18494_42460# a_9313_44734# 0.028817f
C14232 w_1575_34786# a_n3420_39072# 0.024342f
C14233 a_10227_46804# a_15959_42545# 0.152289f
C14234 a_3537_45260# a_3905_42865# 0.258917f
C14235 a_13747_46662# a_15599_45572# 0.041358f
C14236 a_4791_45118# a_5111_44636# 1.11355f
C14237 a_n2497_47436# a_375_42282# 0.018989f
C14238 a_5257_43370# a_6194_45824# 0.029055f
C14239 a_8016_46348# a_9290_44172# 0.020766f
C14240 a_n2293_46098# a_n2956_38680# 0.022177f
C14241 a_743_42282# a_15051_42282# 0.011096f
C14242 a_n2293_43922# a_n3674_39768# 0.018871f
C14243 a_10057_43914# a_10555_44260# 0.041594f
C14244 a_4185_45028# a_1755_42282# 0.023564f
C14245 a_1823_45246# a_3823_42558# 0.137565f
C14246 a_18143_47464# VDD 0.388551f
C14247 a_10809_44734# a_7499_43078# 0.053075f
C14248 a_3090_45724# a_6171_45002# 0.030689f
C14249 a_768_44030# a_2779_44458# 0.014949f
C14250 a_21259_43561# VDD 0.192954f
C14251 a_5342_30871# a_n3420_37440# 0.030303f
C14252 a_n2104_42282# a_n1794_35082# 0.030917f
C14253 COMP_P a_n784_42308# 0.109134f
C14254 a_5534_30871# a_n4064_37440# 0.041703f
C14255 a_13678_32519# C2_N_btm 0.03058f
C14256 a_n961_42308# a_n473_42460# 0.011409f
C14257 a_20205_31679# a_13258_32519# 0.054848f
C14258 a_765_45546# VDD 2.19953f
C14259 a_1467_44172# a_1427_43646# 0.104539f
C14260 a_3090_45724# a_14673_44172# 0.018197f
C14261 a_13661_43548# a_18451_43940# 0.129334f
C14262 a_n755_45592# a_n745_45366# 0.014023f
C14263 a_584_46384# a_3626_43646# 0.195961f
C14264 a_11415_45002# a_14539_43914# 0.010769f
C14265 a_n2293_45546# a_n143_45144# 0.012062f
C14266 a_1138_42852# a_949_44458# 0.013552f
C14267 a_4185_45028# a_n2661_44458# 0.030414f
C14268 a_12549_44172# a_15493_43940# 0.932577f
C14269 a_n1151_42308# a_5385_46902# 0.0125f
C14270 a_11453_44696# a_13661_43548# 0.099457f
C14271 a_21496_47436# a_20916_46384# 0.113102f
C14272 a_n237_47217# a_7715_46873# 0.051915f
C14273 a_n971_45724# a_8145_46902# 0.051701f
C14274 a_n3674_37592# a_n4209_37414# 0.044977f
C14275 a_22400_42852# a_22589_40599# 0.135364f
C14276 a_n2956_37592# a_n4209_39590# 0.090416f
C14277 a_509_45822# VDD 0.190119f
C14278 a_16327_47482# a_18249_42858# 0.315855f
C14279 a_2382_45260# a_3232_43370# 0.239776f
C14280 a_2437_43646# a_1423_45028# 0.023818f
C14281 a_9049_44484# a_8701_44490# 0.100038f
C14282 a_7499_43078# a_5883_43914# 0.100372f
C14283 a_4574_45260# a_4558_45348# 0.19344f
C14284 a_3537_45260# a_5147_45002# 0.092965f
C14285 a_n863_45724# a_n2661_42834# 0.094705f
C14286 a_20916_46384# a_21363_46634# 0.017401f
C14287 a_n1613_43370# a_n1423_46090# 0.15966f
C14288 a_11599_46634# a_13925_46122# 0.549622f
C14289 a_10227_46804# a_10355_46116# 0.022564f
C14290 a_n971_45724# a_5066_45546# 0.045749f
C14291 a_6151_47436# a_6945_45028# 0.335681f
C14292 a_12549_44172# a_12741_44636# 0.090958f
C14293 a_n4209_39304# VDD 1.01306f
C14294 a_n3565_39590# VIN_P 0.067869f
C14295 VDAC_Ni a_5700_37509# 0.079762f
C14296 a_3754_38470# a_4338_37500# 0.473597f
C14297 a_n3565_37414# a_n2302_37690# 0.046906f
C14298 a_n3690_37440# a_n4064_37440# 0.085414f
C14299 a_n3420_37440# a_n2946_37690# 0.236674f
C14300 a_n4209_39590# VREF 0.860047f
C14301 a_n2661_42282# a_n1794_35082# 0.093522f
C14302 a_11967_42832# a_17124_42282# 0.067231f
C14303 a_16751_45260# VDD 0.121848f
C14304 a_13259_45724# a_2982_43646# 0.06616f
C14305 a_4185_45028# a_17364_32525# 0.046035f
C14306 a_8953_45546# a_743_42282# 0.032209f
C14307 a_n913_45002# a_11967_42832# 0.156551f
C14308 a_413_45260# a_17517_44484# 0.013023f
C14309 a_6755_46942# a_8049_45260# 0.035035f
C14310 a_15227_44166# a_10809_44734# 0.034868f
C14311 a_13059_46348# a_13351_46090# 0.074689f
C14312 a_11599_46634# a_15599_45572# 0.26676f
C14313 a_n2497_47436# a_2437_43646# 0.027407f
C14314 a_n2157_46122# a_n1991_46122# 0.614266f
C14315 a_19692_46634# a_21137_46414# 0.242332f
C14316 a_n2293_46634# a_1609_45822# 0.036096f
C14317 a_5807_45002# a_6194_45824# 0.02442f
C14318 a_3626_43646# a_17303_42282# 0.037411f
C14319 a_4223_44672# a_7542_44172# 0.052366f
C14320 a_16922_45042# a_20269_44172# 0.010825f
C14321 a_14815_43914# a_14673_44172# 0.173231f
C14322 a_n2312_38680# a_n4209_39304# 0.062228f
C14323 a_n2497_47436# a_4181_44734# 0.01129f
C14324 a_3877_44458# a_3065_45002# 0.287919f
C14325 a_18597_46090# a_20193_45348# 0.021804f
C14326 a_5164_46348# a_2711_45572# 0.031464f
C14327 a_6452_43396# VDD 0.083252f
C14328 a_4190_30871# a_n4064_37440# 0.032722f
C14329 a_14635_42282# a_14853_42852# 0.01129f
C14330 a_5534_30871# a_n3420_39072# 0.339008f
C14331 a_10193_42453# a_13291_42460# 0.050019f
C14332 a_10623_46897# VDD 0.189083f
C14333 a_5891_43370# a_8791_43396# 0.194389f
C14334 a_n755_45592# a_2123_42473# 0.022891f
C14335 a_18579_44172# a_19319_43548# 0.031277f
C14336 a_8162_45546# a_7499_43078# 0.021916f
C14337 a_768_44030# a_644_44056# 0.177755f
C14338 a_8199_44636# a_1423_45028# 0.088277f
C14339 a_11415_45002# a_14309_45028# 0.040538f
C14340 a_8049_45260# a_19479_31679# 0.022565f
C14341 a_10227_46804# a_20894_47436# 0.010908f
C14342 a_18780_47178# a_18597_46090# 0.175179f
C14343 a_18479_47436# a_19386_47436# 0.219411f
C14344 a_16327_47482# a_4883_46098# 0.096832f
C14345 a_n2497_47436# a_n2661_46634# 0.079801f
C14346 a_2905_45572# a_768_44030# 0.02789f
C14347 a_n1151_42308# a_12891_46348# 0.038292f
C14348 a_5815_47464# a_n1613_43370# 0.360237f
C14349 a_11551_42558# a_11897_42308# 0.013377f
C14350 a_14113_42308# a_15486_42560# 0.039784f
C14351 a_n4318_37592# a_n4064_39072# 0.019896f
C14352 a_1568_43370# a_1756_43548# 0.094732f
C14353 a_n97_42460# a_2896_43646# 0.027089f
C14354 a_2479_44172# a_2075_43172# 0.034186f
C14355 a_15493_43396# a_16664_43396# 0.016417f
C14356 a_375_42282# a_196_42282# 0.165785f
C14357 a_n2293_46098# a_3905_42865# 0.237656f
C14358 a_13661_43548# a_9145_43396# 0.135139f
C14359 a_n2661_45546# a_4223_44672# 0.041115f
C14360 a_8696_44636# a_8953_45002# 0.018854f
C14361 a_22223_45572# a_3357_43084# 0.07533f
C14362 a_2711_45572# a_18494_42460# 0.1183f
C14363 a_8746_45002# a_8560_45348# 0.044092f
C14364 a_12549_44172# a_13607_46688# 0.013421f
C14365 a_10227_46804# a_20411_46873# 0.013631f
C14366 a_2107_46812# a_5257_43370# 0.039927f
C14367 a_n237_47217# a_4419_46090# 0.049065f
C14368 a_584_46384# a_167_45260# 0.0321f
C14369 a_18597_46090# a_18285_46348# 0.012666f
C14370 a_2063_45854# a_2202_46116# 0.026352f
C14371 a_n2946_37984# a_n2860_37984# 0.011479f
C14372 a_22485_38105# a_22889_38993# 0.089418f
C14373 a_20301_43646# a_743_42282# 0.09203f
C14374 a_21513_45002# VDD 0.416919f
C14375 a_4190_30871# a_20556_43646# 0.021112f
C14376 a_21259_43561# a_21487_43396# 0.08444f
C14377 a_17339_46660# a_19095_43396# 0.049229f
C14378 a_5205_44484# a_4223_44672# 0.235572f
C14379 a_n2661_45010# a_n356_44636# 0.091266f
C14380 a_3232_43370# a_5343_44458# 0.654021f
C14381 SMPL_ON_P a_n4318_38216# 0.037528f
C14382 a_n1925_46634# a_8034_45724# 0.206805f
C14383 a_6151_47436# a_6812_45938# 0.018338f
C14384 C6_N_btm VDD 0.210613f
C14385 C7_P_btm VREF_GND 1.61142f
C14386 C8_P_btm VCM 2.61094f
C14387 C6_P_btm VREF 1.41944f
C14388 C8_N_btm C10_N_btm 2.07867f
C14389 C4_P_btm VIN_P 0.50261f
C14390 a_n2810_45572# a_n4318_38680# 0.023234f
C14391 a_22223_45036# a_22315_44484# 0.011923f
C14392 a_14537_43396# a_14955_43940# 0.104291f
C14393 a_1307_43914# a_10949_43914# 0.062121f
C14394 a_n2312_39304# a_n4209_39590# 0.065703f
C14395 a_n2293_42834# a_7542_44172# 0.010138f
C14396 a_22612_30879# a_20447_31679# 0.107874f
C14397 a_10809_44734# a_22959_46124# 0.172346f
C14398 a_2324_44458# a_n1925_42282# 0.018757f
C14399 a_8953_45546# a_8049_45260# 0.156816f
C14400 a_5342_30871# a_14113_42308# 0.203397f
C14401 a_4190_30871# a_n3420_39072# 0.10848f
C14402 a_n1549_44318# a_n1453_44318# 0.013793f
C14403 a_11967_42832# a_18451_43940# 0.01235f
C14404 a_n699_43396# a_n1557_42282# 0.02911f
C14405 a_n913_45002# a_10518_42984# 0.058603f
C14406 a_5807_45002# CLK 0.033646f
C14407 a_n2956_39768# VDD 0.697168f
C14408 a_5257_43370# a_n2661_44458# 0.027109f
C14409 a_10586_45546# a_10907_45822# 0.05477f
C14410 a_n2293_46098# a_5147_45002# 0.211057f
C14411 a_5937_45572# a_3357_43084# 0.257963f
C14412 a_4185_45028# a_n1059_45260# 0.027781f
C14413 a_4791_45118# a_3905_42865# 0.208831f
C14414 a_3316_45546# a_2711_45572# 0.065336f
C14415 a_3218_45724# a_3175_45822# 0.132424f
C14416 a_n443_46116# a_5129_47502# 0.10632f
C14417 a_2063_45854# a_9313_45822# 0.042979f
C14418 a_5342_30871# C8_N_btm 0.093874f
C14419 a_6171_42473# a_5932_42308# 0.224949f
C14420 a_13460_43230# VDD 0.276534f
C14421 a_8349_46414# VDD 0.209819f
C14422 a_n2810_45572# a_n4209_38216# 0.195791f
C14423 a_7499_43078# a_3537_45260# 0.586701f
C14424 a_13259_45724# a_14309_45028# 0.063402f
C14425 a_1823_45246# a_n2661_43922# 0.441151f
C14426 a_5807_45002# a_2107_46812# 1.5594f
C14427 a_n2956_39768# a_n2312_38680# 0.076511f
C14428 a_n2472_46634# a_n2293_46634# 0.163804f
C14429 a_n2661_46634# a_n2104_46634# 0.030211f
C14430 a_n3565_39590# a_n3565_38502# 0.031189f
C14431 a_1169_39587# a_1169_39043# 0.054961f
C14432 a_n4209_39304# a_n2946_39072# 0.022779f
C14433 a_n4209_39590# a_n3420_38528# 0.032196f
C14434 a_1606_42308# C2_P_btm 0.021793f
C14435 a_n3420_39616# a_n4209_38502# 0.028008f
C14436 a_n3565_39304# a_n3690_39392# 0.247167f
C14437 a_n4318_37592# VDD 0.919667f
C14438 a_n97_42460# a_7227_42852# 0.117893f
C14439 a_10341_43396# a_17499_43370# 0.022768f
C14440 a_20202_43084# a_2982_43646# 0.034798f
C14441 a_1138_42852# a_n97_42460# 0.015603f
C14442 a_7499_43078# a_11541_44484# 0.048175f
C14443 a_n1925_46634# a_8016_46348# 0.014574f
C14444 a_12251_46660# a_12347_46660# 0.013793f
C14445 a_n237_47217# a_1848_45724# 0.232571f
C14446 a_584_46384# a_n863_45724# 0.051089f
C14447 a_17609_46634# a_15227_44166# 0.04317f
C14448 a_n2661_46098# a_1138_42852# 0.020229f
C14449 a_13747_46662# a_13759_46122# 0.02887f
C14450 a_n4334_37440# VDD 0.385859f
C14451 VDAC_P C3_P_btm 6.90991f
C14452 a_5534_30871# a_5342_30871# 11.128201f
C14453 a_22959_45036# VDD 0.30999f
C14454 a_3537_45260# a_3600_43914# 0.157156f
C14455 a_18184_42460# a_9313_44734# 0.069472f
C14456 a_10227_46804# a_15803_42450# 0.296174f
C14457 a_10903_43370# a_12379_42858# 0.02509f
C14458 a_n2312_38680# a_n4318_37592# 0.02327f
C14459 a_13661_43548# a_15599_45572# 0.01321f
C14460 a_4791_45118# a_5147_45002# 0.10845f
C14461 a_5257_43370# a_5907_45546# 0.064039f
C14462 a_n2472_46090# a_n2956_38680# 0.157373f
C14463 a_18479_47436# a_3357_43084# 0.292061f
C14464 a_743_42282# a_14113_42308# 0.015227f
C14465 a_n2661_43922# a_n3674_39768# 0.152656f
C14466 a_18989_43940# a_18451_43940# 0.114286f
C14467 a_20835_44721# a_21145_44484# 0.013793f
C14468 a_1823_45246# a_3318_42354# 0.055532f
C14469 a_10227_46804# VDD 2.77567f
C14470 a_5066_45546# a_2711_45572# 0.090644f
C14471 a_3090_45724# a_3232_43370# 0.024183f
C14472 a_11189_46129# a_10907_45822# 0.021145f
C14473 a_5937_45572# a_9159_45572# 0.048183f
C14474 w_1575_34786# w_10694_33990# 0.119791f
C14475 a_n3674_38216# a_n3674_37592# 0.048035f
C14476 a_n4318_38216# a_n1794_35082# 0.031712f
C14477 a_4190_30871# C10_N_btm 0.446355f
C14478 a_n913_45002# a_n2293_42282# 0.028018f
C14479 a_17339_46660# VDD 0.555596f
C14480 a_n356_44636# a_5649_42852# 0.023625f
C14481 a_12741_44636# a_13076_44458# 0.010522f
C14482 a_13661_43548# a_18326_43940# 0.024789f
C14483 a_n2661_45546# a_413_45260# 0.022797f
C14484 a_n755_45592# a_n913_45002# 0.347782f
C14485 a_526_44458# a_2809_45028# 0.033247f
C14486 a_n443_46116# a_1756_43548# 0.046156f
C14487 a_10809_44734# a_n2661_43370# 0.077978f
C14488 a_10907_45822# a_11136_45572# 0.080042f
C14489 a_n2293_45546# a_n467_45028# 0.067105f
C14490 a_1138_42852# a_742_44458# 0.040731f
C14491 a_584_46384# a_3540_43646# 0.045907f
C14492 a_n1151_42308# a_n1557_42282# 0.214486f
C14493 a_n443_42852# a_3357_43084# 0.042246f
C14494 a_n1151_42308# a_4817_46660# 0.029921f
C14495 a_n237_47217# a_7411_46660# 0.033907f
C14496 a_11453_44696# a_5807_45002# 0.050036f
C14497 a_13507_46334# a_20916_46384# 0.123008f
C14498 a_n971_45724# a_7577_46660# 0.523694f
C14499 a_13258_32519# a_21335_42336# 0.022004f
C14500 a_20107_42308# a_7174_31319# 0.175129f
C14501 a_n2810_45028# a_n4209_39590# 0.021994f
C14502 a_7499_43078# a_8701_44490# 0.011795f
C14503 a_22612_30879# a_13467_32519# 0.061222f
C14504 a_8953_45546# a_9028_43914# 0.01093f
C14505 a_3537_45260# a_4558_45348# 0.236111f
C14506 a_4883_46098# a_5204_45822# 0.041898f
C14507 a_11599_46634# a_13759_46122# 0.262969f
C14508 a_n881_46662# a_n1853_46287# 0.229188f
C14509 a_n1613_43370# a_n1991_46122# 0.031697f
C14510 a_4915_47217# a_10809_44734# 0.037616f
C14511 a_12891_46348# a_12741_44636# 0.038901f
C14512 a_10249_46116# a_6755_46942# 0.068878f
C14513 a_n3565_38502# C4_P_btm 0.042623f
C14514 a_1273_38525# VDD 3.23397f
C14515 VDAC_Ni a_5088_37509# 1.70462f
C14516 a_3754_38470# a_3726_37500# 0.554457f
C14517 a_n3565_37414# a_n4064_37440# 0.230258f
C14518 a_743_42282# a_5534_30871# 0.030281f
C14519 a_4190_30871# a_5342_30871# 0.0276f
C14520 a_1307_43914# VDD 3.92807f
C14521 a_4185_45028# a_22959_43396# 0.01521f
C14522 a_n1059_45260# a_11967_42832# 0.627158f
C14523 a_13059_46348# a_12594_46348# 0.03479f
C14524 a_n1613_43370# a_7499_43078# 0.324998f
C14525 a_n2157_46122# a_n1853_46287# 0.617317f
C14526 a_n2293_46098# a_n1991_46122# 0.01544f
C14527 a_19692_46634# a_20708_46348# 0.318388f
C14528 a_5807_45002# a_5907_45546# 0.013402f
C14529 a_n2293_46634# a_n443_42852# 2.09483f
C14530 a_3626_43646# a_4958_30871# 0.087921f
C14531 a_18579_44172# VDD 0.38178f
C14532 a_4223_44672# a_7281_43914# 0.01814f
C14533 a_16922_45042# a_19862_44208# 0.038132f
C14534 a_11453_44696# a_18315_45260# 0.010513f
C14535 a_13059_46348# a_15037_45618# 0.064109f
C14536 a_3090_45724# a_18341_45572# 0.016963f
C14537 a_n881_46662# a_n2661_43370# 0.020731f
C14538 a_9396_43370# VDD 0.288403f
C14539 a_n2293_42282# a_1755_42282# 0.875855f
C14540 a_n2293_42834# a_4520_42826# 0.01065f
C14541 a_18184_42460# a_13887_32519# 0.03303f
C14542 a_5891_43370# a_8147_43396# 0.029069f
C14543 a_10467_46802# VDD 0.401016f
C14544 a_n755_45592# a_1755_42282# 1.52791f
C14545 a_n863_45724# a_2713_42308# 0.044499f
C14546 a_8162_45546# a_8568_45546# 0.078784f
C14547 a_8049_45260# a_22223_45572# 0.013885f
C14548 a_12861_44030# a_15493_43396# 0.254093f
C14549 a_10227_46804# a_19787_47423# 0.03269f
C14550 a_18479_47436# a_18597_46090# 0.473843f
C14551 a_n2833_47464# a_n2661_46634# 0.011033f
C14552 a_n1151_42308# a_11309_47204# 0.546434f
C14553 a_4915_47217# a_n881_46662# 1.23372f
C14554 a_14113_42308# a_15051_42282# 0.077852f
C14555 a_n2661_42282# a_4361_42308# 0.034761f
C14556 a_2479_44172# a_1847_42826# 0.141223f
C14557 a_8034_45724# VDD 0.812726f
C14558 a_19862_44208# a_15743_43084# 0.022478f
C14559 a_4185_45028# a_22959_44484# 0.011365f
C14560 a_n755_45592# a_n2661_44458# 0.023853f
C14561 a_2437_43646# a_3357_43084# 0.424652f
C14562 a_22223_45572# a_19479_31679# 0.155323f
C14563 a_2711_45572# a_18184_42460# 0.367034f
C14564 a_18597_46090# a_4190_30871# 0.022042f
C14565 a_10227_46804# a_20107_46660# 0.312495f
C14566 a_n237_47217# a_4185_45028# 0.074951f
C14567 a_n443_46116# a_n1853_46287# 0.013261f
C14568 a_12465_44636# a_13059_46348# 0.163448f
C14569 a_2063_45854# a_1823_45246# 0.038948f
C14570 a_n4209_39304# a_n4064_37440# 0.029715f
C14571 a_2684_37794# VDAC_Pi 0.133177f
C14572 a_n3565_39304# a_n3420_37440# 0.032339f
C14573 a_n4064_39072# a_n4209_37414# 0.030589f
C14574 a_n3420_39072# a_n3565_37414# 0.031846f
C14575 a_22485_38105# a_22613_38993# 0.253409f
C14576 a_4958_30871# C9_P_btm 0.209166f
C14577 a_4190_30871# a_743_42282# 0.18536f
C14578 a_n2017_45002# a_n2012_44484# 0.013231f
C14579 a_4791_45118# a_7499_43078# 0.024468f
C14580 C5_N_btm VDD 0.267489f
C14581 C8_P_btm VREF_GND 2.58605f
C14582 C9_P_btm VCM 6.06251f
C14583 C7_P_btm VREF 1.818f
C14584 C7_N_btm C10_N_btm 1.39624f
C14585 C8_N_btm C9_N_btm 39.4538f
C14586 C5_P_btm VIN_P 0.502041f
C14587 a_n2810_45572# a_n3674_39304# 0.023379f
C14588 a_11827_44484# a_22315_44484# 0.013f
C14589 a_22223_45036# a_3422_30871# 0.011196f
C14590 a_1307_43914# a_10729_43914# 0.051086f
C14591 a_13076_44458# a_13468_44734# 0.016359f
C14592 a_18494_42460# a_20512_43084# 0.115057f
C14593 a_20202_43084# a_19987_42826# 0.177726f
C14594 a_n443_42852# a_743_42282# 0.03363f
C14595 a_3090_45724# a_10193_42453# 0.027088f
C14596 a_21588_30879# a_20447_31679# 0.055937f
C14597 a_n2661_46634# a_3357_43084# 0.032385f
C14598 a_12465_44636# a_13556_45296# 0.248126f
C14599 a_2324_44458# a_526_44458# 0.279023f
C14600 a_5937_45572# a_8049_45260# 0.103218f
C14601 a_13059_46348# a_2711_45572# 0.075233f
C14602 a_n2293_46634# a_2437_43646# 0.030387f
C14603 a_n443_46116# a_n2661_43370# 0.030763f
C14604 a_11967_42832# a_18326_43940# 0.058879f
C14605 a_2889_44172# a_2998_44172# 0.179664f
C14606 a_n1549_44318# a_n1644_44306# 0.049827f
C14607 a_n913_45002# a_10083_42826# 0.052028f
C14608 a_22612_30879# RST_Z 0.058603f
C14609 a_20916_46384# SINGLE_ENDED 0.020511f
C14610 a_n2840_46634# VDD 0.306342f
C14611 a_13259_45724# a_11962_45724# 0.026896f
C14612 a_4646_46812# a_5343_44458# 0.24395f
C14613 a_6755_46942# a_11691_44458# 0.192426f
C14614 a_768_44030# a_n2293_43922# 0.027199f
C14615 a_10586_45546# a_10210_45822# 0.042978f
C14616 a_n2293_46098# a_4558_45348# 0.030863f
C14617 a_3218_45724# a_2711_45572# 0.1731f
C14618 a_2957_45546# a_3175_45822# 0.08213f
C14619 a_4185_45028# a_n2017_45002# 0.029634f
C14620 a_n443_46116# a_4915_47217# 0.395101f
C14621 a_4791_45118# a_5129_47502# 0.240381f
C14622 a_5755_42308# a_5932_42308# 0.196877f
C14623 a_3823_42558# a_4169_42308# 0.013377f
C14624 a_13635_43156# VDD 0.463701f
C14625 a_3483_46348# CLK 0.408122f
C14626 a_8016_46348# VDD 1.42798f
C14627 a_1138_42852# a_n2661_43922# 0.027736f
C14628 a_768_44030# a_n97_42460# 0.034422f
C14629 a_1823_45246# a_n2661_42834# 0.174801f
C14630 w_10694_33990# a_4190_30871# 0.036996f
C14631 a_n443_42852# a_626_44172# 0.028669f
C14632 a_n2840_46634# a_n2312_38680# 0.040373f
C14633 a_n2661_46634# a_n2293_46634# 0.060962f
C14634 a_n2472_46634# a_n2442_46660# 0.155358f
C14635 a_n1736_42282# VDD 0.227152f
C14636 a_n4209_39304# a_n3420_39072# 0.071714f
C14637 a_n97_42460# a_5755_42852# 0.149651f
C14638 a_10341_43396# a_16759_43396# 0.010617f
C14639 a_11682_45822# VDD 0.316586f
C14640 a_n356_44636# a_1067_42314# 0.019369f
C14641 a_3537_45260# a_n2661_43370# 0.087747f
C14642 a_1307_43914# a_1423_45028# 0.054616f
C14643 a_375_42282# a_626_44172# 0.017957f
C14644 a_18479_47436# a_8049_45260# 0.047429f
C14645 a_2107_46812# a_3483_46348# 0.100707f
C14646 a_n2293_46634# a_8199_44636# 0.029753f
C14647 a_n881_46662# a_10809_44734# 0.026121f
C14648 a_n2661_46098# a_1176_45822# 0.144277f
C14649 a_5807_45002# a_13925_46122# 0.027158f
C14650 a_n4209_37414# VDD 0.819451f
C14651 VDAC_P C4_P_btm 13.8049f
C14652 a_8530_39574# RST_Z 0.431385f
C14653 a_22223_45036# VDD 0.300162f
C14654 a_3537_45260# a_2998_44172# 0.059736f
C14655 a_3065_45002# a_3905_42865# 0.034773f
C14656 a_n443_42852# a_2813_43396# 0.017355f
C14657 a_3232_43370# a_1414_42308# 0.248035f
C14658 a_13259_45724# a_17499_43370# 0.018042f
C14659 a_10227_46804# a_15764_42576# 0.024352f
C14660 a_n2497_47436# a_1307_43914# 0.069365f
C14661 a_8199_44636# a_9625_46129# 0.011574f
C14662 a_5937_45572# a_8953_45546# 0.3871f
C14663 a_4791_45118# a_4558_45348# 0.077256f
C14664 a_5257_43370# a_5263_45724# 0.088982f
C14665 a_n2840_46090# a_n2956_38680# 0.050916f
C14666 a_8016_46348# a_9823_46155# 0.048283f
C14667 a_n1151_42308# a_6171_45002# 0.02292f
C14668 a_5342_30871# COMP_P 0.027184f
C14669 a_n2293_42834# a_n1557_42282# 0.034384f
C14670 a_n2661_43922# a_n4318_39768# 0.010131f
C14671 a_5891_43370# a_n2661_42282# 0.032052f
C14672 a_n2661_42834# a_n3674_39768# 0.150968f
C14673 a_17591_47464# VDD 0.421992f
C14674 a_768_44030# a_742_44458# 0.216263f
C14675 a_9290_44172# a_10907_45822# 0.262972f
C14676 a_765_45546# a_3357_43084# 0.035297f
C14677 a_8199_44636# a_9159_45572# 0.049711f
C14678 a_5534_30871# a_n3420_37440# 0.04166f
C14679 a_n2472_42282# a_n1794_35082# 0.040716f
C14680 a_n357_42282# a_17124_42282# 0.011823f
C14681 a_n1059_45260# a_n2293_42282# 0.033257f
C14682 a_12741_44636# a_12883_44458# 0.073263f
C14683 a_13661_43548# a_18079_43940# 0.028277f
C14684 a_n755_45592# a_n1059_45260# 0.53237f
C14685 a_n357_42282# a_n913_45002# 0.309845f
C14686 a_n443_46116# a_1568_43370# 0.584982f
C14687 a_584_46384# a_2982_43646# 0.057754f
C14688 a_11823_42460# a_8696_44636# 0.026654f
C14689 a_12549_44172# a_11341_43940# 0.406618f
C14690 a_3483_46348# a_n2661_44458# 1.44355f
C14691 VCM VSS 30.7117f
C14692 VREF_GND VSS 17.6497f
C14693 VREF VSS 8.8492f
C14694 VIN_N VSS 13.0509f
C14695 VIN_P VSS 13.027599f
C14696 CLK VSS 1.55797f
C14697 EN_OFFSET_CAL VSS 0.505642f
C14698 DATA[5] VSS 0.561058f
C14699 DATA[4] VSS 0.755679f
C14700 DATA[3] VSS 1.01838f
C14701 DATA[2] VSS 0.536983f
C14702 DATA[1] VSS 0.550109f
C14703 DATA[0] VSS 0.616231f
C14704 CLK_DATA VSS 0.488979f
C14705 SINGLE_ENDED VSS 0.60168f
C14706 START VSS 0.991673f
C14707 RST_Z VSS 11.3723f
C14708 VDD VSS 0.589065p
C14709 C10_N_btm VSS 0.210692p
C14710 C9_N_btm VSS 79.926506f
C14711 C8_N_btm VSS 45.547f
C14712 C7_N_btm VSS 25.886099f
C14713 C6_N_btm VSS 15.5273f
C14714 C5_N_btm VSS 9.624539f
C14715 C4_N_btm VSS 8.794849f
C14716 C3_N_btm VSS 6.38289f
C14717 C2_N_btm VSS 5.46028f
C14718 C1_N_btm VSS 5.26099f
C14719 C0_N_btm VSS 7.20283f
C14720 C0_dummy_N_btm VSS 5.0303f
C14721 C0_dummy_P_btm VSS 5.01806f
C14722 C0_P_btm VSS 7.1984f
C14723 C1_P_btm VSS 5.27428f
C14724 C2_P_btm VSS 5.46972f
C14725 C3_P_btm VSS 6.37616f
C14726 C4_P_btm VSS 8.785789f
C14727 C5_P_btm VSS 9.614769f
C14728 C6_P_btm VSS 15.5172f
C14729 C7_P_btm VSS 25.876501f
C14730 C8_P_btm VSS 45.531998f
C14731 C9_P_btm VSS 79.8995f
C14732 C10_P_btm VSS 0.210676p
C14733 a_21753_35474# VSS 0.730911f
C14734 a_19998_34978# VSS 1.75018f
C14735 a_19250_34978# VSS 1.69804f
C14736 a_18194_34908# VSS 2.11991f
C14737 EN_VIN_BSTR_N VSS 9.06279f
C14738 a_10890_34112# VSS 15.1553f
C14739 a_n217_35014# VSS 1.73445f
C14740 EN_VIN_BSTR_P VSS 9.29511f
C14741 a_n1057_35014# VSS 15.221701f
C14742 a_n1696_34930# VSS 2.16211f
C14743 a_n1550_35448# VSS 1.7497f
C14744 a_n2002_35448# VSS 0.735333f
C14745 a_22737_36887# VSS 0.092029f
C14746 a_22737_37285# VSS 0.095943f
C14747 a_22629_37990# VSS 0.468764f
C14748 a_22725_38406# VSS 0.010928f
C14749 a_22629_38406# VSS 0.583873f
C14750 CAL_P VSS 11.403299f
C14751 a_22537_39537# VSS 2.61801f
C14752 a_22889_38993# VSS 0.497542f
C14753 a_22613_38993# VSS 0.357645f
C14754 a_22581_37893# VSS 1.83807f
C14755 a_22527_39145# VSS 2.28699f
C14756 a_22589_40055# VSS 1.23689f
C14757 a_22537_40625# VSS 1.58437f
C14758 a_22589_40599# VSS 1.83268f
C14759 CAL_N VSS 8.7111f
C14760 a_11206_38545# VSS 0.713084f
C14761 VDAC_P VSS 0.107494p
C14762 a_8912_37509# VSS 3.72815f
C14763 VDAC_N VSS 0.108083p
C14764 a_6886_37412# VSS 3.84933f
C14765 a_5700_37509# VSS 2.08109f
C14766 a_5088_37509# VSS 2.72043f
C14767 a_4338_37500# VSS 2.61032f
C14768 a_3726_37500# VSS 4.51772f
C14769 a_n2302_37690# VSS 0.514517f
C14770 a_n4064_37440# VSS 1.72323f
C14771 a_n2946_37690# VSS 0.517242f
C14772 a_n3420_37440# VSS 5.26673f
C14773 a_n3690_37440# VSS 0.548488f
C14774 a_n3565_37414# VSS 3.17522f
C14775 a_n4334_37440# VSS 0.561497f
C14776 a_n4209_37414# VSS 3.16447f
C14777 a_8530_39574# VSS 2.76298f
C14778 a_7754_38470# VSS 3.2456f
C14779 a_3754_38470# VSS 4.77711f
C14780 VDAC_Ni VSS 2.86578f
C14781 a_7754_38636# VSS 0.353706f
C14782 a_3754_38802# VSS 0.390074f
C14783 a_7754_38968# VSS 0.330037f
C14784 a_3754_39134# VSS 0.401983f
C14785 a_7754_39300# VSS 0.330682f
C14786 a_3754_39466# VSS 0.401172f
C14787 a_7754_39632# VSS 0.340942f
C14788 VDAC_Pi VSS 3.50497f
C14789 a_7754_39964# VSS 2.62481f
C14790 a_7754_40130# VSS 2.84033f
C14791 a_3754_39964# VSS 0.671366f
C14792 a_2113_38308# VSS 2.6473f
C14793 a_n2302_37984# VSS 0.483504f
C14794 a_n4064_37984# VSS 1.65064f
C14795 a_n2946_37984# VSS 0.485942f
C14796 a_n3420_37984# VSS 1.75909f
C14797 a_n3690_38304# VSS 0.517812f
C14798 a_n3565_38216# VSS 1.49099f
C14799 a_n4334_38304# VSS 0.529531f
C14800 a_n4209_38216# VSS 3.0374f
C14801 a_2684_37794# VSS 0.414596f
C14802 a_1107_38525# VSS 0.6415f
C14803 a_n2302_38778# VSS 0.483515f
C14804 a_n4064_38528# VSS 1.69611f
C14805 a_n2946_38778# VSS 0.485895f
C14806 a_n3420_38528# VSS 2.03231f
C14807 a_n3690_38528# VSS 0.516979f
C14808 a_n3565_38502# VSS 1.56051f
C14809 a_n4334_38528# VSS 0.529888f
C14810 a_n4209_38502# VSS 3.02312f
C14811 a_2112_39137# VSS 0.414404f
C14812 comp_n VSS 0.572075f
C14813 a_1666_39043# VSS 0.909399f
C14814 a_1169_39043# VSS 0.615041f
C14815 a_n2302_39072# VSS 0.483504f
C14816 a_n4064_39072# VSS 1.71421f
C14817 a_n2946_39072# VSS 0.486447f
C14818 a_n3420_39072# VSS 2.21234f
C14819 a_n3690_39392# VSS 0.517965f
C14820 a_n3565_39304# VSS 1.4655f
C14821 a_n4334_39392# VSS 0.529516f
C14822 a_n4209_39304# VSS 3.27541f
C14823 a_1273_38525# VSS 3.59416f
C14824 a_1666_39587# VSS 1.1306f
C14825 a_1169_39587# VSS 0.633906f
C14826 a_n2302_39866# VSS 0.483537f
C14827 a_n4064_39616# VSS 2.17427f
C14828 a_n2946_39866# VSS 0.527929f
C14829 a_n3420_39616# VSS 2.10837f
C14830 a_n3690_39616# VSS 0.574329f
C14831 a_n3565_39590# VSS 2.24448f
C14832 a_n4334_39616# VSS 0.529903f
C14833 a_n4209_39590# VSS 4.03213f
C14834 a_n2302_40160# VSS 0.522244f
C14835 a_n4064_40160# VSS 3.30448f
C14836 a_n4334_40480# VSS 0.578721f
C14837 a_n4315_30879# VSS 5.0762f
C14838 a_22485_38105# VSS 1.90993f
C14839 a_22775_42308# VSS 0.602116f
C14840 a_21613_42308# VSS 0.725532f
C14841 a_21887_42336# VSS 0.234022f
C14842 a_21335_42336# VSS 0.259392f
C14843 a_7174_31319# VSS 5.50981f
C14844 a_20712_42282# VSS 0.349662f
C14845 a_20107_42308# VSS 0.344464f
C14846 a_13258_32519# VSS 6.35827f
C14847 a_19647_42308# VSS 0.313304f
C14848 a_19511_42282# VSS 0.751141f
C14849 a_19332_42282# VSS 0.31505f
C14850 a_18907_42674# VSS 0.209311f
C14851 a_18727_42674# VSS 0.233526f
C14852 a_18057_42282# VSS 0.370712f
C14853 a_17531_42308# VSS 0.253358f
C14854 a_17303_42282# VSS 1.19776f
C14855 a_4958_30871# VSS 5.01399f
C14856 a_17124_42282# VSS 0.332693f
C14857 a_16522_42674# VSS 0.073862f
C14858 a_15890_42674# VSS 0.180637f
C14859 a_15959_42545# VSS 0.263128f
C14860 a_15803_42450# VSS 0.566963f
C14861 a_15764_42576# VSS 0.298494f
C14862 a_15486_42560# VSS 0.263746f
C14863 a_15051_42282# VSS 0.790649f
C14864 a_14113_42308# VSS 1.42448f
C14865 a_14456_42282# VSS 0.33927f
C14866 a_13575_42558# VSS 0.370369f
C14867 a_13070_42354# VSS 0.222095f
C14868 a_12563_42308# VSS 0.330976f
C14869 a_11551_42558# VSS 0.372919f
C14870 a_5742_30871# VSS 7.96802f
C14871 a_11323_42473# VSS 0.253445f
C14872 a_10723_42308# VSS 0.342975f
C14873 a_10533_42308# VSS 0.310658f
C14874 a_9803_42558# VSS 0.370474f
C14875 a_9223_42460# VSS 0.236204f
C14876 a_8791_42308# VSS 0.301f
C14877 a_8685_42308# VSS 0.163732f
C14878 a_8325_42308# VSS 0.316205f
C14879 a_8515_42308# VSS 0.250762f
C14880 a_5934_30871# VSS 5.16625f
C14881 a_7963_42308# VSS 0.256292f
C14882 a_6123_31319# VSS 5.02095f
C14883 a_7227_42308# VSS 0.359705f
C14884 a_6761_42308# VSS 0.447596f
C14885 a_5932_42308# VSS 5.1182f
C14886 a_6171_42473# VSS 0.257988f
C14887 a_5755_42308# VSS 0.314735f
C14888 a_4921_42308# VSS 0.511258f
C14889 a_5379_42460# VSS 0.564806f
C14890 a_5267_42460# VSS 0.204309f
C14891 a_3823_42558# VSS 0.381485f
C14892 a_3318_42354# VSS 0.238394f
C14893 a_2903_42308# VSS 0.340659f
C14894 a_2713_42308# VSS 0.31991f
C14895 a_2351_42308# VSS 0.210162f
C14896 a_2123_42473# VSS 0.21778f
C14897 a_1755_42282# VSS 3.17706f
C14898 a_1606_42308# VSS 5.25644f
C14899 a_961_42354# VSS 0.215753f
C14900 a_1184_42692# VSS 0.222827f
C14901 a_1576_42282# VSS 0.327109f
C14902 a_1067_42314# VSS 0.32917f
C14903 a_n1794_35082# VSS 9.32119f
C14904 a_564_42282# VSS 0.36802f
C14905 a_n3674_37592# VSS 3.04613f
C14906 a_n784_42308# VSS 6.50125f
C14907 a_196_42282# VSS 0.343186f
C14908 a_n473_42460# VSS 0.366068f
C14909 a_n961_42308# VSS 0.328065f
C14910 a_n1329_42308# VSS 0.30898f
C14911 COMP_P VSS 10.955f
C14912 a_n4318_37592# VSS 1.00428f
C14913 a_n1736_42282# VSS 0.320711f
C14914 a_n3674_38216# VSS 1.68571f
C14915 a_n2104_42282# VSS 0.346472f
C14916 a_n4318_38216# VSS 0.964502f
C14917 a_n2472_42282# VSS 0.335792f
C14918 a_n3674_38680# VSS 0.881032f
C14919 a_n2840_42282# VSS 0.343361f
C14920 a_14097_32519# VSS 1.90776f
C14921 a_22400_42852# VSS 1.97851f
C14922 a_20256_43172# VSS 0.192089f
C14923 a_18504_43218# VSS 0.078212f
C14924 a_14635_42282# VSS 0.336817f
C14925 a_13291_42460# VSS 0.197331f
C14926 a_12800_43218# VSS 0.073862f
C14927 a_11554_42852# VSS 0.073028f
C14928 a_8292_43218# VSS 0.073862f
C14929 a_n2293_42282# VSS 2.62914f
C14930 a_22959_42860# VSS 0.34332f
C14931 a_22223_42860# VSS 0.328988f
C14932 a_22165_42308# VSS 0.354098f
C14933 a_21671_42860# VSS 0.316857f
C14934 a_21195_42852# VSS 0.277519f
C14935 a_21356_42826# VSS 0.304166f
C14936 a_20922_43172# VSS 0.266814f
C14937 a_19987_42826# VSS 0.378798f
C14938 a_19164_43230# VSS 0.264863f
C14939 a_19339_43156# VSS 0.471496f
C14940 a_18599_43230# VSS 0.266382f
C14941 a_18817_42826# VSS 0.182139f
C14942 a_18249_42858# VSS 0.302863f
C14943 a_17333_42852# VSS 0.29982f
C14944 a_18083_42858# VSS 0.578693f
C14945 a_17701_42308# VSS 0.179963f
C14946 a_17595_43084# VSS 0.205109f
C14947 a_16795_42852# VSS 0.362281f
C14948 a_16414_43172# VSS 0.270304f
C14949 a_15567_42826# VSS 0.316627f
C14950 a_5342_30871# VSS 4.18107f
C14951 a_15279_43071# VSS 0.248252f
C14952 a_5534_30871# VSS 4.58429f
C14953 a_14543_43071# VSS 0.246071f
C14954 a_13460_43230# VSS 0.259861f
C14955 a_13635_43156# VSS 0.7696f
C14956 a_12895_43230# VSS 0.250159f
C14957 a_13113_42826# VSS 0.174096f
C14958 a_12545_42858# VSS 0.287468f
C14959 a_12089_42308# VSS 0.283874f
C14960 a_12379_42858# VSS 0.549229f
C14961 a_10341_42308# VSS 0.317389f
C14962 a_10922_42852# VSS 0.176112f
C14963 a_10991_42826# VSS 0.261283f
C14964 a_10796_42968# VSS 0.29877f
C14965 a_10835_43094# VSS 0.59174f
C14966 a_10518_42984# VSS 0.260322f
C14967 a_10083_42826# VSS 0.762957f
C14968 a_8952_43230# VSS 0.261046f
C14969 a_9127_43156# VSS 0.77314f
C14970 a_8387_43230# VSS 0.255573f
C14971 a_8605_42826# VSS 0.181157f
C14972 a_8037_42858# VSS 0.293593f
C14973 a_7765_42852# VSS 0.252651f
C14974 a_7871_42858# VSS 0.503534f
C14975 a_7227_42852# VSS 0.36607f
C14976 a_5755_42852# VSS 0.383967f
C14977 a_5111_42852# VSS 0.354197f
C14978 a_4520_42826# VSS 0.334784f
C14979 a_3935_42891# VSS 0.26911f
C14980 a_3681_42891# VSS 0.301094f
C14981 a_2905_42968# VSS 0.305424f
C14982 a_2075_43172# VSS 0.537699f
C14983 a_1847_42826# VSS 0.670072f
C14984 a_791_42968# VSS 0.335942f
C14985 a_685_42968# VSS 0.220885f
C14986 a_n1736_43218# VSS 0.073862f
C14987 a_n4318_38680# VSS 1.39087f
C14988 a_n3674_39304# VSS 1.06639f
C14989 a_n13_43084# VSS 0.368998f
C14990 a_n1076_43230# VSS 0.263204f
C14991 a_n901_43156# VSS 0.76245f
C14992 a_n1641_43230# VSS 0.256397f
C14993 a_n1423_42826# VSS 0.1805f
C14994 a_n1991_42858# VSS 0.295941f
C14995 a_n1853_43023# VSS 1.30078f
C14996 a_n2157_42858# VSS 0.556569f
C14997 a_n2472_42826# VSS 0.301801f
C14998 a_n2840_42826# VSS 0.327636f
C14999 a_20749_43396# VSS 0.253248f
C15000 a_17364_32525# VSS 1.89027f
C15001 a_22959_43396# VSS 0.345439f
C15002 a_14209_32519# VSS 2.01073f
C15003 a_22591_43396# VSS 0.335697f
C15004 a_13887_32519# VSS 1.94302f
C15005 a_22223_43396# VSS 0.333609f
C15006 a_5649_42852# VSS 1.95364f
C15007 a_13678_32519# VSS 2.06117f
C15008 a_21855_43396# VSS 0.334538f
C15009 a_4361_42308# VSS 1.30251f
C15010 a_13467_32519# VSS 2.22543f
C15011 a_19095_43396# VSS 0.132304f
C15012 a_21487_43396# VSS 0.293844f
C15013 a_743_42282# VSS 1.36822f
C15014 a_4190_30871# VSS 7.37921f
C15015 a_21259_43561# VSS 0.217667f
C15016 a_16823_43084# VSS 1.23251f
C15017 a_16664_43396# VSS 0.080001f
C15018 a_19700_43370# VSS 0.335707f
C15019 a_19268_43646# VSS 0.242693f
C15020 a_15743_43084# VSS 1.49489f
C15021 a_18783_43370# VSS 0.360096f
C15022 a_18525_43370# VSS 0.361236f
C15023 a_18429_43548# VSS 0.222219f
C15024 a_17324_43396# VSS 0.258017f
C15025 a_17499_43370# VSS 0.762886f
C15026 a_16759_43396# VSS 0.252915f
C15027 a_16977_43638# VSS 0.178776f
C15028 a_16409_43396# VSS 0.290743f
C15029 a_16547_43609# VSS 0.561468f
C15030 a_16243_43396# VSS 0.562369f
C15031 a_16137_43396# VSS 0.635905f
C15032 a_15781_43660# VSS 0.234761f
C15033 a_15681_43442# VSS 0.20154f
C15034 a_12281_43396# VSS 0.691406f
C15035 a_10341_43396# VSS 0.796012f
C15036 a_14955_43396# VSS 0.266041f
C15037 a_15095_43370# VSS 0.436411f
C15038 a_14205_43396# VSS 0.2933f
C15039 a_14358_43442# VSS 0.198188f
C15040 a_14579_43548# VSS 0.293668f
C15041 a_13667_43396# VSS 0.265557f
C15042 a_10695_43548# VSS 0.279385f
C15043 a_9803_43646# VSS 0.371929f
C15044 a_9145_43396# VSS 0.437647f
C15045 a_8685_43396# VSS 1.0146f
C15046 a_3457_43396# VSS 0.379621f
C15047 a_2813_43396# VSS 0.412407f
C15048 a_6452_43396# VSS 0.073862f
C15049 a_9396_43370# VSS 0.338475f
C15050 a_8791_43396# VSS 0.235222f
C15051 a_8147_43396# VSS 0.256103f
C15052 a_7112_43396# VSS 0.256956f
C15053 a_7287_43370# VSS 0.754599f
C15054 a_6547_43396# VSS 0.253718f
C15055 a_6765_43638# VSS 0.174622f
C15056 a_6197_43396# VSS 0.290517f
C15057 a_6293_42852# VSS 0.473619f
C15058 a_6031_43396# VSS 0.541083f
C15059 a_648_43396# VSS 0.231254f
C15060 a_3539_42460# VSS 0.337918f
C15061 a_3626_43646# VSS 1.9807f
C15062 a_2982_43646# VSS 3.25953f
C15063 a_n1557_42282# VSS 0.870257f
C15064 a_4905_42826# VSS 0.781685f
C15065 a_3080_42308# VSS 5.07131f
C15066 a_4699_43561# VSS 0.267684f
C15067 a_4235_43370# VSS 0.33553f
C15068 a_4093_43548# VSS 0.320586f
C15069 a_1756_43548# VSS 0.322408f
C15070 a_1568_43370# VSS 0.63594f
C15071 a_1049_43396# VSS 0.216408f
C15072 a_1209_43370# VSS 0.281234f
C15073 a_458_43396# VSS 0.252302f
C15074 a_n2012_43396# VSS 0.073862f
C15075 a_104_43370# VSS 0.297328f
C15076 a_n97_42460# VSS 6.9914f
C15077 a_n447_43370# VSS 0.269574f
C15078 a_n1352_43396# VSS 0.260107f
C15079 a_n1177_43370# VSS 0.478516f
C15080 a_n1917_43396# VSS 0.258245f
C15081 a_n1699_43638# VSS 0.175452f
C15082 a_n2267_43396# VSS 0.297246f
C15083 a_n2129_43609# VSS 1.07965f
C15084 a_n2433_43396# VSS 0.56533f
C15085 a_n4318_39304# VSS 0.959585f
C15086 a_n2840_43370# VSS 0.316787f
C15087 a_17538_32519# VSS 1.88404f
C15088 a_20974_43370# VSS 0.458091f
C15089 a_14401_32519# VSS 2.31932f
C15090 a_21381_43940# VSS 0.358332f
C15091 a_19319_43548# VSS 0.229395f
C15092 a_14021_43940# VSS 0.387813f
C15093 a_11173_44260# VSS 0.219946f
C15094 a_10555_44260# VSS 0.346315f
C15095 a_22959_43948# VSS 0.341565f
C15096 a_15493_43940# VSS 0.460801f
C15097 a_22223_43948# VSS 0.31992f
C15098 a_11341_43940# VSS 0.365183f
C15099 a_21115_43940# VSS 0.204633f
C15100 a_20935_43940# VSS 0.222887f
C15101 a_20623_43914# VSS 0.371294f
C15102 a_20365_43914# VSS 0.359455f
C15103 a_20269_44172# VSS 0.225063f
C15104 a_19862_44208# VSS 0.562087f
C15105 a_19478_44306# VSS 0.278384f
C15106 a_15493_43396# VSS 0.277875f
C15107 a_19328_44172# VSS 0.2031f
C15108 a_18451_43940# VSS 0.377396f
C15109 a_18326_43940# VSS 0.276559f
C15110 a_18079_43940# VSS 0.21121f
C15111 a_17973_43940# VSS 0.359917f
C15112 a_17737_43940# VSS 0.386318f
C15113 a_15682_43940# VSS 1.9643f
C15114 a_14955_43940# VSS 0.365393f
C15115 a_13483_43940# VSS 0.376442f
C15116 a_12429_44172# VSS 0.389129f
C15117 a_11750_44172# VSS 0.221782f
C15118 a_10807_43548# VSS 0.451031f
C15119 a_10949_43914# VSS 0.257331f
C15120 a_10729_43914# VSS 0.34307f
C15121 a_10405_44172# VSS 0.142993f
C15122 a_9672_43914# VSS 0.323006f
C15123 a_9028_43914# VSS 0.398016f
C15124 a_8333_44056# VSS 0.331632f
C15125 a_n2661_42282# VSS 1.51789f
C15126 a_3499_42826# VSS 0.380221f
C15127 a_n1644_44306# VSS 0.080042f
C15128 a_n3674_39768# VSS 0.890487f
C15129 a_n4318_39768# VSS 1.09976f
C15130 a_7845_44172# VSS 0.239173f
C15131 a_7542_44172# VSS 0.283767f
C15132 a_7281_43914# VSS 0.271121f
C15133 a_6453_43914# VSS 0.26639f
C15134 a_5663_43940# VSS 0.488325f
C15135 a_5495_43940# VSS 0.212229f
C15136 a_5013_44260# VSS 0.279924f
C15137 a_5244_44056# VSS 0.216368f
C15138 a_3905_42865# VSS 0.9893f
C15139 a_3600_43914# VSS 0.422049f
C15140 a_2998_44172# VSS 0.503048f
C15141 a_2889_44172# VSS 0.217034f
C15142 a_2675_43914# VSS 0.2974f
C15143 a_895_43940# VSS 0.237723f
C15144 a_2479_44172# VSS 0.817462f
C15145 a_2127_44172# VSS 0.517911f
C15146 a_453_43940# VSS 0.285192f
C15147 a_1414_42308# VSS 1.07452f
C15148 a_1467_44172# VSS 0.187431f
C15149 a_1115_44172# VSS 0.52592f
C15150 a_644_44056# VSS 0.227493f
C15151 a_175_44278# VSS 0.226801f
C15152 a_n984_44318# VSS 0.27358f
C15153 a_n809_44244# VSS 0.785904f
C15154 a_n1549_44318# VSS 0.264547f
C15155 a_n1331_43914# VSS 0.185087f
C15156 a_n1899_43946# VSS 0.299008f
C15157 a_n1761_44111# VSS 0.392075f
C15158 a_n2065_43946# VSS 0.658803f
C15159 a_n2472_43914# VSS 0.3103f
C15160 a_n2840_43914# VSS 0.345355f
C15161 a_19237_31679# VSS 1.48495f
C15162 a_22959_44484# VSS 0.343897f
C15163 a_17730_32519# VSS 2.44967f
C15164 a_22591_44484# VSS 0.315361f
C15165 a_22485_44484# VSS 0.590119f
C15166 a_20512_43084# VSS 0.561552f
C15167 a_22315_44484# VSS 0.238239f
C15168 a_3422_30871# VSS 8.519179f
C15169 a_21398_44850# VSS 0.073862f
C15170 a_18579_44172# VSS 0.812679f
C15171 a_19279_43940# VSS 1.69633f
C15172 a_20766_44850# VSS 0.177656f
C15173 a_20835_44721# VSS 0.260406f
C15174 a_20679_44626# VSS 0.58931f
C15175 a_20640_44752# VSS 0.296084f
C15176 a_20362_44736# VSS 0.255907f
C15177 a_20159_44458# VSS 0.483669f
C15178 a_19615_44636# VSS 0.238459f
C15179 a_11967_42832# VSS 6.11191f
C15180 a_19006_44850# VSS 0.073862f
C15181 a_17517_44484# VSS 0.244051f
C15182 a_14673_44172# VSS 0.290001f
C15183 a_11541_44484# VSS 0.139071f
C15184 a_15433_44458# VSS 0.301508f
C15185 a_14815_43914# VSS 0.445698f
C15186 a_n2293_43922# VSS 3.31971f
C15187 a_n2661_43922# VSS 1.51991f
C15188 a_n2661_42834# VSS 1.20196f
C15189 a_9159_44484# VSS 0.158168f
C15190 a_10617_44484# VSS 0.119149f
C15191 a_5708_44484# VSS 0.231649f
C15192 a_3363_44484# VSS 0.27629f
C15193 a_556_44484# VSS 0.201935f
C15194 a_9313_44734# VSS 1.31461f
C15195 a_5891_43370# VSS 2.82295f
C15196 a_8375_44464# VSS 0.211867f
C15197 a_7640_43914# VSS 0.542377f
C15198 a_6109_44484# VSS 0.648821f
C15199 a_n23_44458# VSS 0.278255f
C15200 a_n356_44636# VSS 2.91333f
C15201 a_n2012_44484# VSS 0.080001f
C15202 a_18989_43940# VSS 0.423174f
C15203 a_18374_44850# VSS 0.179731f
C15204 a_18443_44721# VSS 0.253971f
C15205 a_18287_44626# VSS 0.507939f
C15206 a_18248_44752# VSS 0.294917f
C15207 a_17970_44736# VSS 0.26161f
C15208 a_17767_44458# VSS 0.474097f
C15209 a_16979_44734# VSS 0.363013f
C15210 a_14539_43914# VSS 1.18088f
C15211 a_16112_44458# VSS 0.326339f
C15212 a_15004_44636# VSS 0.254778f
C15213 a_13720_44458# VSS 0.403209f
C15214 a_13076_44458# VSS 0.38829f
C15215 a_12883_44458# VSS 0.287544f
C15216 a_12607_44458# VSS 0.499331f
C15217 a_8975_43940# VSS 0.652857f
C15218 a_10057_43914# VSS 0.654189f
C15219 a_10440_44484# VSS 0.210149f
C15220 a_10334_44484# VSS 0.210217f
C15221 a_10157_44484# VSS 0.208916f
C15222 a_9838_44484# VSS 0.276258f
C15223 a_5883_43914# VSS 0.792825f
C15224 a_8701_44490# VSS 0.358059f
C15225 a_8103_44636# VSS 0.340824f
C15226 a_6298_44484# VSS 1.93814f
C15227 a_5518_44484# VSS 0.242995f
C15228 a_5343_44458# VSS 1.28071f
C15229 a_4743_44484# VSS 0.327178f
C15230 a_n699_43396# VSS 1.82142f
C15231 a_4223_44672# VSS 0.659279f
C15232 a_2779_44458# VSS 0.532137f
C15233 a_949_44458# VSS 1.97734f
C15234 a_742_44458# VSS 1.02263f
C15235 a_n452_44636# VSS 0.254732f
C15236 a_n1352_44484# VSS 0.269853f
C15237 a_n1177_44458# VSS 0.493891f
C15238 a_n1917_44484# VSS 0.280038f
C15239 a_n1699_44726# VSS 0.197478f
C15240 a_n2267_44484# VSS 0.308908f
C15241 a_n2129_44697# VSS 0.307327f
C15242 a_n2433_44484# VSS 0.679598f
C15243 a_n2661_44458# VSS 0.487677f
C15244 a_n4318_40392# VSS 0.995833f
C15245 a_n2840_44458# VSS 0.316322f
C15246 a_19721_31679# VSS 1.61824f
C15247 a_18114_32519# VSS 3.11898f
C15248 a_16237_45028# VSS 0.017944f
C15249 a_20193_45348# VSS 1.70015f
C15250 a_11691_44458# VSS 1.78467f
C15251 a_19113_45348# VSS 0.367248f
C15252 a_22959_45036# VSS 0.345334f
C15253 a_22223_45036# VSS 0.354178f
C15254 a_11827_44484# VSS 1.28091f
C15255 a_21359_45002# VSS 0.397791f
C15256 a_21101_45002# VSS 0.35202f
C15257 a_21005_45260# VSS 0.212992f
C15258 a_20567_45036# VSS 0.31908f
C15259 a_18494_42460# VSS 1.15626f
C15260 a_18184_42460# VSS 0.838573f
C15261 a_19778_44110# VSS 0.599421f
C15262 a_18911_45144# VSS 0.307008f
C15263 a_18587_45118# VSS 0.214925f
C15264 a_18315_45260# VSS 0.334834f
C15265 a_17719_45144# VSS 0.331229f
C15266 a_17613_45144# VSS 0.244364f
C15267 a_17023_45118# VSS 0.20885f
C15268 a_16922_45042# VSS 0.818675f
C15269 a_n2661_43370# VSS 0.820606f
C15270 a_8560_45348# VSS 0.185033f
C15271 a_n2293_42834# VSS 1.1151f
C15272 a_2304_45348# VSS 0.182367f
C15273 a_1423_45028# VSS 0.980773f
C15274 a_626_44172# VSS 0.67926f
C15275 a_375_42282# VSS 0.447027f
C15276 a_16751_45260# VSS 0.316547f
C15277 a_1307_43914# VSS 2.30311f
C15278 a_16019_45002# VSS 0.25377f
C15279 a_15595_45028# VSS 0.214111f
C15280 a_15415_45028# VSS 0.221991f
C15281 a_14797_45144# VSS 0.249222f
C15282 a_14537_43396# VSS 1.73146f
C15283 a_14180_45002# VSS 0.327485f
C15284 a_13777_45326# VSS 0.272936f
C15285 a_13556_45296# VSS 1.01916f
C15286 a_9482_43914# VSS 3.42654f
C15287 a_13348_45260# VSS 0.243533f
C15288 a_13159_45002# VSS 0.265737f
C15289 a_13017_45260# VSS 0.362048f
C15290 a_11963_45334# VSS 0.226884f
C15291 a_11787_45002# VSS 0.212512f
C15292 a_10951_45334# VSS 0.228638f
C15293 a_10775_45002# VSS 0.204487f
C15294 a_8953_45002# VSS 1.94941f
C15295 a_8191_45002# VSS 0.325964f
C15296 a_7705_45326# VSS 0.273009f
C15297 a_6709_45028# VSS 0.354418f
C15298 a_7229_43940# VSS 0.786182f
C15299 a_7276_45260# VSS 0.251523f
C15300 a_5205_44484# VSS 0.546179f
C15301 a_6431_45366# VSS 0.233718f
C15302 a_6171_45002# VSS 0.700605f
C15303 a_3232_43370# VSS 2.99721f
C15304 a_5691_45260# VSS 0.370273f
C15305 a_4927_45028# VSS 0.520892f
C15306 a_5111_44636# VSS 3.44603f
C15307 a_5147_45002# VSS 0.803306f
C15308 a_4558_45348# VSS 0.446148f
C15309 a_4574_45260# VSS 0.208274f
C15310 a_3537_45260# VSS 2.45782f
C15311 a_3429_45260# VSS 0.274034f
C15312 a_3065_45002# VSS 0.864786f
C15313 a_2680_45002# VSS 0.321351f
C15314 a_2382_45260# VSS 1.03422f
C15315 a_2274_45254# VSS 0.187307f
C15316 a_1667_45002# VSS 0.345429f
C15317 a_327_44734# VSS 0.419171f
C15318 a_413_45260# VSS 4.87522f
C15319 a_n37_45144# VSS 0.321746f
C15320 a_n143_45144# VSS 0.209896f
C15321 a_n467_45028# VSS 0.311181f
C15322 a_n967_45348# VSS 0.453992f
C15323 en_comp VSS 7.84057f
C15324 a_n2956_37592# VSS 2.90302f
C15325 a_n2810_45028# VSS 1.52635f
C15326 a_n745_45366# VSS 0.257282f
C15327 a_n913_45002# VSS 5.04725f
C15328 a_n1059_45260# VSS 2.30619f
C15329 a_n2017_45002# VSS 1.09013f
C15330 a_n2109_45247# VSS 0.252392f
C15331 a_n2293_45010# VSS 0.614925f
C15332 a_n2472_45002# VSS 0.298945f
C15333 a_n2661_45010# VSS 0.839496f
C15334 a_n2840_45002# VSS 0.340687f
C15335 a_20447_31679# VSS 1.49378f
C15336 a_22959_45572# VSS 0.34535f
C15337 a_19963_31679# VSS 1.43825f
C15338 a_22591_45572# VSS 0.363695f
C15339 a_3357_43084# VSS 2.42707f
C15340 a_19479_31679# VSS 1.67203f
C15341 a_22223_45572# VSS 0.334964f
C15342 a_2437_43646# VSS 6.25635f
C15343 a_21513_45002# VSS 0.669089f
C15344 a_20528_45572# VSS 0.073082f
C15345 a_21188_45572# VSS 0.284872f
C15346 a_21363_45546# VSS 0.515994f
C15347 a_20623_45572# VSS 0.256236f
C15348 a_20841_45814# VSS 0.180037f
C15349 a_20273_45572# VSS 0.288513f
C15350 a_20107_45572# VSS 0.541125f
C15351 a_17668_45572# VSS 0.217142f
C15352 a_18596_45572# VSS 0.073862f
C15353 a_19256_45572# VSS 0.257674f
C15354 a_19431_45546# VSS 0.487121f
C15355 a_18691_45572# VSS 0.255356f
C15356 a_18909_45814# VSS 0.178658f
C15357 a_18341_45572# VSS 0.291608f
C15358 a_18479_45785# VSS 1.15946f
C15359 a_18175_45572# VSS 0.516981f
C15360 a_16147_45260# VSS 0.506229f
C15361 a_16020_45572# VSS 0.073862f
C15362 a_17478_45572# VSS 0.232341f
C15363 a_15861_45028# VSS 0.449058f
C15364 a_8696_44636# VSS 0.917254f
C15365 a_16680_45572# VSS 0.258674f
C15366 a_16855_45546# VSS 0.471485f
C15367 a_16115_45572# VSS 0.253972f
C15368 a_16333_45814# VSS 0.178165f
C15369 a_15765_45572# VSS 0.291326f
C15370 a_15903_45785# VSS 0.4164f
C15371 a_15599_45572# VSS 0.50233f
C15372 a_15037_45618# VSS 0.209713f
C15373 a_11136_45572# VSS 0.17156f
C15374 a_9159_45572# VSS 0.151638f
C15375 a_8192_45572# VSS 0.17002f
C15376 a_11682_45822# VSS 0.010374f
C15377 a_10907_45822# VSS 0.547001f
C15378 a_10210_45822# VSS 0.012573f
C15379 a_15143_45578# VSS 0.315994f
C15380 a_14495_45572# VSS 0.325874f
C15381 a_13249_42308# VSS 1.08648f
C15382 a_13904_45546# VSS 0.327907f
C15383 a_13527_45546# VSS 0.245514f
C15384 a_13163_45724# VSS 0.180841f
C15385 a_12791_45546# VSS 0.237787f
C15386 a_11823_42460# VSS 2.45644f
C15387 a_12427_45724# VSS 0.190531f
C15388 a_11962_45724# VSS 0.218739f
C15389 a_11652_45724# VSS 0.258015f
C15390 a_11525_45546# VSS 0.346102f
C15391 a_11322_45546# VSS 0.62914f
C15392 a_10490_45724# VSS 0.972668f
C15393 a_8746_45002# VSS 0.547616f
C15394 a_10193_42453# VSS 3.59848f
C15395 a_10180_45724# VSS 0.281135f
C15396 a_10053_45546# VSS 0.373668f
C15397 a_9049_44484# VSS 0.249658f
C15398 a_7499_43078# VSS 3.22587f
C15399 a_8568_45546# VSS 0.317032f
C15400 a_8162_45546# VSS 0.376225f
C15401 a_7230_45938# VSS 0.078992f
C15402 a_4880_45572# VSS 0.182839f
C15403 a_3775_45552# VSS 0.209244f
C15404 a_7227_45028# VSS 0.439395f
C15405 a_6598_45938# VSS 0.185967f
C15406 a_6667_45809# VSS 0.264656f
C15407 a_6511_45714# VSS 0.647716f
C15408 a_6472_45840# VSS 0.310105f
C15409 a_6194_45824# VSS 0.2717f
C15410 a_5907_45546# VSS 0.592148f
C15411 a_5263_45724# VSS 0.250928f
C15412 a_4099_45572# VSS 0.33915f
C15413 a_2711_45572# VSS 1.77517f
C15414 a_2277_45546# VSS 0.303704f
C15415 a_1609_45822# VSS 0.5528f
C15416 a_n443_42852# VSS 4.64762f
C15417 a_509_45822# VSS 0.010571f
C15418 a_n23_45546# VSS 0.281189f
C15419 a_n356_45724# VSS 0.32306f
C15420 a_3503_45724# VSS 0.322319f
C15421 a_3316_45546# VSS 0.336134f
C15422 a_3218_45724# VSS 0.379893f
C15423 a_2957_45546# VSS 0.276358f
C15424 a_1848_45724# VSS 0.245258f
C15425 a_997_45618# VSS 0.248122f
C15426 a_n755_45592# VSS 5.8889f
C15427 a_n357_42282# VSS 2.46134f
C15428 a_310_45028# VSS 0.207165f
C15429 a_n1099_45572# VSS 0.339525f
C15430 a_380_45546# VSS 0.337145f
C15431 a_n452_45724# VSS 0.253614f
C15432 a_n863_45724# VSS 3.49288f
C15433 a_n1079_45724# VSS 0.289271f
C15434 a_n2293_45546# VSS 0.879703f
C15435 a_n2956_38216# VSS 1.49846f
C15436 a_n2472_45546# VSS 0.340801f
C15437 a_n2661_45546# VSS 1.58481f
C15438 a_n2810_45572# VSS 1.43198f
C15439 a_n2840_45546# VSS 0.344757f
C15440 a_20692_30879# VSS 1.62176f
C15441 a_20205_31679# VSS 1.45875f
C15442 a_19240_46482# VSS 0.073862f
C15443 a_16375_45002# VSS 1.44161f
C15444 a_13259_45724# VSS 4.49032f
C15445 a_14180_46482# VSS 0.073862f
C15446 a_12638_46436# VSS 0.162178f
C15447 a_12379_46436# VSS 0.275423f
C15448 a_10586_45546# VSS 0.542658f
C15449 a_8049_45260# VSS 0.741927f
C15450 a_8034_45724# VSS 0.299594f
C15451 a_5066_45546# VSS 0.436834f
C15452 a_n1925_42282# VSS 1.34109f
C15453 a_526_44458# VSS 6.44493f
C15454 a_2981_46116# VSS 0.091491f
C15455 a_n1736_46482# VSS 0.07565f
C15456 a_n2956_38680# VSS 1.34225f
C15457 a_n2956_39304# VSS 1.60721f
C15458 a_22959_46124# VSS 0.345245f
C15459 a_10809_44734# VSS 1.05002f
C15460 a_22223_46124# VSS 0.354467f
C15461 a_6945_45028# VSS 0.978274f
C15462 a_21137_46414# VSS 0.340736f
C15463 a_20708_46348# VSS 0.268156f
C15464 a_19900_46494# VSS 0.26164f
C15465 a_20075_46420# VSS 0.475201f
C15466 a_19335_46494# VSS 0.260378f
C15467 a_19553_46090# VSS 0.179968f
C15468 a_18985_46122# VSS 0.297132f
C15469 a_18819_46122# VSS 0.545109f
C15470 a_17957_46116# VSS 0.309446f
C15471 a_18189_46348# VSS 0.296366f
C15472 a_17715_44484# VSS 0.55862f
C15473 a_17583_46090# VSS 0.307562f
C15474 a_15682_46116# VSS 1.96743f
C15475 a_2324_44458# VSS 6.12227f
C15476 a_14840_46494# VSS 0.263367f
C15477 a_15015_46420# VSS 0.472948f
C15478 a_14275_46494# VSS 0.258968f
C15479 a_14493_46090# VSS 0.176122f
C15480 a_13925_46122# VSS 0.294602f
C15481 a_13759_46122# VSS 0.518292f
C15482 a_13351_46090# VSS 0.304427f
C15483 a_12594_46348# VSS 0.284494f
C15484 a_12005_46116# VSS 0.381711f
C15485 a_10903_43370# VSS 2.66576f
C15486 a_11387_46155# VSS 0.260117f
C15487 a_11133_46155# VSS 0.299642f
C15488 a_11189_46129# VSS 0.32558f
C15489 a_9290_44172# VSS 4.78398f
C15490 a_10355_46116# VSS 0.290668f
C15491 a_9823_46155# VSS 0.261206f
C15492 a_9569_46155# VSS 0.304755f
C15493 a_9625_46129# VSS 0.369694f
C15494 a_8953_45546# VSS 1.00397f
C15495 a_5937_45572# VSS 1.8333f
C15496 a_8199_44636# VSS 2.29742f
C15497 a_8349_46414# VSS 0.273442f
C15498 a_8016_46348# VSS 0.539696f
C15499 a_7920_46348# VSS 0.269852f
C15500 a_6419_46155# VSS 0.273686f
C15501 a_6165_46155# VSS 0.303989f
C15502 a_5497_46414# VSS 0.304684f
C15503 a_5204_45822# VSS 0.338817f
C15504 a_5164_46348# VSS 0.419282f
C15505 a_5068_46348# VSS 0.25855f
C15506 a_4704_46090# VSS 0.296767f
C15507 a_4419_46090# VSS 0.357571f
C15508 a_4185_45028# VSS 2.50496f
C15509 a_3699_46348# VSS 0.226584f
C15510 a_3483_46348# VSS 4.80498f
C15511 a_3147_46376# VSS 0.52775f
C15512 a_2804_46116# VSS 0.222855f
C15513 a_2698_46116# VSS 0.215567f
C15514 a_2521_46116# VSS 0.220999f
C15515 a_167_45260# VSS 1.32487f
C15516 a_2202_46116# VSS 0.273578f
C15517 a_1823_45246# VSS 2.36307f
C15518 a_1138_42852# VSS 0.456566f
C15519 a_1176_45822# VSS 0.278365f
C15520 a_1208_46090# VSS 0.348206f
C15521 a_805_46414# VSS 0.27506f
C15522 a_472_46348# VSS 0.32751f
C15523 a_376_46348# VSS 0.285607f
C15524 a_n1076_46494# VSS 0.262147f
C15525 a_n901_46420# VSS 0.762523f
C15526 a_n1641_46494# VSS 0.256945f
C15527 a_n1423_46090# VSS 0.176189f
C15528 a_n1991_46122# VSS 0.305274f
C15529 a_n1853_46287# VSS 0.341802f
C15530 a_n2157_46122# VSS 0.525314f
C15531 a_n2293_46098# VSS 0.690447f
C15532 a_n2472_46090# VSS 0.290925f
C15533 a_n2840_46090# VSS 0.340313f
C15534 a_21076_30879# VSS 2.20404f
C15535 a_22959_46660# VSS 0.338967f
C15536 a_12741_44636# VSS 0.979225f
C15537 a_20820_30879# VSS 1.70591f
C15538 a_22591_46660# VSS 0.292786f
C15539 a_11415_45002# VSS 1.63684f
C15540 a_20202_43084# VSS 1.05073f
C15541 a_22365_46825# VSS 0.208388f
C15542 a_18280_46660# VSS 0.29316f
C15543 a_17639_46660# VSS 0.308795f
C15544 a_20528_46660# VSS 0.07565f
C15545 a_22000_46634# VSS 0.295895f
C15546 a_21188_46660# VSS 0.261124f
C15547 a_21363_46634# VSS 0.488515f
C15548 a_20623_46660# VSS 0.258464f
C15549 a_20841_46902# VSS 0.180869f
C15550 a_20273_46660# VSS 0.309206f
C15551 a_20411_46873# VSS 0.393328f
C15552 a_20107_46660# VSS 0.575208f
C15553 a_19123_46287# VSS 0.477642f
C15554 a_18285_46348# VSS 0.577053f
C15555 a_765_45546# VSS 0.902406f
C15556 a_17339_46660# VSS 0.927636f
C15557 a_16721_46634# VSS 0.305539f
C15558 a_16388_46812# VSS 1.42609f
C15559 a_13059_46348# VSS 2.36107f
C15560 a_14513_46634# VSS 0.29862f
C15561 a_14180_46812# VSS 0.368158f
C15562 a_14035_46660# VSS 0.322858f
C15563 a_13885_46660# VSS 0.297377f
C15564 a_12156_46660# VSS 0.074642f
C15565 a_19692_46634# VSS 1.97188f
C15566 a_19466_46812# VSS 0.675335f
C15567 a_19333_46634# VSS 0.289568f
C15568 a_15227_44166# VSS 2.80559f
C15569 a_18834_46812# VSS 0.198054f
C15570 a_17609_46634# VSS 0.205547f
C15571 a_16292_46812# VSS 0.271203f
C15572 a_15559_46634# VSS 0.394779f
C15573 a_15368_46634# VSS 0.278142f
C15574 a_14976_45028# VSS 0.479565f
C15575 a_3090_45724# VSS 2.6372f
C15576 a_15009_46634# VSS 0.270859f
C15577 a_14084_46812# VSS 0.251005f
C15578 a_13607_46688# VSS 0.218935f
C15579 a_12816_46660# VSS 0.260317f
C15580 a_12991_46634# VSS 0.475827f
C15581 a_12251_46660# VSS 0.270927f
C15582 a_12469_46902# VSS 0.193369f
C15583 a_11901_46660# VSS 0.303844f
C15584 a_11813_46116# VSS 0.563718f
C15585 a_11735_46660# VSS 0.520568f
C15586 a_11186_47026# VSS 0.078586f
C15587 a_8270_45546# VSS 0.779033f
C15588 a_7832_46660# VSS 0.073862f
C15589 a_6969_46634# VSS 0.289597f
C15590 a_6755_46942# VSS 3.33348f
C15591 a_10249_46116# VSS 0.414443f
C15592 a_10554_47026# VSS 0.191251f
C15593 a_10623_46897# VSS 0.283572f
C15594 a_10467_46802# VSS 0.523954f
C15595 a_10428_46928# VSS 0.314538f
C15596 a_10150_46912# VSS 0.276624f
C15597 a_9863_46634# VSS 0.607398f
C15598 a_8492_46660# VSS 0.283316f
C15599 a_8667_46634# VSS 0.596387f
C15600 a_7927_46660# VSS 0.269867f
C15601 a_8145_46902# VSS 0.179735f
C15602 a_7577_46660# VSS 0.314978f
C15603 a_7715_46873# VSS 0.546182f
C15604 a_7411_46660# VSS 0.532412f
C15605 a_5257_43370# VSS 1.42323f
C15606 a_5072_46660# VSS 0.073862f
C15607 a_6540_46812# VSS 0.248814f
C15608 a_5732_46660# VSS 0.260482f
C15609 a_5907_46634# VSS 0.473347f
C15610 a_5167_46660# VSS 0.263586f
C15611 a_5385_46902# VSS 0.17737f
C15612 a_4817_46660# VSS 0.296797f
C15613 a_4955_46873# VSS 0.365781f
C15614 a_4651_46660# VSS 0.548065f
C15615 a_4646_46812# VSS 2.12519f
C15616 a_3877_44458# VSS 2.8543f
C15617 a_2864_46660# VSS 0.080001f
C15618 a_3524_46660# VSS 0.267612f
C15619 a_3699_46634# VSS 0.499647f
C15620 a_2959_46660# VSS 0.261026f
C15621 a_3177_46902# VSS 0.184239f
C15622 a_2609_46660# VSS 0.302878f
C15623 a_2443_46660# VSS 0.657702f
C15624 a_n2661_46098# VSS 2.05975f
C15625 a_1799_45572# VSS 0.30194f
C15626 a_491_47026# VSS 0.010533f
C15627 a_288_46660# VSS 0.075217f
C15628 a_1983_46706# VSS 0.205951f
C15629 a_2107_46812# VSS 1.13475f
C15630 a_948_46660# VSS 0.263413f
C15631 a_1123_46634# VSS 0.776627f
C15632 a_383_46660# VSS 0.269735f
C15633 a_601_46902# VSS 0.192316f
C15634 a_33_46660# VSS 0.309712f
C15635 a_171_46873# VSS 0.579977f
C15636 a_n133_46660# VSS 0.576523f
C15637 a_n2438_43548# VSS 2.99787f
C15638 a_n743_46660# VSS 3.29885f
C15639 a_n1021_46688# VSS 0.271211f
C15640 a_n1925_46634# VSS 1.33202f
C15641 a_n2312_38680# VSS 2.0221f
C15642 a_n2104_46634# VSS 0.340006f
C15643 a_n2293_46634# VSS 1.52366f
C15644 a_n2442_46660# VSS 1.32617f
C15645 a_n2472_46634# VSS 0.323981f
C15646 a_n2661_46634# VSS 0.742038f
C15647 a_n2956_39768# VSS 1.30197f
C15648 a_n2840_46634# VSS 0.328049f
C15649 a_22612_30879# VSS 3.41585f
C15650 a_21588_30879# VSS 2.80238f
C15651 a_20916_46384# VSS 0.827544f
C15652 a_20843_47204# VSS 0.121976f
C15653 a_19594_46812# VSS 0.277274f
C15654 a_19321_45002# VSS 1.15234f
C15655 a_13747_46662# VSS 2.11905f
C15656 a_13661_43548# VSS 2.82749f
C15657 a_5807_45002# VSS 2.5828f
C15658 a_15928_47570# VSS 0.075455f
C15659 a_768_44030# VSS 3.03052f
C15660 a_12549_44172# VSS 2.68201f
C15661 a_12891_46348# VSS 1.22195f
C15662 a_11309_47204# VSS 0.423399f
C15663 a_9804_47204# VSS 0.528639f
C15664 a_8128_46384# VSS 0.573494f
C15665 a_n881_46662# VSS 4.56296f
C15666 a_n1613_43370# VSS 4.90074f
C15667 a_2747_46873# VSS 0.287894f
C15668 a_n2312_39304# VSS 1.49307f
C15669 a_n2312_40392# VSS 2.25565f
C15670 a_22959_47212# VSS 0.322938f
C15671 a_11453_44696# VSS 0.689179f
C15672 SMPL_ON_N VSS 2.63208f
C15673 a_22731_47423# VSS 0.227778f
C15674 a_22223_47212# VSS 0.332189f
C15675 a_12465_44636# VSS 5.61685f
C15676 a_21811_47423# VSS 0.23358f
C15677 a_4883_46098# VSS 1.54736f
C15678 a_21496_47436# VSS 0.249536f
C15679 a_13507_46334# VSS 4.83848f
C15680 a_21177_47436# VSS 0.223524f
C15681 a_20990_47178# VSS 0.224581f
C15682 a_20894_47436# VSS 0.233111f
C15683 a_19787_47423# VSS 0.258015f
C15684 a_19386_47436# VSS 0.209882f
C15685 a_18597_46090# VSS 2.82344f
C15686 a_18780_47178# VSS 0.319719f
C15687 a_18479_47436# VSS 1.19826f
C15688 a_18143_47464# VSS 0.579061f
C15689 a_10227_46804# VSS 8.12328f
C15690 a_17591_47464# VSS 0.576556f
C15691 a_16588_47582# VSS 0.263715f
C15692 a_16763_47508# VSS 0.587861f
C15693 a_16023_47582# VSS 0.264352f
C15694 a_16327_47482# VSS 5.17799f
C15695 a_16241_47178# VSS 0.18232f
C15696 a_15673_47210# VSS 0.315684f
C15697 a_15811_47375# VSS 0.349499f
C15698 a_15507_47210# VSS 0.556554f
C15699 a_11599_46634# VSS 2.84967f
C15700 a_14955_47212# VSS 0.358339f
C15701 a_14311_47204# VSS 0.248858f
C15702 a_13487_47204# VSS 0.643275f
C15703 a_12861_44030# VSS 3.64545f
C15704 a_13717_47436# VSS 1.02478f
C15705 a_n1435_47204# VSS 9.72476f
C15706 a_13381_47204# VSS 0.225132f
C15707 a_11459_47204# VSS 0.553679f
C15708 a_9313_45822# VSS 1.04727f
C15709 a_11031_47542# VSS 0.247302f
C15710 a_9863_47436# VSS 0.265619f
C15711 a_9067_47204# VSS 0.606182f
C15712 a_6575_47204# VSS 0.798434f
C15713 a_7903_47542# VSS 0.258657f
C15714 a_7227_47204# VSS 0.610401f
C15715 a_6851_47204# VSS 0.346433f
C15716 a_6491_46660# VSS 0.343406f
C15717 a_6545_47178# VSS 0.597936f
C15718 a_6151_47436# VSS 2.12954f
C15719 a_5815_47464# VSS 0.594449f
C15720 a_5129_47502# VSS 0.361487f
C15721 a_4915_47217# VSS 2.79467f
C15722 a_n443_46116# VSS 4.167f
C15723 a_4791_45118# VSS 2.65418f
C15724 a_4700_47436# VSS 0.271201f
C15725 a_4007_47204# VSS 0.628996f
C15726 a_3815_47204# VSS 0.440491f
C15727 a_3785_47178# VSS 0.541893f
C15728 a_3381_47502# VSS 0.320926f
C15729 a_n1151_42308# VSS 3.78206f
C15730 a_3160_47472# VSS 0.607125f
C15731 a_2905_45572# VSS 0.47073f
C15732 a_2952_47436# VSS 0.275026f
C15733 a_2553_47502# VSS 0.294118f
C15734 a_2063_45854# VSS 1.92678f
C15735 a_584_46384# VSS 2.10508f
C15736 a_2124_47436# VSS 0.276508f
C15737 a_1431_47204# VSS 0.595895f
C15738 a_1239_47204# VSS 0.33333f
C15739 a_1209_47178# VSS 0.474725f
C15740 a_327_47204# VSS 0.581187f
C15741 a_n785_47204# VSS 0.361759f
C15742 a_n23_47502# VSS 0.278861f
C15743 a_n237_47217# VSS 3.05697f
C15744 a_n746_45260# VSS 0.993718f
C15745 a_n971_45724# VSS 4.81311f
C15746 a_n452_47436# VSS 0.28781f
C15747 a_n815_47178# VSS 0.513835f
C15748 a_n1605_47204# VSS 0.250546f
C15749 SMPL_ON_P VSS 4.99224f
C15750 a_n1741_47186# VSS 1.81488f
C15751 a_n1920_47178# VSS 0.310881f
C15752 a_n2109_47186# VSS 0.936844f
C15753 a_n2288_47178# VSS 0.346995f
C15754 a_n2497_47436# VSS 2.31207f
C15755 a_n2833_47464# VSS 0.602779f
C15756 w_10694_33990# VSS 53.0313f
C15757 w_1575_34786# VSS 53.144802f
.ends

