* NGSPICE file created from state_machine.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends


.subckt state_machine VDD VSS RST_Z START COMP_P COMP_N SAMPLE_O VCM_O[10] VCM_O[9] VCM_O[8] VCM_O[7] VCM_O[6] VCM_O[5] VCM_O[4] VCM_O[3] VCM_O[2]
+ VCM_O[1] VCM_O[0] EN_COMP VIN_P_SW_ON VIN_N_SW_ON VCM_DUMMY_O EN_VCM_SW_O EN_OFFSET_CAL OFFSET_CAL_CYCLE EN_OFFSET_CAL_O CLK_DATA DATA[5]
+ DATA[4] DATA[3] DATA[2] DATA[1] DATA[0] DEBUG_MUX[3] DEBUG_MUX[2] DEBUG_MUX[1] DEBUG_MUX[0] DEBUG_OUT VSS_N_O[10] VSS_N_O[9] VSS_N_O[8]
+ VSS_N_O[7] VSS_N_O[6] VSS_N_O[5] VSS_N_O[4] VSS_N_O[3] VSS_N_O[2] VSS_N_O[1] VSS_N_O[0] VREF_Z_N_O[10] VREF_Z_N_O[9] VREF_Z_N_O[8]
+ VREF_Z_N_O[7] VREF_Z_N_O[6] VREF_Z_N_O[5] VREF_Z_N_O[4] VREF_Z_N_O[3] VREF_Z_N_O[2] VREF_Z_N_O[1] VREF_Z_N_O[0] VSS_P_O[10] VSS_P_O[9]
+ VSS_P_O[8] VSS_P_O[7] VSS_P_O[6] VSS_P_O[5] VSS_P_O[4] VSS_P_O[3] VSS_P_O[2] VSS_P_O[1] VSS_P_O[0] VREF_Z_P_O[10] VREF_Z_P_O[9]
+ VREF_Z_P_O[8] VREF_Z_P_O[7] VREF_Z_P_O[6] VREF_Z_P_O[5] VREF_Z_P_O[4] VREF_Z_P_O[3] VREF_Z_P_O[2] VREF_Z_P_O[1] VREF_Z_P_O[0] CLK EN_VCM_SW_O_I
+ VCM_O_I[10] VCM_O_I[9] VCM_O_I[8] VCM_O_I[7] VCM_O_I[6] VCM_O_I[5] VCM_O_I[4] VCM_O_I[3] VCM_O_I[2] VCM_O_I[1] VCM_O_I[0] SINGLE_ENDED
X_363_ result\[11\] _106_ _141_ _142_ net105 VSS VSS VDD VDD _003_ sky130_fd_sc_hd__a32o_1
X_294_ _087_ _101_ VSS VSS VDD VDD net69 sky130_fd_sc_hd__or2_1
X_432_ net117 _000_ net112 VSS VSS VDD VDD counter_sample sky130_fd_sc_hd__dfrtp_1
Xfanout116 net118 VSS VSS VDD VDD net116 sky130_fd_sc_hd__buf_2
Xfanout105 _027_ VSS VSS VDD VDD net105 sky130_fd_sc_hd__buf_2
X_346_ counter\[5\] net100 VSS VSS VDD VDD net26 sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_8_66 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_415_ net116 _003_ net112 VSS VSS VDD VDD result\[11\] sky130_fd_sc_hd__dfrtp_1
X_277_ _029_ result\[9\] net98 net109 VSS VSS VDD VDD _094_ sky130_fd_sc_hd__o211a_1
X_200_ result\[1\] result\[7\] _051_ VSS VSS VDD VDD _053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_82 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_329_ _047_ _119_ _050_ net116 VSS VSS VDD VDD net34 sky130_fd_sc_hd__a211oi_2
XFILLER_0_6_17 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
*XANTENNA_5 net80 VSS VSS VDD VDD sky130_fd_sc_hd__diode_2
Xoutput31 net31 VSS VSS VDD VDD data[4] sky130_fd_sc_hd__clkbuf_4
Xoutput42 net42 VSS VSS VDD VDD vcm_o[1] sky130_fd_sc_hd__buf_2
Xoutput86 net86 VSS VSS VDD VDD vss_p_o[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_35 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput64 net64 VSS VSS VDD VDD vref_z_p_o[1] sky130_fd_sc_hd__buf_2
Xoutput53 net53 VSS VSS VDD VDD vref_z_n_o[1] sky130_fd_sc_hd__buf_2
Xoutput75 net75 VSS VSS VDD VDD vss_n_o[1] sky130_fd_sc_hd__buf_2
X_362_ net102 _075_ _140_ VSS VSS VDD VDD _142_ sky130_fd_sc_hd__and3_1
X_293_ result\[7\] result\[6\] net108 VSS VSS VDD VDD _101_ sky130_fd_sc_hd__mux2_1
X_431_ net117 _019_ net112 VSS VSS VDD VDD counter\[11\] sky130_fd_sc_hd__dfrtp_4
Xfanout117 net118 VSS VSS VDD VDD net117 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout106 net109 VSS VSS VDD VDD net106 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_120 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_9_275 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_67 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_414_ net115 _002_ net111 VSS VSS VDD VDD result\[2\] sky130_fd_sc_hd__dfrtp_1
X_345_ _050_ _132_ _107_ counter_sample VSS VSS VDD VDD _171_ sky130_fd_sc_hd__a2bb2o_1
X_276_ counter\[11\] net96 _074_ VSS VSS VDD VDD _093_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_256 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_14 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_4_94 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_259_ net56 _085_ VSS VSS VDD VDD net89 sky130_fd_sc_hd__nand2_1
X_328_ net105 counter\[1\] _118_ VSS VSS VDD VDD _119_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_6_Right_6 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
Xoutput32 net32 VSS VSS VDD VDD data[5] sky130_fd_sc_hd__clkbuf_4
Xoutput54 net54 VSS VSS VDD VDD vref_z_n_o[2] sky130_fd_sc_hd__buf_2
XFILLER_0_7_192 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
Xoutput43 net43 VSS VSS VDD VDD vcm_o[2] sky130_fd_sc_hd__buf_2
Xoutput87 net87 VSS VSS VDD VDD vss_p_o[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_36 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput76 net76 VSS VSS VDD VDD vss_n_o[2] sky130_fd_sc_hd__buf_2
Xoutput65 net65 VSS VSS VDD VDD vref_z_p_o[2] sky130_fd_sc_hd__buf_2
XFILLER_0_4_151 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_361_ net102 _075_ VSS VSS VDD VDD _141_ sky130_fd_sc_hd__nand2_1
X_292_ _068_ _100_ VSS VSS VDD VDD net68 sky130_fd_sc_hd__or2_1
XFILLER_0_7_61 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_430_ net117 _018_ net112 VSS VSS VDD VDD counter\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_195 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xfanout118 net1 VSS VSS VDD VDD net118 sky130_fd_sc_hd__clkbuf_2
Xfanout107 net109 VSS VSS VDD VDD net107 sky130_fd_sc_hd__clkbuf_2
X_413_ net115 _001_ net114 VSS VSS VDD VDD result\[6\] sky130_fd_sc_hd__dfrtp_2
X_275_ result\[10\] _074_ VSS VSS VDD VDD net61 sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_8_68 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_344_ _118_ _131_ counter\[7\] counter\[2\] VSS VSS VDD VDD _132_ sky130_fd_sc_hd__and4b_1
X_189_ net18 VSS VSS VDD VDD _043_ sky130_fd_sc_hd__inv_2
X_258_ result\[4\] _084_ net95 VSS VSS VDD VDD _085_ sky130_fd_sc_hd__o21ai_1
X_327_ net107 counter\[0\] VSS VSS VDD VDD _118_ sky130_fd_sc_hd__nor2_1
Xoutput33 net33 VSS VSS VDD VDD debug_out sky130_fd_sc_hd__clkbuf_4
Xoutput55 net55 VSS VSS VDD VDD vref_z_n_o[3] sky130_fd_sc_hd__buf_2
Xoutput44 net44 VSS VSS VDD VDD vcm_o[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_37 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput88 net88 VSS VSS VDD VDD vss_p_o[3] sky130_fd_sc_hd__buf_2
Xoutput77 net77 VSS VSS VDD VDD vss_n_o[3] sky130_fd_sc_hd__buf_2
Xoutput66 net66 VSS VSS VDD VDD vref_z_p_o[3] sky130_fd_sc_hd__buf_2
X_291_ result\[6\] result\[5\] net107 VSS VSS VDD VDD _100_ sky130_fd_sc_hd__mux2_1
X_360_ net3 _106_ VSS VSS VDD VDD _140_ sky130_fd_sc_hd__and2_1
Xfanout108 net109 VSS VSS VDD VDD net108 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_8_69 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_412_ _140_ _169_ _168_ VSS VSS VDD VDD _025_ sky130_fd_sc_hd__mux2_1
X_343_ counter\[1\] counter\[10\] counter\[8\] _130_ VSS VSS VDD VDD _131_ sky130_fd_sc_hd__and4_1
X_274_ result\[9\] _072_ _092_ VSS VSS VDD VDD net93 sky130_fd_sc_hd__a21o_1
XFILLER_0_6_225 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_326_ net7 _112_ _116_ VSS VSS VDD VDD _117_ sky130_fd_sc_hd__and3_1
X_188_ net15 VSS VSS VDD VDD _042_ sky130_fd_sc_hd__inv_2
X_257_ counter\[6\] net105 VSS VSS VDD VDD _084_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_209 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_309_ counter\[7\] _105_ VSS VSS VDD VDD net47 sky130_fd_sc_hd__nor2_1
Xoutput56 net56 VSS VSS VDD VDD vref_z_n_o[4] sky130_fd_sc_hd__buf_2
Xoutput45 net45 VSS VSS VDD VDD vcm_o[4] sky130_fd_sc_hd__buf_2
Xoutput34 net34 VSS VSS VDD VDD en_comp sky130_fd_sc_hd__buf_2
Xoutput89 net89 VSS VSS VDD VDD vss_p_o[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_38 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput78 net78 VSS VSS VDD VDD vss_n_o[4] sky130_fd_sc_hd__buf_2
Xoutput67 net67 VSS VSS VDD VDD vref_z_p_o[4] sky130_fd_sc_hd__buf_2
X_290_ _066_ _084_ _099_ VSS VSS VDD VDD net67 sky130_fd_sc_hd__or3_1
XFILLER_0_9_223 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xfanout109 single_ended_reg VSS VSS VDD VDD net109 sky130_fd_sc_hd__clkbuf_2
X_342_ net103 _033_ _129_ counter\[5\] counter\[6\] VSS VSS VDD VDD _130_ sky130_fd_sc_hd__o2111a_1
X_273_ _030_ result\[8\] net98 net108 VSS VSS VDD VDD _092_ sky130_fd_sc_hd__o211a_1
X_411_ _039_ _107_ VSS VSS VDD VDD _169_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_281 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_325_ net5 _113_ _115_ VSS VSS VDD VDD _116_ sky130_fd_sc_hd__a21bo_1
X_256_ result\[5\] _065_ VSS VSS VDD VDD net56 sky130_fd_sc_hd__nand2_1
X_187_ result\[10\] VSS VSS VDD VDD _041_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_8_Left_18 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_239_ result\[11\] net14 _075_ _059_ VSS VSS VDD VDD net74 sky130_fd_sc_hd__o31ai_1
X_308_ counter\[6\] _105_ VSS VSS VDD VDD net46 sky130_fd_sc_hd__nor2_1
XFILLER_0_1_54 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
Xoutput57 net57 VSS VSS VDD VDD vref_z_n_o[5] sky130_fd_sc_hd__buf_2
Xoutput46 net46 VSS VSS VDD VDD vcm_o[5] sky130_fd_sc_hd__buf_2
Xoutput35 net35 VSS VSS VDD VDD en_offset_cal_o sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_2_39 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput68 net68 VSS VSS VDD VDD vref_z_p_o[5] sky130_fd_sc_hd__buf_2
Xoutput79 net79 VSS VSS VDD VDD vss_n_o[5] sky130_fd_sc_hd__buf_2
XFILLER_0_7_97 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_4_187 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_0_1_179 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_1_157 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
X_272_ counter\[10\] net96 _072_ VSS VSS VDD VDD _091_ sky130_fd_sc_hd__a21o_1
X_410_ _137_ _158_ net107 VSS VSS VDD VDD _168_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_190 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_341_ counter\[3\] counter\[11\] net110 counter\[4\] VSS VSS VDD VDD _129_ sky130_fd_sc_hd__and4_1
X_324_ _034_ net5 _045_ net6 _114_ VSS VSS VDD VDD _115_ sky130_fd_sc_hd__o311a_1
X_186_ result\[9\] VSS VSS VDD VDD _040_ sky130_fd_sc_hd__inv_2
X_255_ net55 _083_ VSS VSS VDD VDD net88 sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_9_70 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_238_ net105 counter\[11\] VSS VSS VDD VDD _075_ sky130_fd_sc_hd__nand2_1
X_307_ counter\[5\] _105_ VSS VSS VDD VDD net45 sky130_fd_sc_hd__nor2_1
XFILLER_0_1_33 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xoutput58 net58 VSS VSS VDD VDD vref_z_n_o[6] sky130_fd_sc_hd__buf_2
Xoutput47 net47 VSS VSS VDD VDD vcm_o[6] sky130_fd_sc_hd__buf_2
Xoutput36 net36 VSS VSS VDD VDD en_vcm_sw_o sky130_fd_sc_hd__buf_2
Xoutput69 net69 VSS VSS VDD VDD vref_z_p_o[6] sky130_fd_sc_hd__buf_2
XFILLER_0_4_166 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_9_225 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_271_ result\[9\] _072_ VSS VSS VDD VDD net60 sky130_fd_sc_hd__nand2_1
X_340_ net12 _127_ _000_ VSS VSS VDD VDD _170_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_55 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_323_ net5 net4 counter\[6\] VSS VSS VDD VDD _114_ sky130_fd_sc_hd__or3b_1
X_254_ result\[3\] _082_ net95 VSS VSS VDD VDD _083_ sky130_fd_sc_hd__o21ai_1
X_185_ result\[3\] VSS VSS VDD VDD _039_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_9_71 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_275 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_306_ counter\[4\] _105_ VSS VSS VDD VDD net44 sky130_fd_sc_hd__nor2_1
X_237_ _041_ _074_ net96 VSS VSS VDD VDD net83 sky130_fd_sc_hd__a21o_1
Xoutput26 net26 VSS VSS VDD VDD clk_data sky130_fd_sc_hd__clkbuf_4
Xoutput59 net59 VSS VSS VDD VDD vref_z_n_o[7] sky130_fd_sc_hd__buf_2
Xoutput48 net48 VSS VSS VDD VDD vcm_o[7] sky130_fd_sc_hd__buf_2
Xoutput37 net37 VSS VSS VDD VDD offset_cal_cycle sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_7_11 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_40 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_270_ result\[8\] net97 _090_ VSS VSS VDD VDD net92 sky130_fd_sc_hd__a21o_1
X_399_ counter\[6\] net101 _082_ _159_ VSS VSS VDD VDD _160_ sky130_fd_sc_hd__a31o_1
X_322_ counter\[2\] counter\[0\] net4 VSS VSS VDD VDD _113_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_72 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_253_ net103 counter\[5\] VSS VSS VDD VDD _082_ sky130_fd_sc_hd__nor2_1
X_184_ result\[8\] VSS VSS VDD VDD _038_ sky130_fd_sc_hd__inv_2
X_305_ counter\[3\] _105_ VSS VSS VDD VDD net43 sky130_fd_sc_hd__nor2_1
X_236_ net23 _073_ VSS VSS VDD VDD _074_ sky130_fd_sc_hd__nor2_1
X_219_ _039_ _063_ net95 VSS VSS VDD VDD net76 sky130_fd_sc_hd__a21o_1
Xoutput27 net27 VSS VSS VDD VDD data[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_143 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xoutput49 net49 VSS VSS VDD VDD vcm_o[8] sky130_fd_sc_hd__buf_2
Xoutput38 net38 VSS VSS VDD VDD sample_o sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_135 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_41 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_160 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
X_398_ net106 _158_ VSS VSS VDD VDD _159_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_9_73 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_321_ _111_ _110_ _109_ VSS VSS VDD VDD _112_ sky130_fd_sc_hd__or3b_1
Xfanout95 _058_ VSS VSS VDD VDD net95 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_20 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_183_ result\[2\] VSS VSS VDD VDD _037_ sky130_fd_sc_hd__inv_2
X_252_ net107 _034_ net17 result\[4\] VSS VSS VDD VDD net55 sky130_fd_sc_hd__or4b_2
X_304_ counter\[2\] _105_ VSS VSS VDD VDD net42 sky130_fd_sc_hd__nor2_1
X_235_ net104 counter\[10\] VSS VSS VDD VDD _073_ sky130_fd_sc_hd__nand2_1
X_218_ net16 _062_ VSS VSS VDD VDD _063_ sky130_fd_sc_hd__nor2_1
Xoutput28 net28 VSS VSS VDD VDD data[1] sky130_fd_sc_hd__clkbuf_4
Xoutput39 net39 VSS VSS VDD VDD vcm_dummy_o sky130_fd_sc_hd__buf_2
XFILLER_0_1_106 VSS VSS VDD VDD sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_42 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_250 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_0_172 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_397_ counter\[4\] _050_ counter\[5\] VSS VSS VDD VDD _158_ sky130_fd_sc_hd__or3b_1
X_320_ counter\[7\] net5 net4 net6 VSS VSS VDD VDD _111_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_0_21 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout96 _058_ VSS VSS VDD VDD net96 sky130_fd_sc_hd__clkbuf_2
X_182_ result\[7\] VSS VSS VDD VDD _036_ sky130_fd_sc_hd__inv_2
X_251_ result\[3\] _063_ _081_ VSS VSS VDD VDD net87 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_9_74 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_13 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_303_ counter\[1\] _105_ VSS VSS VDD VDD net40 sky130_fd_sc_hd__nor2_1
X_234_ _040_ _072_ net96 VSS VSS VDD VDD net82 sky130_fd_sc_hd__a21o_1
X_217_ net103 counter\[3\] VSS VSS VDD VDD _062_ sky130_fd_sc_hd__nand2_1
Xoutput29 net29 VSS VSS VDD VDD data[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_91 VSS VSS VDD VDD sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_5_Right_5 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_43 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_396_ _157_ _140_ _156_ VSS VSS VDD VDD _021_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_22 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_181_ result\[1\] VSS VSS VDD VDD _035_ sky130_fd_sc_hd__inv_2
X_250_ _034_ result\[2\] net98 net106 VSS VSS VDD VDD _081_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_9_75 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_379_ _154_ net3 _153_ VSS VSS VDD VDD _007_ sky130_fd_sc_hd__mux2_1
X_302_ net104 net98 VSS VSS VDD VDD _105_ sky130_fd_sc_hd__nand2_4
X_233_ net22 _071_ VSS VSS VDD VDD _072_ sky130_fd_sc_hd__nor2_1
X_216_ _037_ _061_ net95 VSS VSS VDD VDD net75 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_3_44 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_141 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_395_ _036_ _107_ VSS VSS VDD VDD _157_ sky130_fd_sc_hd__nor2_1
X_180_ counter\[4\] VSS VSS VDD VDD _034_ sky130_fd_sc_hd__inv_2
Xfanout98 net39 VSS VSS VDD VDD net98 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_9_76 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_23 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_378_ result\[0\] _106_ VSS VSS VDD VDD _154_ sky130_fd_sc_hd__and2_1
X_301_ net104 _041_ net74 VSS VSS VDD VDD net63 sky130_fd_sc_hd__o21ai_1
X_232_ net104 net110 VSS VSS VDD VDD _071_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_6_55 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_215_ net103 counter\[2\] _042_ VSS VSS VDD VDD _061_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_169 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_4_128 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_7_38 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_394_ net108 net110 _032_ net102 _155_ VSS VSS VDD VDD _156_ sky130_fd_sc_hd__a41o_1
XFILLER_0_5_267 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_77 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout99 _133_ VSS VSS VDD VDD net99 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_0_24 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_377_ counter\[1\] net100 _118_ _152_ VSS VSS VDD VDD _153_ sky130_fd_sc_hd__a31o_1
X_231_ _038_ _070_ net96 VSS VSS VDD VDD net81 sky130_fd_sc_hd__a21o_1
XFILLER_0_5_82 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_300_ _093_ _104_ VSS VSS VDD VDD net72 sky130_fd_sc_hd__nand2_1
X_429_ net116 _017_ net112 VSS VSS VDD VDD counter\[9\] sky130_fd_sc_hd__dfrtp_1
Xinput1 clk VSS VSS VDD VDD net1 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_7_Left_17 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_56 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_214_ result\[1\] _060_ _059_ VSS VSS VDD VDD net73 sky130_fd_sc_hd__o21ai_2
XFILLER_0_7_126 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_4_118 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Right_9 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_393_ _026_ net103 counter\[8\] net101 VSS VSS VDD VDD _155_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_9_78 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_25 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_376_ counter\[1\] net100 net106 counter\[2\] VSS VSS VDD VDD _152_ sky130_fd_sc_hd__and4b_1
X_230_ net108 _032_ net21 VSS VSS VDD VDD _070_ sky130_fd_sc_hd__nor3_1
X_428_ net116 _016_ net113 VSS VSS VDD VDD counter\[8\] sky130_fd_sc_hd__dfrtp_4
X_359_ net3 _139_ _138_ VSS VSS VDD VDD _002_ sky130_fd_sc_hd__mux2_1
Xinput2 comp_n VSS VSS VDD VDD net2 sky130_fd_sc_hd__buf_1
XFILLER_0_9_190 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_57 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_213_ net106 net13 counter\[1\] VSS VSS VDD VDD _060_ sky130_fd_sc_hd__or3b_1
XFILLER_0_2_40 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xmax_cap97 _070_ VSS VSS VDD VDD net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_100 VSS VSS VDD VDD sky130_fd_sc_hd__decap_6
X_392_ net109 net11 _127_ VSS VSS VDD VDD _020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_203 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_26 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_280 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_79 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_375_ net3 _151_ _150_ VSS VSS VDD VDD _006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_228 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_5_51 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_358_ _037_ _107_ VSS VSS VDD VDD _139_ sky130_fd_sc_hd__nor2_1
X_427_ net116 _015_ net113 VSS VSS VDD VDD counter\[7\] sky130_fd_sc_hd__dfrtp_4
X_289_ result\[5\] result\[4\] net107 VSS VSS VDD VDD _099_ sky130_fd_sc_hd__mux2_1
Xinput3 comp_p VSS VSS VDD VDD net3 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_58 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_212_ net108 net98 VSS VSS VDD VDD _059_ sky130_fd_sc_hd__nand2_4
XFILLER_0_6_172 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_3_142 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_0_Right_0 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_8_256 VDD VSS VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_0_0_123 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_391_ state\[1\] counter\[11\] net102 VSS VSS VDD VDD _019_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_0_27 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_374_ _038_ _107_ VSS VSS VDD VDD _151_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_74 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
Xinput4 debug_mux[0] VSS VSS VDD VDD net4 sky130_fd_sc_hd__buf_2
X_288_ net103 result\[4\] _098_ VSS VSS VDD VDD net66 sky130_fd_sc_hd__a21o_1
X_357_ counter\[2\] _050_ _062_ _137_ net103 VSS VSS VDD VDD _138_ sky130_fd_sc_hd__o32a_1
X_426_ net118 _014_ net114 VSS VSS VDD VDD counter\[6\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_6_59 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_211_ net106 net98 VSS VSS VDD VDD _058_ sky130_fd_sc_hd__and2_1
X_409_ _106_ _167_ VSS VSS VDD VDD _024_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_20 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_0_135 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_8_268 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
X_390_ counter\[11\] _049_ _133_ counter\[10\] VSS VSS VDD VDD _018_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_28 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_373_ counter\[8\] _050_ _071_ _149_ net110 VSS VSS VDD VDD _150_ sky130_fd_sc_hd__o32a_1
XFILLER_0_5_97 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
Xinput5 debug_mux[1] VSS VSS VDD VDD net5 sky130_fd_sc_hd__buf_2
X_425_ net115 _013_ net111 VSS VSS VDD VDD counter\[5\] sky130_fd_sc_hd__dfrtp_2
X_287_ net106 result\[3\] _059_ _064_ _082_ VSS VSS VDD VDD _098_ sky130_fd_sc_hd__a221o_1
X_356_ counter\[3\] _051_ VSS VSS VDD VDD _137_ sky130_fd_sc_hd__or2_1
X_210_ net24 net25 _050_ VSS VSS VDD VDD net39 sky130_fd_sc_hd__nor3_1
X_408_ result\[5\] net3 _166_ VSS VSS VDD VDD _167_ sky130_fd_sc_hd__mux2_1
X_339_ _117_ _121_ _126_ _128_ VSS VSS VDD VDD net33 sky130_fd_sc_hd__o31a_1
XFILLER_0_2_76 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_3_111 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_3_122 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_5_217 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_29 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_372_ net105 _030_ _050_ VSS VSS VDD VDD _149_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_87 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_355_ _136_ net3 _135_ VSS VSS VDD VDD _001_ sky130_fd_sc_hd__mux2_1
X_424_ net115 _012_ net111 VSS VSS VDD VDD counter\[4\] sky130_fd_sc_hd__dfrtp_4
X_286_ _080_ _097_ VSS VSS VDD VDD net65 sky130_fd_sc_hd__nand2_1
Xinput6 debug_mux[2] VSS VSS VDD VDD net6 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_2_Left_12 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_338_ net5 net4 _127_ _120_ VSS VSS VDD VDD _128_ sky130_fd_sc_hd__or4b_1
X_269_ _031_ result\[7\] net98 net108 VSS VSS VDD VDD _090_ sky130_fd_sc_hd__o211a_1
X_407_ counter\[7\] net101 _084_ _165_ VSS VSS VDD VDD _166_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_7_60 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput20 vcm_o_i[6] VSS VSS VDD VDD net20 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_4_Right_4 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_7_281 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_371_ _140_ _148_ _147_ VSS VSS VDD VDD _005_ sky130_fd_sc_hd__mux2_1
X_440_ net118 _025_ net111 VSS VSS VDD VDD result\[3\] sky130_fd_sc_hd__dfrtp_2
X_354_ result\[6\] _106_ VSS VSS VDD VDD _136_ sky130_fd_sc_hd__and2_1
X_423_ net115 _011_ net111 VSS VSS VDD VDD counter\[3\] sky130_fd_sc_hd__dfrtp_4
X_285_ _037_ _039_ net103 VSS VSS VDD VDD _097_ sky130_fd_sc_hd__mux2_1
Xinput7 debug_mux[3] VSS VSS VDD VDD net7 sky130_fd_sc_hd__buf_1
XFILLER_0_9_162 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_199_ _052_ VSS VSS VDD VDD net27 sky130_fd_sc_hd__inv_2
X_406_ net107 counter\[5\] net101 counter\[6\] VSS VSS VDD VDD _165_ sky130_fd_sc_hd__and4bb_1
X_337_ state\[1\] state\[0\] VSS VSS VDD VDD _127_ sky130_fd_sc_hd__nor2_2
X_268_ net110 net96 net97 VSS VSS VDD VDD _089_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_7_61 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput10 rst_z VSS VSS VDD VDD net10 sky130_fd_sc_hd__clkbuf_1
Xinput21 vcm_o_i[7] VSS VSS VDD VDD net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_88 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_4_274 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_370_ _040_ _107_ VSS VSS VDD VDD _148_ sky130_fd_sc_hd__nor2_1
X_422_ net115 _010_ net111 VSS VSS VDD VDD counter\[2\] sky130_fd_sc_hd__dfrtp_4
X_284_ _078_ _096_ VSS VSS VDD VDD net64 sky130_fd_sc_hd__or2_1
X_353_ _026_ net108 counter\[8\] net101 _134_ VSS VSS VDD VDD _135_ sky130_fd_sc_hd__a41o_1
Xinput8 en_offset_cal VSS VSS VDD VDD net8 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_1_30 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_198_ result\[0\] result\[6\] _051_ VSS VSS VDD VDD _052_ sky130_fd_sc_hd__mux2_1
X_336_ _046_ net6 _123_ _125_ VSS VSS VDD VDD _126_ sky130_fd_sc_hd__a31o_1
X_405_ _164_ _140_ _163_ VSS VSS VDD VDD _023_ sky130_fd_sc_hd__mux2_1
X_267_ result\[8\] _070_ VSS VSS VDD VDD net59 sky130_fd_sc_hd__nand2_1
XFILLER_0_6_166 VSS VSS VDD VDD sky130_fd_sc_hd__decap_6
Xinput11 single_ended VSS VSS VDD VDD net11 sky130_fd_sc_hd__clkbuf_1
X_319_ net110 _044_ net4 VSS VSS VDD VDD _110_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_7_62 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput22 vcm_o_i[8] VSS VSS VDD VDD net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_169 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_8_228 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_8_206 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_421_ net115 _009_ net111 VSS VSS VDD VDD counter\[1\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_1_31 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 en_vcm_sw_o_i VSS VSS VDD VDD net9 sky130_fd_sc_hd__clkbuf_1
X_283_ result\[2\] result\[1\] net106 VSS VSS VDD VDD _096_ sky130_fd_sc_hd__mux2_1
X_352_ counter\[6\] net105 net101 counter\[7\] VSS VSS VDD VDD _134_ sky130_fd_sc_hd__and4b_1
X_335_ _044_ net102 _120_ _124_ VSS VSS VDD VDD _125_ sky130_fd_sc_hd__o211a_1
X_197_ counter\[4\] net100 VSS VSS VDD VDD _051_ sky130_fd_sc_hd__nand2_2
X_404_ result\[1\] _106_ VSS VSS VDD VDD _164_ sky130_fd_sc_hd__and2_1
X_266_ net58 _088_ VSS VSS VDD VDD net91 sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_6_Left_16 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
Xinput12 start VSS VSS VDD VDD net12 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_63 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_318_ _032_ net5 net4 _108_ VSS VSS VDD VDD _109_ sky130_fd_sc_hd__a211o_1
Xinput23 vcm_o_i[9] VSS VSS VDD VDD net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_126 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_249_ counter\[4\] net95 _063_ VSS VSS VDD VDD _080_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_129 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Right_8 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_0_80 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_1_9 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_32 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_420_ net116 _008_ net114 VSS VSS VDD VDD counter\[0\] sky130_fd_sc_hd__dfrtp_1
X_351_ net102 _119_ _107_ VSS VSS VDD VDD net36 sky130_fd_sc_hd__a21o_1
X_282_ net103 result\[1\] _095_ VSS VSS VDD VDD net62 sky130_fd_sc_hd__a21o_1
XFILLER_0_9_154 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_334_ net4 _106_ VSS VSS VDD VDD _124_ sky130_fd_sc_hd__nand2_1
X_403_ counter\[3\] net100 _076_ _162_ VSS VSS VDD VDD _163_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_135 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_2_15 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_196_ state\[0\] state\[1\] VSS VSS VDD VDD _050_ sky130_fd_sc_hd__nand2b_4
X_265_ _032_ result\[6\] net98 net108 VSS VSS VDD VDD _088_ sky130_fd_sc_hd__o211ai_1
Xinput24 vin_n_sw_on VSS VSS VDD VDD net24 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_64 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_317_ counter\[10\] net5 VSS VSS VDD VDD _108_ sky130_fd_sc_hd__nor2_1
Xinput13 vcm_o_i[0] VSS VSS VDD VDD net13 sky130_fd_sc_hd__clkbuf_1
X_179_ counter\[0\] VSS VSS VDD VDD _033_ sky130_fd_sc_hd__inv_2
X_248_ result\[3\] _063_ VSS VSS VDD VDD net54 sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_33 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_350_ state\[1\] state\[0\] VSS VSS VDD VDD _133_ sky130_fd_sc_hd__and2_1
X_281_ net106 result\[0\] _059_ _060_ _076_ VSS VSS VDD VDD _095_ sky130_fd_sc_hd__a221o_1
X_333_ net3 _044_ _045_ net2 _122_ VSS VSS VDD VDD _123_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_27 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_195_ state\[0\] state\[1\] VSS VSS VDD VDD _049_ sky130_fd_sc_hd__and2b_1
X_402_ net106 counter\[1\] net100 counter\[2\] VSS VSS VDD VDD _162_ sky130_fd_sc_hd__and4bb_1
X_264_ counter\[8\] net95 _069_ VSS VSS VDD VDD _087_ sky130_fd_sc_hd__a21oi_1
Xinput25 vin_p_sw_on VSS VSS VDD VDD net25 sky130_fd_sc_hd__buf_1
X_316_ counter_sample _106_ VSS VSS VDD VDD _000_ sky130_fd_sc_hd__nor2_1
Xinput14 vcm_o_i[10] VSS VSS VDD VDD net14 sky130_fd_sc_hd__clkbuf_1
X_247_ net53 _079_ VSS VSS VDD VDD net86 sky130_fd_sc_hd__nand2_1
X_178_ counter\[8\] VSS VSS VDD VDD _032_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_109 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_2_194 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_3_70 VSS VSS VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_7_264 VDD VSS VDD VSS sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_9_91 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_1_215 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_34 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_281 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_280_ _041_ _059_ net52 VSS VSS VDD VDD net85 sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_167 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_9_145 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_401_ _161_ net3 _160_ VSS VSS VDD VDD _022_ sky130_fd_sc_hd__mux2_1
X_332_ counter\[11\] net5 net4 VSS VSS VDD VDD _122_ sky130_fd_sc_hd__and3_1
X_194_ net9 VSS VSS VDD VDD _048_ sky130_fd_sc_hd__inv_2
X_263_ result\[7\] _069_ VSS VSS VDD VDD net58 sky130_fd_sc_hd__nand2_1
XFILLER_0_5_181 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
X_315_ _106_ VSS VSS VDD VDD _107_ sky130_fd_sc_hd__inv_2
Xinput15 vcm_o_i[1] VSS VSS VDD VDD net15 sky130_fd_sc_hd__clkbuf_1
X_246_ _028_ result\[1\] net98 net106 VSS VSS VDD VDD _079_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_3_118 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
X_177_ net110 VSS VSS VDD VDD _031_ sky130_fd_sc_hd__inv_2
X_229_ _036_ _069_ net95 VSS VSS VDD VDD net80 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_4_45 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_72 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_331_ net5 net4 net34 _120_ VSS VSS VDD VDD _121_ sky130_fd_sc_hd__and4_1
X_400_ result\[4\] _106_ VSS VSS VDD VDD _161_ sky130_fd_sc_hd__and2_1
X_193_ net8 VSS VSS VDD VDD _047_ sky130_fd_sc_hd__inv_2
X_262_ net57 _086_ VSS VSS VDD VDD net90 sky130_fd_sc_hd__nand2_1
Xinput16 vcm_o_i[2] VSS VSS VDD VDD net16 sky130_fd_sc_hd__clkbuf_1
X_245_ counter\[3\] net95 _061_ VSS VSS VDD VDD _078_ sky130_fd_sc_hd__a21oi_1
X_176_ counter\[10\] VSS VSS VDD VDD _030_ sky130_fd_sc_hd__inv_2
X_314_ state\[1\] state\[0\] VSS VSS VDD VDD _106_ sky130_fd_sc_hd__nand2b_4
X_228_ net20 counter\[7\] net104 VSS VSS VDD VDD _069_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_4_46 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_330_ net7 net6 VSS VSS VDD VDD _120_ sky130_fd_sc_hd__nor2_1
X_192_ net7 VSS VSS VDD VDD _046_ sky130_fd_sc_hd__inv_2
X_261_ _026_ result\[5\] net98 net107 VSS VSS VDD VDD _086_ sky130_fd_sc_hd__o211ai_1
X_175_ counter\[11\] VSS VSS VDD VDD _029_ sky130_fd_sc_hd__inv_2
X_313_ counter\[11\] _105_ VSS VSS VDD VDD net41 sky130_fd_sc_hd__nor2_1
Xinput17 vcm_o_i[3] VSS VSS VDD VDD net17 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_1_Left_11 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_244_ result\[2\] _061_ VSS VSS VDD VDD net53 sky130_fd_sc_hd__nand2_1
XFILLER_0_2_186 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_3_95 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_8_18 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_7_223 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_227_ result\[6\] _068_ _059_ VSS VSS VDD VDD net79 sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_234 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_47 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_85 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Right_3 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_260_ result\[6\] _067_ VSS VSS VDD VDD net57 sky130_fd_sc_hd__nand2_1
X_191_ net4 VSS VSS VDD VDD _045_ sky130_fd_sc_hd__inv_2
X_389_ counter\[10\] net102 _133_ counter\[9\] VSS VSS VDD VDD _017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_162 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_312_ counter\[10\] _105_ VSS VSS VDD VDD net50 sky130_fd_sc_hd__nor2_1
Xinput18 vcm_o_i[4] VSS VSS VDD VDD net18 sky130_fd_sc_hd__clkbuf_1
X_174_ counter\[3\] VSS VSS VDD VDD _028_ sky130_fd_sc_hd__inv_2
X_243_ net51 _077_ VSS VSS VDD VDD net84 sky130_fd_sc_hd__nand2_1
XFILLER_0_2_176 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_226_ counter\[7\] net96 _067_ VSS VSS VDD VDD _068_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_4_48 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_209_ _057_ VSS VSS VDD VDD net32 sky130_fd_sc_hd__inv_2
XFILLER_0_0_64 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_6_74 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_190_ net5 VSS VSS VDD VDD _044_ sky130_fd_sc_hd__inv_2
X_388_ net110 net102 net99 counter\[8\] VSS VSS VDD VDD _016_ sky130_fd_sc_hd__a22o_1
X_311_ net110 _105_ VSS VSS VDD VDD net49 sky130_fd_sc_hd__nor2_1
Xinput19 vcm_o_i[5] VSS VSS VDD VDD net19 sky130_fd_sc_hd__clkbuf_1
X_173_ net108 VSS VSS VDD VDD _027_ sky130_fd_sc_hd__inv_2
X_242_ result\[0\] _076_ net95 VSS VSS VDD VDD _077_ sky130_fd_sc_hd__o21ai_1
X_225_ net19 counter\[6\] net104 VSS VSS VDD VDD _067_ sky130_fd_sc_hd__and3b_1
XFILLER_0_7_225 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_49 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_208_ result\[5\] result\[11\] _051_ VSS VSS VDD VDD _057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_106 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_6_64 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_387_ counter\[8\] net102 net99 counter\[7\] VSS VSS VDD VDD _015_ sky130_fd_sc_hd__a22o_1
X_310_ counter\[8\] _105_ VSS VSS VDD VDD net48 sky130_fd_sc_hd__nor2_1
X_439_ net118 _024_ net114 VSS VSS VDD VDD result\[5\] sky130_fd_sc_hd__dfrtp_2
X_172_ counter\[7\] VSS VSS VDD VDD _026_ sky130_fd_sc_hd__inv_2
X_241_ net103 counter\[2\] VSS VSS VDD VDD _076_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_76 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_15 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_224_ result\[5\] _059_ _066_ VSS VSS VDD VDD net78 sky130_fd_sc_hd__a21oi_1
X_207_ _056_ VSS VSS VDD VDD net31 sky130_fd_sc_hd__inv_2
XFILLER_0_4_218 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_0_55 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Right_7 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_8_173 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_386_ counter\[7\] net101 net99 counter\[6\] VSS VSS VDD VDD _014_ sky130_fd_sc_hd__a22o_1
Xoutput90 net90 VSS VSS VDD VDD vss_p_o[5] sky130_fd_sc_hd__buf_2
XFILLER_0_5_110 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_5_198 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_240_ _035_ _060_ VSS VSS VDD VDD net51 sky130_fd_sc_hd__or2_1
XFILLER_0_3_44 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_3_66 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_3_99 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_369_ net110 _050_ _073_ _146_ counter\[10\] VSS VSS VDD VDD _147_ sky130_fd_sc_hd__o32a_1
X_438_ net115 _023_ net111 VSS VSS VDD VDD result\[1\] sky130_fd_sc_hd__dfrtp_4
Xfanout110 counter\[9\] VSS VSS VDD VDD net110 sky130_fd_sc_hd__buf_2
X_223_ net95 _065_ VSS VSS VDD VDD _066_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_260 VDD VSS VDD VSS sky130_ef_sc_hd__decap_12
X_206_ result\[4\] result\[10\] _051_ VSS VSS VDD VDD _056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_285 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_0_244 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_50 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_11 VSS VSS VDD VDD sky130_fd_sc_hd__decap_6
X_385_ counter\[6\] net100 net99 counter\[5\] VSS VSS VDD VDD _013_ sky130_fd_sc_hd__a22o_1
Xoutput80 net80 VSS VSS VDD VDD vss_n_o[6] sky130_fd_sc_hd__buf_2
Xoutput91 net91 VSS VSS VDD VDD vss_p_o[6] sky130_fd_sc_hd__buf_2
X_437_ net115 _022_ net111 VSS VSS VDD VDD result\[4\] sky130_fd_sc_hd__dfrtp_2
X_299_ _040_ _041_ net104 VSS VSS VDD VDD _104_ sky130_fd_sc_hd__mux2_1
X_368_ net104 _029_ _050_ VSS VSS VDD VDD _146_ sky130_fd_sc_hd__or3_1
Xfanout111 net114 VSS VSS VDD VDD net111 sky130_fd_sc_hd__clkbuf_4
Xfanout100 net101 VSS VSS VDD VDD net100 sky130_fd_sc_hd__buf_2
X_222_ net105 counter\[5\] _043_ VSS VSS VDD VDD _065_ sky130_fd_sc_hd__and3_1
X_205_ _055_ VSS VSS VDD VDD net30 sky130_fd_sc_hd__inv_2
XFILLER_0_9_44 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_0_201 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_51 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_120 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_8_186 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_384_ counter\[4\] net99 net26 VSS VSS VDD VDD _012_ sky130_fd_sc_hd__a21o_1
Xoutput70 net70 VSS VSS VDD VDD vref_z_p_o[7] sky130_fd_sc_hd__buf_2
Xoutput81 net81 VSS VSS VDD VDD vss_n_o[7] sky130_fd_sc_hd__buf_2
Xoutput92 net92 VSS VSS VDD VDD vss_p_o[7] sky130_fd_sc_hd__buf_2
X_367_ _140_ result\[10\] _145_ VSS VSS VDD VDD _004_ sky130_fd_sc_hd__mux2_1
X_436_ net116 _021_ net113 VSS VSS VDD VDD result\[7\] sky130_fd_sc_hd__dfrtp_2
X_298_ _091_ _103_ VSS VSS VDD VDD net71 sky130_fd_sc_hd__nand2_1
Xfanout112 net113 VSS VSS VDD VDD net112 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_57 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
Xfanout101 _049_ VSS VSS VDD VDD net101 sky130_fd_sc_hd__clkbuf_2
X_221_ result\[4\] _064_ _059_ VSS VSS VDD VDD net77 sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_9_Left_19 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
X_419_ net115 _007_ net111 VSS VSS VDD VDD result\[0\] sky130_fd_sc_hd__dfrtp_1
X_204_ result\[3\] result\[9\] _051_ VSS VSS VDD VDD _055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_34 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_52 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
*XANTENNA_1 net51 VSS VSS VDD VDD sky130_fd_sc_hd__diode_2
X_383_ counter\[4\] net100 net99 counter\[3\] VSS VSS VDD VDD _011_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_7 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xoutput60 net60 VSS VSS VDD VDD vref_z_n_o[8] sky130_fd_sc_hd__buf_2
Xoutput71 net71 VSS VSS VDD VDD vref_z_p_o[8] sky130_fd_sc_hd__buf_2
Xoutput82 net82 VSS VSS VDD VDD vss_n_o[8] sky130_fd_sc_hd__buf_2
Xoutput93 net93 VSS VSS VDD VDD vss_p_o[8] sky130_fd_sc_hd__buf_2
XFILLER_0_5_113 VSS VSS VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_0_5_135 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_366_ _127_ net99 _144_ VSS VSS VDD VDD _145_ sky130_fd_sc_hd__or3_1
X_435_ net117 _020_ net112 VSS VSS VDD VDD single_ended_reg sky130_fd_sc_hd__dfrtp_1
X_297_ _038_ _040_ net104 VSS VSS VDD VDD _103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_149 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
Xfanout113 net114 VSS VSS VDD VDD net113 sky130_fd_sc_hd__buf_2
Xfanout102 _049_ VSS VSS VDD VDD net102 sky130_fd_sc_hd__buf_2
X_220_ net107 _034_ net17 VSS VSS VDD VDD _064_ sky130_fd_sc_hd__or3_1
X_349_ net8 _119_ VSS VSS VDD VDD net37 sky130_fd_sc_hd__and2_1
X_418_ net116 _006_ net113 VSS VSS VDD VDD result\[8\] sky130_fd_sc_hd__dfrtp_2
X_203_ _054_ VSS VSS VDD VDD net29 sky130_fd_sc_hd__inv_2
XFILLER_0_3_244 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_3_277 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_53 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_225 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
*XANTENNA_2 net54 VSS VSS VDD VDD sky130_fd_sc_hd__diode_2
Xoutput61 net61 VSS VSS VDD VDD vref_z_n_o[9] sky130_fd_sc_hd__buf_2
Xoutput72 net72 VSS VSS VDD VDD vref_z_p_o[9] sky130_fd_sc_hd__buf_2
X_382_ counter\[3\] net100 net99 counter\[2\] VSS VSS VDD VDD _010_ sky130_fd_sc_hd__a22o_1
Xoutput50 net50 VSS VSS VDD VDD vcm_o[9] sky130_fd_sc_hd__buf_2
Xoutput94 net94 VSS VSS VDD VDD vss_p_o[9] sky130_fd_sc_hd__buf_2
Xoutput83 net83 VSS VSS VDD VDD vss_n_o[9] sky130_fd_sc_hd__buf_2
XFILLER_0_5_158 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
X_365_ counter\[10\] _075_ _143_ net102 VSS VSS VDD VDD _144_ sky130_fd_sc_hd__o211a_1
X_434_ net117 _171_ net113 VSS VSS VDD VDD state\[1\] sky130_fd_sc_hd__dfrtp_4
X_296_ _089_ _102_ VSS VSS VDD VDD net70 sky130_fd_sc_hd__nand2_1
XFILLER_0_3_15 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_9_261 VSS VSS VDD VDD sky130_fd_sc_hd__decap_8
Xfanout114 net10 VSS VSS VDD VDD net114 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_0_Left_10 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
Xfanout103 net105 VSS VSS VDD VDD net103 sky130_fd_sc_hd__buf_2
X_417_ net116 _005_ net112 VSS VSS VDD VDD result\[9\] sky130_fd_sc_hd__dfrtp_2
X_348_ net8 net112 VSS VSS VDD VDD net35 sky130_fd_sc_hd__and2_1
X_279_ net14 _075_ result\[11\] VSS VSS VDD VDD net52 sky130_fd_sc_hd__or3b_1
X_202_ result\[2\] result\[8\] _051_ VSS VSS VDD VDD _054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_234 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_54 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Right_2 VSS VSS VDD VDD sky130_fd_sc_hd__decap_3
*XANTENNA_3 net56 VSS VSS VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_0_8_156 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
Xoutput84 net84 VSS VSS VDD VDD vss_p_o[0] sky130_fd_sc_hd__buf_2
Xoutput40 net40 VSS VSS VDD VDD vcm_o[0] sky130_fd_sc_hd__buf_2
X_381_ counter\[2\] net100 net99 counter\[1\] VSS VSS VDD VDD _009_ sky130_fd_sc_hd__a22o_1
Xoutput73 net73 VSS VSS VDD VDD vss_n_o[0] sky130_fd_sc_hd__buf_2
Xoutput51 net51 VSS VSS VDD VDD vref_z_n_o[0] sky130_fd_sc_hd__buf_2
Xoutput62 net62 VSS VSS VDD VDD vref_z_p_o[0] sky130_fd_sc_hd__buf_2
X_433_ net117 _170_ net112 VSS VSS VDD VDD state\[0\] sky130_fd_sc_hd__dfrtp_2
X_295_ _036_ _038_ net104 VSS VSS VDD VDD _102_ sky130_fd_sc_hd__mux2_1
X_364_ net108 _029_ VSS VSS VDD VDD _143_ sky130_fd_sc_hd__nand2_1
Xfanout115 net118 VSS VSS VDD VDD net115 sky130_fd_sc_hd__buf_2
Xfanout104 net105 VSS VSS VDD VDD net104 sky130_fd_sc_hd__clkbuf_4
X_416_ net116 _004_ net112 VSS VSS VDD VDD result\[10\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_8_65 VSS VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_3 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
X_347_ state\[1\] _048_ _127_ counter\[11\] VSS VSS VDD VDD net38 sky130_fd_sc_hd__a211oi_2
X_278_ result\[10\] _074_ _094_ VSS VSS VDD VDD net94 sky130_fd_sc_hd__a21o_1
X_201_ _053_ VSS VSS VDD VDD net28 sky130_fd_sc_hd__inv_2
XFILLER_0_4_70 VSS VSS VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_9_26 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_0_8_146 VSS VSS VDD VDD sky130_fd_sc_hd__fill_2
*XANTENNA_4 net58 VSS VSS VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_0_6_38 VSS VSS VDD VDD sky130_fd_sc_hd__fill_1
Xoutput52 net52 VSS VSS VDD VDD vref_z_n_o[10] sky130_fd_sc_hd__buf_2
Xoutput30 net30 VSS VSS VDD VDD data[3] sky130_fd_sc_hd__clkbuf_4
X_380_ counter\[1\] net101 net99 counter\[0\] VSS VSS VDD VDD _008_ sky130_fd_sc_hd__a22o_1
Xoutput41 net41 VSS VSS VDD VDD vcm_o[10] sky130_fd_sc_hd__buf_2
Xoutput63 net63 VSS VSS VDD VDD vref_z_p_o[10] sky130_fd_sc_hd__buf_2
Xoutput85 net85 VSS VSS VDD VDD vss_p_o[10] sky130_fd_sc_hd__buf_2
Xoutput74 net74 VSS VSS VDD VDD vss_n_o[10] sky130_fd_sc_hd__buf_2
.ends

